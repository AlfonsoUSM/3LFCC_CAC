* NGSPICE file created from mag_files/POSTLAYOUT/pmos_flat_48x48.ext - technology: sky130A

.subckt mag_files/POSTLAYOUT/pmos_flat_48x48 G D PW S
X0 S.t4606 G.t0 D.t4511 S.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1 S.t4605 G.t1 D.t4510 S.t218 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2 S.t4604 G.t2 D.t4509 S.t218 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3 S.t4603 G.t3 D.t4508 S.t216 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4 S.t4602 G.t4 D.t4507 S.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X5 D.t4506 G.t5 S.t4601 S.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X6 S.t4600 G.t6 D.t4505 S.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X7 S.t4599 G.t7 D.t4504 S.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X8 S.t4598 G.t8 D.t4503 S.t158 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X9 S.t4597 G.t9 D.t4502 S.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X10 S.t4596 G.t10 D.t4501 S.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X11 S.t4595 G.t11 D.t4500 S.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X12 D.t4499 G.t12 S.t4594 S.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X13 D.t4498 G.t13 S.t4593 S.t139 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X14 D.t4497 G.t14 S.t4592 S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X15 S.t4591 G.t15 D.t4496 S.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X16 S.t4590 G.t16 D.t4495 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X17 S.t4589 G.t17 D.t4494 S.t209 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X18 D.t4493 G.t18 S.t4588 S.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X19 S.t4587 G.t19 D.t4492 S.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X20 S.t4586 G.t20 D.t4491 S.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X21 D.t4490 G.t21 S.t4585 S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X22 S.t4584 G.t22 D.t4489 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X23 D.t4488 G.t23 S.t4583 S.t406 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X24 D.t4487 G.t24 S.t4582 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X25 S.t4581 G.t25 D.t4486 S.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X26 D.t4485 G.t26 S.t4580 S.t538 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X27 D.t4484 G.t27 S.t4579 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X28 D.t4483 G.t28 S.t4578 S.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X29 S.t4577 G.t29 D.t4482 S.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X30 S.t4576 G.t30 D.t4481 S.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X31 D.t4480 G.t31 S.t4575 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X32 D.t4479 G.t32 S.t4574 S.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X33 S.t4573 G.t33 D.t4478 S.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X34 S.t4572 G.t34 D.t4477 S.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X35 S.t4571 G.t35 D.t4476 S.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X36 S.t4570 G.t36 D.t4475 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X37 S.t4569 G.t37 D.t4474 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X38 D.t4473 G.t38 S.t4568 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X39 S.t4567 G.t39 D.t4472 S.t176 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X40 D.t4471 G.t40 S.t4566 S.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X41 S.t4565 G.t41 D.t4470 S.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X42 D.t4469 G.t42 S.t4564 S.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X43 D.t4468 G.t43 S.t4563 S.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X44 D.t4467 G.t44 S.t4562 S.t270 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X45 D.t4466 G.t45 S.t4561 S.t332 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X46 D.t4465 G.t46 S.t4560 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X47 S.t4559 G.t47 D.t4464 S.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X48 D.t4463 G.t48 S.t4558 S.t231 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X49 D.t4462 G.t49 S.t4557 S.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X50 S.t4556 G.t50 D.t4461 S.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X51 D.t2208 G.t51 S.t4555 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X52 D.t2207 G.t52 S.t4554 S.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X53 D.t2206 G.t53 S.t4553 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X54 S.t4552 G.t54 D.t2205 S.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X55 S.t4551 G.t55 D.t2204 S.t158 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X56 D.t2203 G.t56 S.t4550 S.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X57 D.t2202 G.t57 S.t4549 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X58 D.t2201 G.t58 S.t4548 S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X59 D.t2200 G.t59 S.t4547 S.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X60 S.t4546 G.t60 D.t2199 S.t388 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X61 D.t2198 G.t61 S.t4545 S.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X62 S.t4544 G.t62 D.t2197 S.t150 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X63 D.t2196 G.t63 S.t4543 S.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X64 S.t4542 G.t64 D.t2195 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X65 D.t2194 G.t65 S.t4541 S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X66 D.t2193 G.t66 S.t4540 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X67 S.t4539 G.t67 D.t2192 S.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X68 S.t4538 G.t68 D.t2191 S.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X69 S.t4537 G.t69 D.t2190 S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X70 S.t4536 G.t70 D.t2189 S.t357 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X71 D.t2188 G.t71 S.t4535 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X72 S.t4534 G.t72 D.t2187 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X73 D.t2186 G.t73 S.t4533 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X74 D.t2185 G.t74 S.t4532 S.t79 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X75 S.t4531 G.t75 D.t2184 S.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X76 D.t2183 G.t76 S.t4530 S.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X77 D.t2182 G.t77 S.t4529 S.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X78 S.t4528 G.t78 D.t2181 S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X79 S.t4527 G.t79 D.t2180 S.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X80 S.t4526 G.t80 D.t2179 S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X81 S.t4525 G.t81 D.t2178 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X82 S.t4524 G.t82 D.t2177 S.t321 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X83 D.t2176 G.t83 S.t4523 S.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X84 S.t4522 G.t84 D.t2175 S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X85 S.t4521 G.t85 D.t2174 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X86 D.t2173 G.t86 S.t4520 S.t79 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X87 S.t4519 G.t87 D.t2172 S.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X88 S.t4518 G.t88 D.t2171 S.t218 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X89 S.t4517 G.t89 D.t2170 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X90 D.t2169 G.t90 S.t4516 S.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X91 S.t4515 G.t91 D.t2168 S.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X92 S.t4514 G.t92 D.t2167 S.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X93 S.t4513 G.t93 D.t2166 S.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X94 D.t2165 G.t94 S.t4512 S.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X95 S.t4511 G.t95 D.t2164 S.t183 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X96 D.t2163 G.t96 S.t4510 S.t139 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X97 D.t2162 G.t97 S.t4509 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X98 D.t2161 G.t98 S.t4508 S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X99 S.t4507 G.t99 D.t2160 S.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X100 D.t2159 G.t100 S.t4506 S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X101 S.t4505 G.t101 D.t2158 S.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X102 D.t2157 G.t102 S.t4504 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X103 D.t2156 G.t103 S.t4503 S.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X104 S.t4502 G.t104 D.t2155 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X105 D.t2154 G.t105 S.t4501 S.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X106 S.t4500 G.t106 D.t2153 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X107 S.t4499 G.t107 D.t2152 S.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X108 D.t2151 G.t108 S.t4498 S.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X109 D.t4042 G.t109 S.t4497 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X110 D.t4041 G.t110 S.t4496 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X111 S.t4495 G.t111 D.t4040 S.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X112 S.t4494 G.t112 D.t4039 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X113 D.t4038 G.t113 S.t4493 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X114 S.t4492 G.t114 D.t4037 S.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X115 S.t4491 G.t115 D.t4036 S.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X116 D.t4035 G.t116 S.t4490 S.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X117 D.t4034 G.t117 S.t4489 S.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X118 S.t4488 G.t118 D.t4033 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X119 S.t4487 G.t119 D.t4032 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X120 S.t4486 G.t120 D.t4031 S.t79 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X121 S.t4485 G.t121 D.t4030 S.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X122 S.t4484 G.t122 D.t4029 S.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X123 S.t4483 G.t123 D.t4028 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X124 D.t4027 G.t124 S.t4482 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X125 S.t4481 G.t125 D.t4026 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X126 S.t4480 G.t126 D.t4025 S.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X127 D.t4024 G.t127 S.t4479 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X128 D.t4023 G.t128 S.t4478 S.t150 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X129 S.t4477 G.t129 D.t4022 S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X130 S.t4476 G.t130 D.t4021 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X131 D.t4020 G.t131 S.t4475 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X132 D.t4019 G.t132 S.t4474 S.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X133 S.t4473 G.t133 D.t4018 S.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X134 D.t4017 G.t134 S.t4472 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X135 S.t4471 G.t135 D.t4016 S.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X136 D.t4015 G.t136 S.t4470 S.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X137 D.t4014 G.t137 S.t4469 S.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X138 S.t4468 G.t138 D.t4013 S.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X139 D.t4012 G.t139 S.t4467 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X140 D.t4011 G.t140 S.t4466 S.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X141 D.t4010 G.t141 S.t4465 S.t218 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X142 S.t4464 G.t142 D.t4009 S.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X143 S.t4463 G.t143 D.t4008 S.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X144 D.t4007 G.t144 S.t4462 S.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X145 S.t4461 G.t145 D.t4006 S.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X146 D.t4005 G.t146 S.t4460 S.t443 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X147 D.t4004 G.t147 S.t4459 S.t158 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X148 D.t4003 G.t148 S.t4458 S.t270 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X149 D.t4002 G.t149 S.t4457 S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X150 S.t4456 G.t150 D.t4001 S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X151 D.t4000 G.t151 S.t4455 S.t209 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X152 D.t3999 G.t152 S.t4454 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X153 S.t4453 G.t153 D.t3998 S.t388 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X154 S.t4452 G.t154 D.t3997 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X155 D.t3996 G.t155 S.t4451 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X156 D.t3995 G.t156 S.t4450 S.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X157 D.t3994 G.t157 S.t4449 S.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X158 D.t3993 G.t158 S.t4448 S.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X159 S.t4447 G.t159 D.t3992 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X160 D.t3991 G.t160 S.t4446 S.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X161 D.t3990 G.t161 S.t4445 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X162 D.t3989 G.t162 S.t4444 S.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X163 D.t3988 G.t163 S.t4443 S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X164 S.t4442 G.t164 D.t3987 S.t538 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X165 D.t3986 G.t165 S.t4441 S.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X166 S.t4440 G.t166 D.t2548 S.t218 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X167 D.t2547 G.t167 S.t4439 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X168 D.t2546 G.t168 S.t4438 S.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X169 D.t2545 G.t169 S.t4437 S.t79 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X170 D.t2544 G.t170 S.t4436 S.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X171 S.t4435 G.t171 D.t2543 S.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X172 D.t2542 G.t172 S.t4434 S.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X173 D.t2541 G.t173 S.t4433 S.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X174 S.t4432 G.t174 D.t2540 S.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X175 S.t4431 G.t175 D.t2539 S.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X176 S.t4430 G.t176 D.t2538 S.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X177 S.t4429 G.t177 D.t2537 S.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X178 S.t4428 G.t178 D.t2536 S.t321 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X179 D.t2535 G.t179 S.t4427 S.t139 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X180 S.t4426 G.t180 D.t2534 S.t158 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X181 D.t2533 G.t181 S.t4425 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X182 D.t2532 G.t182 S.t4424 S.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X183 S.t4423 G.t183 D.t2531 S.t209 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X184 D.t2530 G.t184 S.t4422 S.t79 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X185 S.t4421 G.t185 D.t2529 S.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X186 D.t2528 G.t186 S.t4420 S.t216 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X187 S.t4419 G.t187 D.t2527 S.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X188 S.t4418 G.t188 D.t2526 S.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X189 D.t2525 G.t189 S.t4417 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X190 S.t4416 G.t190 D.t2524 S.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X191 D.t2523 G.t191 S.t4415 S.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X192 D.t2070 G.t192 S.t4414 S.t406 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X193 D.t2069 G.t193 S.t4413 S.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X194 D.t2068 G.t194 S.t4412 S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X195 D.t2067 G.t195 S.t4411 S.t198 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X196 S.t4410 G.t196 D.t2066 S.t176 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X197 D.t2065 G.t197 S.t4409 S.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X198 D.t2064 G.t198 S.t4408 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X199 D.t2063 G.t199 S.t4407 S.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X200 S.t4406 G.t200 D.t2062 S.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X201 D.t2061 G.t201 S.t4405 S.t332 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X202 S.t4404 G.t202 D.t2060 S.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X203 D.t2059 G.t203 S.t4403 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X204 D.t2058 G.t204 S.t4402 S.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X205 D.t2057 G.t205 S.t4401 S.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X206 D.t2056 G.t206 S.t4400 S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X207 D.t2055 G.t207 S.t4399 S.t150 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X208 S.t4398 G.t208 D.t2054 S.t176 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X209 D.t2053 G.t209 S.t4397 S.t198 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X210 D.t2052 G.t210 S.t4396 S.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X211 S.t4395 G.t211 D.t2051 S.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X212 D.t2050 G.t212 S.t4394 S.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X213 S.t4393 G.t213 D.t2049 S.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X214 D.t2048 G.t214 S.t4392 S.t332 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X215 D.t2047 G.t215 S.t4391 S.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X216 D.t2046 G.t216 S.t4390 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X217 S.t4389 G.t217 D.t779 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X218 D.t778 G.t218 S.t4388 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X219 D.t777 G.t219 S.t4387 S.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X220 D.t776 G.t220 S.t4386 S.t231 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X221 S.t4385 G.t221 D.t775 S.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X222 D.t774 G.t222 S.t4384 S.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X223 S.t4383 G.t223 D.t773 S.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X224 D.t772 G.t224 S.t4382 S.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X225 S.t4381 G.t225 D.t771 S.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X226 D.t770 G.t226 S.t4380 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X227 D.t769 G.t227 S.t4379 S.t443 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X228 D.t768 G.t228 S.t4378 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X229 D.t767 G.t229 S.t4377 S.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X230 S.t4376 G.t230 D.t766 S.t158 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X231 D.t765 G.t231 S.t4375 S.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X232 D.t764 G.t232 S.t4374 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X233 D.t763 G.t233 S.t4373 S.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X234 D.t762 G.t234 S.t4372 S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X235 D.t761 G.t235 S.t4371 S.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X236 D.t760 G.t236 S.t4370 S.t218 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X237 S.t4369 G.t237 D.t759 S.t388 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X238 D.t717 G.t238 S.t4368 S.t218 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X239 S.t4367 G.t239 D.t716 S.t443 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X240 S.t4366 G.t240 D.t715 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X241 D.t714 G.t241 S.t4365 S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X242 D.t713 G.t242 S.t4364 S.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X243 D.t712 G.t243 S.t4363 S.t158 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X244 S.t4362 G.t244 D.t711 S.t209 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X245 S.t4361 G.t245 D.t710 S.t139 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X246 D.t709 G.t246 S.t4360 S.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X247 D.t708 G.t247 S.t4359 S.t209 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X248 S.t4358 G.t248 D.t707 S.t357 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X249 D.t706 G.t249 S.t4357 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X250 S.t4356 G.t250 D.t705 S.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X251 D.t704 G.t251 S.t4355 S.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X252 D.t703 G.t252 S.t4354 S.t79 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X253 D.t702 G.t253 S.t4353 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X254 S.t4352 G.t254 D.t701 S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X255 D.t700 G.t255 S.t4351 S.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X256 D.t699 G.t256 S.t4350 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X257 S.t4349 G.t257 D.t698 S.t321 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X258 D.t64 G.t258 S.t4348 S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X259 D.t63 G.t259 S.t4347 S.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X260 D.t62 G.t260 S.t4346 S.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X261 D.t61 G.t261 S.t4345 S.t79 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X262 D.t60 G.t262 S.t4344 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X263 S.t4343 G.t263 D.t59 S.t332 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X264 D.t58 G.t264 S.t4342 S.t216 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X265 D.t57 G.t265 S.t4341 S.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X266 D.t56 G.t266 S.t4340 S.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X267 D.t55 G.t267 S.t4339 S.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X268 D.t54 G.t268 S.t4338 S.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X269 S.t4337 G.t269 D.t53 S.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X270 D.t52 G.t270 S.t4336 S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X271 S.t4335 G.t271 D.t51 S.t183 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X272 S.t4334 G.t272 D.t50 S.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X273 D.t49 G.t273 S.t4333 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X274 S.t4332 G.t274 D.t48 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X275 S.t4331 G.t275 D.t47 S.t198 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X276 D.t46 G.t276 S.t4330 S.t176 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X277 D.t1701 G.t277 S.t4329 S.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X278 D.t1700 G.t278 S.t4328 S.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X279 S.t4327 G.t279 D.t1699 S.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X280 S.t4326 G.t280 D.t1698 S.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X281 S.t4325 G.t281 D.t1697 S.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X282 D.t1696 G.t282 S.t4324 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X283 D.t1695 G.t283 S.t4323 S.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X284 S.t4322 G.t284 D.t1694 S.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X285 S.t4321 G.t285 D.t1693 S.t176 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X286 D.t1692 G.t286 S.t4320 S.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X287 D.t1691 G.t287 S.t4319 S.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X288 S.t4318 G.t288 D.t1690 S.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X289 S.t4317 G.t289 D.t1689 S.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X290 D.t1688 G.t290 S.t4316 S.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X291 S.t4315 G.t291 D.t1687 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X292 D.t1686 G.t292 S.t4314 S.t158 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X293 S.t4313 G.t293 D.t1685 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X294 D.t1684 G.t294 S.t4312 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X295 D.t1683 G.t295 S.t4311 S.t332 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X296 D.t1384 G.t296 S.t4310 S.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X297 D.t1383 G.t297 S.t4309 S.t388 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X298 S.t4308 G.t298 D.t1382 S.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X299 D.t1381 G.t299 S.t4307 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X300 D.t1380 G.t300 S.t4306 S.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X301 S.t4305 G.t301 D.t1379 S.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X302 D.t1378 G.t302 S.t4304 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X303 S.t4303 G.t303 D.t1377 S.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X304 D.t1376 G.t304 S.t4302 S.t150 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X305 S.t4301 G.t305 D.t1375 S.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X306 D.t1374 G.t306 S.t4300 S.t198 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X307 D.t1373 G.t307 S.t4299 S.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X308 D.t1372 G.t308 S.t4298 S.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X309 S.t4297 G.t309 D.t1371 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X310 D.t1370 G.t310 S.t4296 S.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X311 S.t4295 G.t311 D.t3900 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X312 D.t3899 G.t312 S.t4294 S.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X313 D.t3898 G.t313 S.t4293 S.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X314 S.t4292 G.t314 D.t3897 S.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X315 S.t4291 G.t315 D.t3896 S.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X316 D.t3895 G.t316 S.t4290 S.t443 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X317 S.t4289 G.t317 D.t3894 S.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X318 D.t3893 G.t318 S.t4288 S.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X319 D.t3892 G.t319 S.t4287 S.t158 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X320 D.t3891 G.t320 S.t4286 S.t332 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X321 D.t3890 G.t321 S.t4285 S.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X322 D.t3889 G.t322 S.t4284 S.t270 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X323 D.t3888 G.t323 S.t4283 S.t321 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X324 S.t4282 G.t324 D.t3887 S.t216 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X325 D.t426 G.t325 S.t4281 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X326 D.t425 G.t326 S.t4280 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X327 D.t424 G.t327 S.t4279 S.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X328 D.t423 G.t328 S.t4278 S.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X329 S.t4277 G.t329 D.t422 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X330 S.t4276 G.t330 D.t421 S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X331 S.t4275 G.t331 D.t420 S.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X332 D.t419 G.t332 S.t4274 S.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X333 S.t4273 G.t333 D.t418 S.t406 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X334 D.t417 G.t334 S.t4272 S.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X335 D.t416 G.t335 S.t4271 S.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X336 S.t4270 G.t336 D.t415 S.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X337 D.t799 G.t337 S.t4269 S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X338 D.t798 G.t338 S.t4268 S.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X339 S.t4267 G.t339 D.t797 S.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X340 D.t796 G.t340 S.t4266 S.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X341 S.t4265 G.t341 D.t795 S.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X342 S.t4264 G.t342 D.t794 S.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X343 D.t793 G.t343 S.t4263 S.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X344 S.t4262 G.t344 D.t792 S.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X345 D.t791 G.t345 S.t4261 S.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X346 D.t790 G.t346 S.t4260 S.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X347 S.t4259 G.t347 D.t789 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X348 D.t788 G.t348 S.t4258 S.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X349 S.t4257 G.t349 D.t358 S.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X350 S.t4256 G.t350 D.t357 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X351 S.t4255 G.t351 D.t356 S.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X352 D.t355 G.t352 S.t4254 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X353 D.t354 G.t353 S.t4253 S.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X354 D.t353 G.t354 S.t4252 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X355 D.t352 G.t355 S.t4251 S.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X356 S.t4250 G.t356 D.t351 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X357 D.t350 G.t357 S.t4249 S.t176 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X358 S.t4248 G.t358 D.t349 S.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X359 D.t348 G.t359 S.t4247 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X360 D.t2562 G.t360 S.t4246 S.t216 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X361 S.t4245 G.t361 D.t2561 S.t332 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X362 D.t2560 G.t362 S.t4244 S.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X363 S.t4243 G.t363 D.t2559 S.t150 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X364 D.t2558 G.t364 S.t4242 S.t406 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X365 D.t2557 G.t365 S.t4241 S.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X366 D.t2556 G.t366 S.t4240 S.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X367 S.t4239 G.t367 D.t2555 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X368 S.t4238 G.t368 D.t2554 S.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X369 D.t2553 G.t369 S.t4237 S.t158 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X370 S.t4236 G.t370 D.t758 S.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X371 S.t4235 G.t371 D.t757 S.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X372 D.t756 G.t372 S.t4234 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X373 S.t4233 G.t373 D.t755 S.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X374 D.t754 G.t374 S.t4232 S.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X375 D.t753 G.t375 S.t4231 S.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X376 D.t752 G.t376 S.t4230 S.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X377 D.t751 G.t377 S.t4229 S.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X378 D.t750 G.t378 S.t4228 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X379 S.t4227 G.t379 D.t1045 S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X380 S.t4226 G.t380 D.t1044 S.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X381 D.t1043 G.t381 S.t4225 S.t270 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X382 D.t1042 G.t382 S.t4224 S.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X383 D.t1041 G.t383 S.t4223 S.t209 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X384 D.t1040 G.t384 S.t4222 S.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X385 S.t4221 G.t385 D.t1039 S.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X386 D.t1038 G.t386 S.t4220 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X387 S.t4219 G.t387 D.t3512 S.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X388 D.t3511 G.t388 S.t4218 S.t357 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X389 S.t4217 G.t389 D.t3510 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X390 S.t4216 G.t390 D.t3509 S.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X391 S.t4215 G.t391 D.t3352 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X392 S.t4214 G.t392 D.t3351 S.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X393 S.t4213 G.t393 D.t3350 S.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X394 D.t3349 G.t394 S.t4212 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X395 D.t3458 G.t395 S.t4211 S.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X396 D.t3457 G.t396 S.t4210 S.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X397 D.t3456 G.t397 S.t4209 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X398 S.t4208 G.t398 D.t3455 S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X399 D.t3495 G.t399 S.t4207 S.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X400 D.t3494 G.t400 S.t4206 S.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X401 D.t3493 G.t401 S.t4205 S.t218 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X402 D.t3492 G.t402 S.t4204 S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X403 D.t3232 G.t403 S.t4203 S.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X404 S.t4202 G.t404 D.t3231 S.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X405 D.t3230 G.t405 S.t4201 S.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X406 S.t4200 G.t406 D.t3229 S.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X407 D.t3356 G.t407 S.t4199 S.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X408 D.t3355 G.t408 S.t4198 S.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X409 S.t4197 G.t409 D.t3354 S.t139 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X410 D.t3353 G.t410 S.t4196 S.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X411 D.t3299 G.t411 S.t4195 S.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X412 S.t4194 G.t412 D.t3298 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X413 S.t4193 G.t413 D.t3297 S.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X414 S.t4192 G.t414 D.t3296 S.t357 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X415 D.t3788 G.t415 S.t4191 S.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X416 S.t4190 G.t416 D.t3787 S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X417 D.t3786 G.t417 S.t4189 S.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X418 S.t4188 G.t418 D.t3785 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X419 S.t4187 G.t419 D.t3762 S.t406 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X420 S.t4186 G.t420 D.t3761 S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X421 D.t3760 G.t421 S.t4185 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X422 S.t4184 G.t422 D.t3759 S.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X423 S.t4183 G.t423 D.t3792 S.t198 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X424 D.t3791 G.t424 S.t4182 S.t176 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X425 D.t3790 G.t425 S.t4181 S.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X426 D.t3789 G.t426 S.t4180 S.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X427 S.t4179 G.t427 D.t3967 S.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X428 D.t3966 G.t428 S.t4178 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X429 S.t4177 G.t429 D.t3965 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X430 S.t4176 G.t430 D.t3964 S.t332 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X431 S.t4175 G.t431 D.t1501 S.t406 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X432 S.t4174 G.t432 D.t1500 S.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X433 S.t4173 G.t433 D.t1499 S.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X434 D.t1498 G.t434 S.t4172 S.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X435 D.t3450 G.t435 S.t4171 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X436 D.t3449 G.t436 S.t4170 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X437 S.t4169 G.t437 D.t3448 S.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X438 D.t3447 G.t438 S.t4168 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X439 S.t4167 G.t439 D.t3643 S.t150 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X440 S.t4166 G.t440 D.t3642 S.t198 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X441 S.t4165 G.t441 D.t3641 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X442 D.t3640 G.t442 S.t4164 S.t176 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X443 S.t4163 G.t443 D.t3222 S.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X444 S.t4162 G.t444 D.t3221 S.t332 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X445 S.t4161 G.t445 D.t3220 S.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X446 D.t3219 G.t446 S.t4160 S.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X447 D.t3589 G.t447 S.t4159 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X448 S.t4158 G.t448 D.t3588 S.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X449 S.t4157 G.t449 D.t3587 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X450 S.t4156 G.t450 D.t3617 S.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X451 D.t3616 G.t451 S.t4155 S.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X452 S.t4154 G.t452 D.t3615 S.t443 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X453 D.t3536 G.t453 S.t4153 S.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X454 D.t3535 G.t454 S.t4152 S.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X455 S.t4151 G.t455 D.t3534 S.t270 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X456 D.t4113 G.t456 S.t4150 S.t158 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X457 S.t4149 G.t457 D.t4112 S.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X458 D.t4111 G.t458 S.t4148 S.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X459 S.t4147 G.t459 D.t3468 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X460 D.t3467 G.t460 S.t4146 S.t388 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X461 S.t4145 G.t461 D.t3466 S.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X462 D.t3744 G.t462 S.t4144 S.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X463 S.t4143 G.t463 D.t3743 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X464 S.t4142 G.t464 D.t3712 S.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X465 D.t3711 G.t465 S.t4141 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X466 S.t4140 G.t466 D.t4135 S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X467 S.t4139 G.t467 D.t4134 S.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X468 S.t4138 G.t468 D.t3486 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X469 S.t4137 G.t469 D.t3485 S.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X470 D.t3324 G.t470 S.t4136 S.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X471 D.t3323 G.t471 S.t4135 S.t357 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X472 S.t4134 G.t472 D.t4155 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X473 D.t4154 G.t473 S.t4133 S.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X474 S.t4132 G.t474 D.t3602 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X475 D.t3601 G.t475 S.t4131 S.t79 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X476 D.t3326 G.t476 S.t4130 S.t216 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X477 S.t4129 G.t477 D.t3325 S.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X478 D.t4099 G.t478 S.t4128 S.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X479 S.t4127 G.t479 D.t4098 S.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X480 D.t3902 G.t480 S.t4126 S.t270 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X481 D.t3901 G.t481 S.t4125 S.t321 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X482 D.t4115 G.t482 S.t4124 S.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X483 S.t4123 G.t483 D.t4114 S.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X484 D.t3446 G.t484 S.t4122 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X485 D.t3445 G.t485 S.t4121 S.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X486 S.t4120 G.t486 D.t3569 S.t216 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X487 S.t4119 G.t487 D.t3568 S.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X488 D.t4067 G.t488 S.t4118 S.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X489 S.t4117 G.t489 D.t4066 S.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X490 D.t3343 G.t490 S.t4116 S.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X491 D.t3342 G.t491 S.t4115 S.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X492 D.t4084 G.t492 S.t4114 S.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X493 D.t4083 G.t493 S.t4113 S.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X494 S.t4112 G.t494 D.t3596 S.t406 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X495 D.t3595 G.t495 S.t4111 S.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X496 S.t4110 G.t496 D.t3260 S.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X497 D.t3259 G.t497 S.t4109 S.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X498 D.t4096 G.t498 S.t4108 S.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X499 S.t4107 G.t499 D.t4095 S.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X500 S.t4106 G.t500 D.t4076 S.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X501 D.t4075 G.t501 S.t4105 S.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X502 D.t3565 G.t502 S.t4104 S.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X503 S.t4103 G.t503 D.t3564 S.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X504 S.t4102 G.t504 D.t3465 S.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X505 S.t4101 G.t505 D.t3464 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X506 D.t4400 G.t506 S.t4100 S.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X507 D.t4399 G.t507 S.t4099 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X508 S.t4098 G.t508 D.t3291 S.t270 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X509 D.t3290 G.t509 S.t4097 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X510 S.t4096 G.t510 D.t4103 S.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X511 S.t4095 G.t511 D.t4102 S.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X512 S.t4094 G.t512 D.t3856 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X513 D.t3855 G.t513 S.t4093 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X514 D.t3737 G.t514 S.t4092 S.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X515 D.t3736 G.t515 S.t4091 S.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X516 S.t4090 G.t516 D.t3331 S.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X517 D.t3330 G.t517 S.t4089 S.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X518 S.t4088 G.t518 D.t4101 S.t150 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X519 S.t4087 G.t519 D.t4100 S.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X520 S.t4086 G.t520 D.t3705 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X521 S.t4085 G.t521 D.t3704 S.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X522 S.t4084 G.t522 D.t3764 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X523 S.t4083 G.t523 D.t3763 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X524 D.t4304 G.t524 S.t4082 S.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X525 D.t4303 G.t525 S.t4081 S.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X526 S.t4080 G.t526 D.t4300 S.t357 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X527 D.t4299 G.t527 S.t4079 S.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X528 S.t4078 G.t528 D.t3767 S.t216 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X529 S.t4077 G.t529 D.t3766 S.t443 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X530 S.t4076 G.t530 D.t4210 S.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X531 D.t4209 G.t531 S.t4075 S.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X532 S.t4074 G.t532 D.t3963 S.t270 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X533 S.t4073 G.t533 D.t3962 S.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X534 S.t4072 G.t534 D.t4319 S.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X535 D.t4318 G.t535 S.t4071 S.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X536 D.t4263 G.t536 S.t4070 S.t357 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X537 S.t4069 G.t537 D.t4262 S.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X538 S.t4068 G.t538 D.t4223 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X539 D.t4222 G.t539 S.t4067 S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X540 S.t4066 G.t540 D.t4307 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X541 S.t4065 G.t541 D.t4306 S.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X542 S.t4064 G.t542 D.t4330 S.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X543 S.t4063 G.t543 D.t4329 S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X544 S.t4062 G.t544 D.t3169 S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X545 S.t4061 G.t545 D.t3168 S.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X546 S.t4060 G.t546 D.t3859 S.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X547 S.t4059 G.t547 D.t3858 S.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X548 D.t4081 G.t548 S.t4058 S.t216 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X549 S.t4057 G.t549 D.t4080 S.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X550 S.t4056 G.t550 D.t3441 S.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X551 D.t3440 G.t551 S.t4055 S.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X552 D.t3752 G.t552 S.t4054 S.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X553 S.t4053 G.t553 D.t3751 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X554 D.t4058 G.t554 S.t4052 S.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X555 S.t4051 G.t555 D.t4057 S.t139 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X556 D.t4120 G.t556 S.t4050 S.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X557 D.t4119 G.t557 S.t4049 S.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X558 S.t4048 G.t558 D.t3584 S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X559 D.t3583 G.t559 S.t4047 S.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X560 S.t4046 G.t560 D.t3322 S.t79 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X561 S.t4045 G.t561 D.t3321 S.t198 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X562 D.t3913 G.t562 S.t4044 S.t176 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X563 S.t4043 G.t563 D.t3912 S.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X564 S.t4042 G.t564 D.t4394 S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X565 S.t4041 G.t565 D.t3069 S.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X566 D.t3112 G.t566 S.t4040 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X567 D.t2821 G.t567 S.t4039 S.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X568 S.t4038 G.t568 D.t4409 S.t332 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X569 S.t4037 G.t569 D.t2728 S.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X570 S.t4036 G.t570 D.t1313 S.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X571 S.t4035 G.t571 D.t3843 S.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X572 S.t4034 G.t572 D.t3808 S.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X573 D.t3626 G.t573 S.t4033 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X574 S.t4032 G.t574 D.t2995 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X575 S.t4031 G.t575 D.t4157 S.t198 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X576 S.t4030 G.t576 D.t3333 S.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X577 S.t4029 G.t577 D.t4437 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X578 D.t3657 G.t578 S.t4028 S.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X579 S.t4027 G.t579 D.t3773 S.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X580 D.t3916 G.t580 S.t4026 S.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X581 D.t141 G.t581 S.t4025 S.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X582 D.t3605 G.t582 S.t4024 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X583 S.t4023 G.t583 D.t3854 S.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X584 S.t4022 G.t584 D.t3932 S.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X585 S.t4021 G.t585 D.t4130 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X586 S.t4020 G.t586 D.t3638 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X587 D.t4097 G.t587 S.t4019 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X588 D.t4091 G.t588 S.t4018 S.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X589 D.t3289 G.t589 S.t4017 S.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X590 S.t4016 G.t590 D.t3635 S.t443 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X591 S.t4015 G.t591 D.t3707 S.t270 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X592 S.t4014 G.t592 D.t3907 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X593 D.t4093 G.t593 S.t4013 S.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X594 S.t4012 G.t594 D.t4124 S.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X595 D.t3571 G.t595 S.t4011 S.t388 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X596 D.t3285 G.t596 S.t4010 S.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X597 S.t4009 G.t597 D.t3245 S.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X598 S.t4008 G.t598 D.t3634 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X599 D.t3319 G.t599 S.t4007 S.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X600 S.t4006 G.t600 D.t3316 S.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X601 D.t3329 G.t601 S.t4005 S.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X602 S.t4004 G.t602 D.t4122 S.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X603 D.t4446 G.t603 S.t4003 S.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X604 S.t4002 G.t604 D.t3443 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X605 D.t3985 G.t605 S.t4001 S.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X606 S.t4000 G.t606 D.t3706 S.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X607 S.t3999 G.t607 D.t4090 S.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X608 D.t4138 G.t608 S.t3998 S.t216 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X609 S.t3997 G.t609 D.t4450 S.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X610 S.t3996 G.t610 D.t3851 S.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X611 S.t3995 G.t611 D.t3604 S.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X612 D.t4077 G.t612 S.t3994 S.t321 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X613 S.t3993 G.t613 D.t3739 S.t216 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X614 D.t4432 G.t614 S.t3992 S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X615 S.t3991 G.t615 D.t4285 S.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X616 D.t3972 G.t616 S.t3990 S.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X617 S.t3989 G.t617 D.t4385 S.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X618 S.t3988 G.t618 D.t4440 S.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X619 D.t4406 G.t619 S.t3987 S.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X620 D.t4182 G.t620 S.t3986 S.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X621 D.t4055 G.t621 S.t3985 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X622 D.t3532 G.t622 S.t3984 S.t150 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X623 S.t3983 G.t623 D.t4429 S.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X624 D.t3421 G.t624 S.t3982 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X625 S.t3981 G.t625 D.t4455 S.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X626 D.t4435 G.t626 S.t3980 S.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X627 S.t3979 G.t627 D.t4360 S.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X628 D.t3235 G.t628 S.t3978 S.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X629 S.t3977 G.t629 D.t3244 S.t79 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X630 D.t4397 G.t630 S.t3976 S.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X631 S.t3975 G.t631 D.t3800 S.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X632 D.t4320 G.t632 S.t3974 S.t538 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X633 S.t3973 G.t633 D.t4248 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X634 S.t3972 G.t634 D.t4217 S.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X635 S.t3971 G.t635 D.t4220 S.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X636 D.t4189 G.t636 S.t3970 S.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X637 D.t4177 G.t637 S.t3969 S.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X638 S.t3968 G.t638 D.t4380 S.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X639 D.t4310 G.t639 S.t3967 S.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X640 S.t3966 G.t640 D.t3852 S.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X641 D.t4284 G.t641 S.t3965 S.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X642 S.t3964 G.t642 D.t3579 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X643 S.t3963 G.t643 D.t4290 S.t231 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X644 D.t4180 G.t644 S.t3962 S.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X645 D.t4188 G.t645 S.t3961 S.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X646 S.t3960 G.t646 D.t4213 S.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X647 S.t3959 G.t647 D.t4270 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X648 S.t3958 G.t648 D.t4271 S.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X649 S.t3957 G.t649 D.t4339 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X650 D.t4305 G.t650 S.t3956 S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X651 S.t3955 G.t651 D.t4275 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X652 S.t3954 G.t652 D.t4276 S.t357 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X653 S.t3953 G.t653 D.t4281 S.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X654 S.t3952 G.t654 D.t4322 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X655 D.t4321 G.t655 S.t3951 S.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X656 S.t3950 G.t656 D.t4245 S.t216 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X657 S.t3949 G.t657 D.t4252 S.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X658 S.t3948 G.t658 D.t4312 S.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X659 S.t3947 G.t659 D.t4298 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X660 D.t4324 G.t660 S.t3946 S.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X661 S.t3945 G.t661 D.t4362 S.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X662 D.t4219 G.t662 S.t3944 S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X663 S.t3943 G.t663 D.t4247 S.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X664 D.t4162 G.t664 S.t3942 S.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X665 S.t3941 G.t665 D.t4206 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X666 S.t3940 G.t666 D.t4216 S.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X667 S.t3939 G.t667 D.t4185 S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X668 D.t4181 G.t668 S.t3938 S.t538 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X669 D.t4175 G.t669 S.t3937 S.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X670 D.t3578 G.t670 S.t3936 S.t443 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X671 D.t3933 G.t671 S.t3935 S.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X672 D.t3774 G.t672 S.t3934 S.t158 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X673 S.t3933 G.t673 D.t3755 S.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X674 S.t3932 G.t674 D.t3812 S.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X675 D.t3658 G.t675 S.t3931 S.t183 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X676 D.t3659 G.t676 S.t3930 S.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X677 S.t3929 G.t677 D.t4121 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X678 S.t3928 G.t678 D.t3582 S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X679 D.t3320 G.t679 S.t3927 S.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X680 D.t3624 G.t680 S.t3926 S.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X681 D.t2709 G.t681 S.t3925 S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X682 S.t3924 G.t682 D.t4110 S.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X683 D.t157 G.t683 S.t3923 S.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X684 D.t4414 G.t684 S.t3922 S.t216 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X685 D.t3344 G.t685 S.t3921 S.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X686 D.t4390 G.t686 S.t3920 S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X687 D.t2926 G.t687 S.t3919 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X688 D.t4402 G.t688 S.t3918 S.t231 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X689 D.t4343 G.t689 S.t3917 S.t150 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X690 D.t2911 G.t690 S.t3916 S.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X691 S.t3915 G.t691 D.t3163 S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X692 D.t2932 G.t692 S.t3914 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X693 S.t3913 G.t693 D.t2773 S.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X694 S.t3912 G.t694 D.t3067 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X695 S.t3911 G.t695 D.t2877 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X696 D.t3026 G.t696 S.t3910 S.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X697 S.t3909 G.t697 D.t3017 S.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X698 D.t2976 G.t698 S.t3908 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X699 S.t3907 G.t699 D.t2867 S.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X700 D.t2833 G.t700 S.t3906 S.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X701 S.t3905 G.t701 D.t3081 S.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X702 S.t3904 G.t702 D.t2972 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X703 D.t3028 G.t703 S.t3903 S.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X704 D.t2880 G.t704 S.t3902 S.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X705 D.t3099 G.t705 S.t3901 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X706 S.t3900 G.t706 D.t3159 S.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X707 S.t3899 G.t707 D.t2896 S.t231 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X708 D.t2984 G.t708 S.t3898 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X709 D.t3022 G.t709 S.t3897 S.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X710 D.t2801 G.t710 S.t3896 S.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X711 S.t3895 G.t711 D.t2930 S.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X712 D.t2922 G.t712 S.t3894 S.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X713 S.t3893 G.t713 D.t3107 S.t218 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X714 D.t2830 G.t714 S.t3892 S.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X715 S.t3891 G.t715 D.t3075 S.t388 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X716 S.t3890 G.t716 D.t3070 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X717 S.t3889 G.t717 D.t3043 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X718 S.t3888 G.t718 D.t2858 S.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X719 D.t2834 G.t719 S.t3887 S.t406 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X720 D.t2963 G.t720 S.t3886 S.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X721 S.t3885 G.t721 D.t2954 S.t183 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X722 S.t3884 G.t722 D.t2902 S.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X723 D.t2875 G.t723 S.t3883 S.t538 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X724 D.t2818 G.t724 S.t3882 S.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X725 D.t2802 G.t725 S.t3881 S.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X726 S.t3880 G.t726 D.t3104 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X727 D.t3024 G.t727 S.t3879 S.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X728 D.t3130 G.t728 S.t3878 S.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X729 S.t3877 G.t729 D.t3033 S.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X730 D.t3077 G.t730 S.t3876 S.t79 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X731 S.t3875 G.t731 D.t2999 S.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X732 S.t3874 G.t732 D.t3098 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X733 S.t3873 G.t733 D.t2933 S.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X734 S.t3872 G.t734 D.t2958 S.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X735 S.t3871 G.t735 D.t2947 S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X736 S.t3870 G.t736 D.t2881 S.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X737 D.t2860 G.t737 S.t3869 S.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X738 D.t2789 G.t738 S.t3868 S.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X739 D.t2771 G.t739 S.t3867 S.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X740 S.t3866 G.t740 D.t2927 S.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X741 D.t2913 G.t741 S.t3865 S.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X742 D.t4407 G.t742 S.t3864 S.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X743 S.t3863 G.t743 D.t2979 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X744 D.t3006 G.t744 S.t3862 S.t183 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X745 D.t4388 G.t745 S.t3861 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X746 D.t4401 G.t746 S.t3860 S.t150 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X747 D.t3116 G.t747 S.t3859 S.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X748 D.t3012 G.t748 S.t3858 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X749 D.t3014 G.t749 S.t3857 S.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X750 D.t3076 G.t750 S.t3856 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X751 D.t2907 G.t751 S.t3855 S.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X752 S.t3854 G.t752 D.t4337 S.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X753 D.t3555 G.t753 S.t3853 S.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X754 D.t2892 G.t754 S.t3852 S.t357 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X755 D.t140 G.t755 S.t3851 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X756 D.t4443 G.t756 S.t3850 S.t538 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X757 S.t3849 G.t757 D.t3710 S.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X758 S.t3848 G.t758 D.t3427 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X759 D.t4448 G.t759 S.t3847 S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X760 S.t3846 G.t760 D.t4211 S.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X761 S.t3845 G.t761 D.t3332 S.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X762 S.t3844 G.t762 D.t4089 S.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X763 D.t4137 G.t763 S.t3843 S.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X764 S.t3842 G.t764 D.t3470 S.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X765 S.t3841 G.t765 D.t3748 S.t231 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X766 D.t3254 G.t766 S.t3840 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X767 S.t3839 G.t767 D.t3709 S.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X768 D.t4117 G.t768 S.t3838 S.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X769 S.t3837 G.t769 D.t3977 S.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X770 D.t4456 G.t770 S.t3836 S.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X771 S.t3835 G.t771 D.t4104 S.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X772 D.t3292 G.t772 S.t3834 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X773 S.t3833 G.t773 D.t3508 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X774 S.t3832 G.t774 D.t3567 S.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X775 D.t103 G.t775 S.t3831 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X776 S.t3830 G.t776 D.t3021 S.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X777 S.t3829 G.t777 D.t4426 S.t357 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X778 S.t3828 G.t778 D.t3429 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X779 D.t4107 G.t779 S.t3827 S.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X780 D.t3740 G.t780 S.t3826 S.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X781 S.t3825 G.t781 D.t3869 S.t216 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X782 D.t3769 G.t782 S.t3824 S.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X783 S.t3823 G.t783 D.t4131 S.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X784 S.t3822 G.t784 D.t3725 S.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X785 D.t3772 G.t785 S.t3821 S.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X786 D.t3713 G.t786 S.t3820 S.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X787 D.t4404 G.t787 S.t3819 S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X788 S.t3818 G.t788 D.t4129 S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X789 D.t3572 G.t789 S.t3817 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X790 S.t3816 G.t790 D.t3537 S.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X791 D.t4158 G.t791 S.t3815 S.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X792 S.t3814 G.t792 D.t2838 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X793 S.t3813 G.t793 D.t4371 S.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X794 S.t3812 G.t794 D.t3531 S.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X795 D.t3914 G.t795 S.t3811 S.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X796 D.t4379 G.t796 S.t3810 S.t538 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X797 S.t3809 G.t797 D.t3853 S.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X798 D.t3433 G.t798 S.t3808 S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X799 D.t3328 G.t799 S.t3807 S.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X800 S.t3806 G.t800 D.t3444 S.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X801 D.t3866 G.t801 S.t3805 S.t443 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X802 S.t3804 G.t802 D.t4161 S.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X803 D.t4128 G.t803 S.t3803 S.t183 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X804 S.t3802 G.t804 D.t4327 S.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X805 S.t3801 G.t805 D.t4460 S.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X806 S.t3800 G.t806 D.t4444 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X807 D.t3453 G.t807 S.t3799 S.t139 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X808 S.t3798 G.t808 D.t3585 S.t158 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X809 D.t3867 G.t809 S.t3797 S.t209 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X810 S.t3796 G.t810 D.t4358 S.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X811 S.t3795 G.t811 D.t3654 S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X812 D.t3284 G.t812 S.t3794 S.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X813 S.t3793 G.t813 D.t3915 S.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X814 D.t3708 G.t814 S.t3792 S.t332 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X815 D.t4125 G.t815 S.t3791 S.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X816 S.t3790 G.t816 D.t3768 S.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X817 D.t4374 G.t817 S.t3789 S.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X818 D.t3653 G.t818 S.t3788 S.t231 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X819 D.t4160 G.t819 S.t3787 S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X820 S.t3786 G.t820 D.t3879 S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X821 D.t3652 G.t821 S.t3785 S.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X822 S.t3784 G.t822 D.t3586 S.t321 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X823 D.t4408 G.t823 S.t3783 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X824 S.t3782 G.t824 D.t3327 S.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X825 D.t3530 G.t825 S.t3781 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X826 D.t4436 G.t826 S.t3780 S.t357 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X827 S.t3779 G.t827 D.t4412 S.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X828 S.t3778 G.t828 D.t4215 S.t388 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X829 D.t3496 G.t829 S.t3777 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X830 D.t4045 G.t830 S.t3776 S.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X831 S.t3775 G.t831 D.t3504 S.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X832 D.t3825 G.t832 S.t3774 S.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X833 S.t3773 G.t833 D.t3317 S.t209 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X834 S.t3772 G.t834 D.t3246 S.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X835 D.t4457 G.t835 S.t3771 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X836 S.t3770 G.t836 D.t3594 S.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X837 D.t4288 G.t837 S.t3769 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X838 S.t3768 G.t838 D.t3563 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X839 D.t4441 G.t839 S.t3767 S.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X840 D.t4428 G.t840 S.t3766 S.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X841 S.t3765 G.t841 D.t4054 S.t231 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X842 D.t3606 G.t842 S.t3764 S.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X843 S.t3763 G.t843 D.t3283 S.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X844 D.t3505 G.t844 S.t3762 S.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X845 D.t3905 G.t845 S.t3761 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X846 D.t4421 G.t846 S.t3760 S.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X847 D.t3281 G.t847 S.t3759 S.t443 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X848 S.t3758 G.t848 D.t3703 S.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X849 D.t4078 G.t849 S.t3757 S.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X850 D.t4116 G.t850 S.t3756 S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X851 S.t3755 G.t851 D.t4143 S.t218 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X852 S.t3754 G.t852 D.t2962 S.t388 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X853 D.t4422 G.t853 S.t3753 S.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X854 D.t4346 G.t854 S.t3752 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X855 S.t3751 G.t855 D.t4424 S.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X856 S.t3750 G.t856 D.t4198 S.t321 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X857 D.t3502 G.t857 S.t3749 S.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X858 S.t3748 G.t858 D.t3451 S.t183 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X859 D.t3422 G.t859 S.t3747 S.t406 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X860 S.t3746 G.t860 D.t3428 S.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X861 S.t3745 G.t861 D.t4454 S.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X862 D.t4425 G.t862 S.t3744 S.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X863 S.t3743 G.t863 D.t4419 S.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X864 D.t4416 G.t864 S.t3742 S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X865 S.t3741 G.t865 D.t4405 S.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X866 D.t4186 G.t866 S.t3740 S.t79 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X867 S.t3739 G.t867 D.t3603 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X868 D.t4348 G.t868 S.t3738 S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X869 S.t3737 G.t869 D.t3688 S.t176 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X870 D.t4118 G.t870 S.t3736 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X871 S.t3735 G.t871 D.t4289 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X872 S.t3734 G.t872 D.t4184 S.t321 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X873 S.t3733 G.t873 D.t3282 S.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X874 S.t3732 G.t874 D.t3655 S.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X875 D.t3656 G.t875 S.t3731 S.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X876 D.t4453 G.t876 S.t3730 S.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X877 D.t4445 G.t877 S.t3729 S.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X878 S.t3728 G.t878 D.t4439 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X879 S.t3727 G.t879 D.t4442 S.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X880 S.t3726 G.t880 D.t4438 S.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X881 S.t3725 G.t881 D.t4434 S.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X882 D.t4431 G.t882 S.t3724 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X883 S.t3723 G.t883 D.t4403 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X884 D.t4393 G.t884 S.t3722 S.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X885 D.t4359 G.t885 S.t3721 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X886 S.t3720 G.t886 D.t4375 S.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X887 D.t4153 G.t887 S.t3719 S.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X888 S.t3718 G.t888 D.t3463 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X889 D.t3503 G.t889 S.t3717 S.t332 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X890 S.t3716 G.t890 D.t4254 S.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X891 S.t3715 G.t891 D.t4178 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X892 D.t4123 G.t892 S.t3714 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X893 D.t4433 G.t893 S.t3713 S.t357 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X894 S.t3712 G.t894 D.t4423 S.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X895 D.t4415 G.t895 S.t3711 S.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X896 S.t3710 G.t896 D.t4351 S.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X897 S.t3709 G.t897 D.t4345 S.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X898 S.t3708 G.t898 D.t4250 S.t321 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X899 S.t3707 G.t899 D.t3276 S.t388 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X900 D.t3275 G.t900 S.t3706 S.t538 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X901 S.t3705 G.t901 D.t3947 S.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X902 S.t3704 G.t902 D.t3765 S.t209 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X903 D.t3454 G.t903 S.t3703 S.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X904 S.t3702 G.t904 D.t4212 S.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X905 S.t3701 G.t905 D.t4342 S.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X906 D.t4336 G.t906 S.t3700 S.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X907 S.t3699 G.t907 D.t4382 S.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X908 D.t4283 G.t908 S.t3698 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X909 D.t3452 G.t909 S.t3697 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X910 S.t3696 G.t910 D.t3233 S.t231 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X911 D.t3318 G.t911 S.t3695 S.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X912 D.t4228 G.t912 S.t3694 S.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X913 S.t3693 G.t913 D.t4381 S.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X914 S.t3692 G.t914 D.t4378 S.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X915 D.t4243 G.t915 S.t3691 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X916 S.t3690 G.t916 D.t4176 S.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X917 S.t3689 G.t917 D.t4376 S.t538 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X918 D.t4364 G.t918 S.t3688 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X919 D.t3234 G.t919 S.t3687 S.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X920 D.t4258 G.t920 S.t3686 S.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X921 S.t3685 G.t921 D.t4056 S.t443 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X922 D.t3689 G.t922 S.t3684 S.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X923 D.t4152 G.t923 S.t3683 S.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X924 D.t4315 G.t924 S.t3682 S.t443 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X925 S.t3681 G.t925 D.t4297 S.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X926 D.t4277 G.t926 S.t3680 S.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X927 D.t4230 G.t927 S.t3679 S.t158 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X928 S.t3678 G.t928 D.t4383 S.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X929 S.t3677 G.t929 D.t4183 S.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X930 S.t3676 G.t930 D.t4065 S.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X931 S.t3675 G.t931 D.t4377 S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X932 D.t4365 G.t932 S.t3674 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X933 S.t3673 G.t933 D.t4373 S.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X934 D.t4372 G.t934 S.t3672 S.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X935 D.t4159 G.t935 S.t3671 S.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X936 S.t3670 G.t936 D.t4331 S.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X937 S.t3669 G.t937 D.t3738 S.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X938 S.t3668 G.t938 D.t4253 S.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X939 D.t4308 G.t939 S.t3667 S.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X940 S.t3666 G.t940 D.t4309 S.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X941 D.t4317 G.t941 S.t3665 S.t198 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X942 S.t3664 G.t942 D.t4396 S.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X943 S.t3663 G.t943 D.t4413 S.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X944 D.t4452 G.t944 S.t3662 S.t443 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X945 S.t3661 G.t945 D.t4449 S.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X946 S.t3660 G.t946 D.t4420 S.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X947 D.t4417 G.t947 S.t3659 S.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X948 D.t4341 G.t948 S.t3658 S.t270 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X949 D.t4278 G.t949 S.t3657 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X950 S.t3656 G.t950 D.t4287 S.t538 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X951 D.t4294 G.t951 S.t3655 S.t388 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X952 S.t3654 G.t952 D.t4295 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X953 D.t4313 G.t953 S.t3653 S.t139 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X954 S.t3652 G.t954 D.t4311 S.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X955 D.t4316 G.t955 S.t3651 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X956 D.t4350 G.t956 S.t3650 S.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X957 S.t3649 G.t957 D.t4314 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X958 D.t4227 G.t958 S.t3648 S.t332 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X959 S.t3647 G.t959 D.t4249 S.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X960 S.t3646 G.t960 D.t4268 S.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X961 D.t4280 G.t961 S.t3645 S.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X962 D.t4352 G.t962 S.t3644 S.t231 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X963 S.t3643 G.t963 D.t4302 S.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X964 D.t4301 G.t964 S.t3642 S.t406 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X965 S.t3641 G.t965 D.t4323 S.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X966 D.t4325 G.t966 S.t3640 S.t231 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X967 S.t3639 G.t967 D.t4326 S.t321 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X968 S.t3638 G.t968 D.t4363 S.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X969 S.t3637 G.t969 D.t4361 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X970 S.t3636 G.t970 D.t4366 S.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X971 D.t4369 G.t971 S.t3635 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X972 D.t4367 G.t972 S.t3634 S.t218 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X973 D.t4368 G.t973 S.t3633 S.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X974 S.t3632 G.t974 D.t4370 S.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X975 S.t3631 G.t975 D.t4357 S.t388 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X976 S.t3630 G.t976 D.t4349 S.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X977 S.t3629 G.t977 D.t4286 S.t406 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X978 D.t4273 G.t978 S.t3628 S.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X979 S.t3627 G.t979 D.t4251 S.t209 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X980 S.t3626 G.t980 D.t4179 S.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X981 D.t4194 G.t981 S.t3625 S.t139 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X982 S.t3624 G.t982 D.t4214 S.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X983 S.t3623 G.t983 D.t4231 S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X984 D.t4241 G.t984 S.t3622 S.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X985 S.t3621 G.t985 D.t4244 S.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X986 D.t4257 G.t986 S.t3620 S.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X987 S.t3619 G.t987 D.t4296 S.t231 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X988 D.t4282 G.t988 S.t3618 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X989 S.t3617 G.t989 D.t4279 S.t198 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X990 D.t4272 G.t990 S.t3616 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X991 S.t3615 G.t991 D.t4291 S.t198 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X992 S.t3614 G.t992 D.t4292 S.t538 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X993 D.t4269 G.t993 S.t3613 S.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X994 D.t4274 G.t994 S.t3612 S.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X995 S.t3611 G.t995 D.t4265 S.t443 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X996 S.t3610 G.t996 D.t4061 S.t218 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X997 D.t4236 G.t997 S.t3609 S.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X998 S.t3608 G.t998 D.t4208 S.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X999 D.t4256 G.t999 S.t3607 S.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1000 S.t3606 G.t1000 D.t4246 S.t388 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1001 D.t4261 G.t1001 S.t3605 S.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1002 D.t4255 G.t1002 S.t3604 S.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1003 D.t4259 G.t1003 S.t3603 S.t406 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1004 S.t3602 G.t1004 D.t4260 S.t183 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1005 S.t3601 G.t1005 D.t4264 S.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1006 S.t3600 G.t1006 D.t4266 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1007 S.t3599 G.t1007 D.t4267 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1008 D.t4233 G.t1008 S.t3598 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1009 D.t4226 G.t1009 S.t3597 S.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1010 S.t3596 G.t1010 D.t4192 S.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1011 S.t3595 G.t1011 D.t4187 S.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1012 S.t3594 G.t1012 D.t4064 S.t332 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1013 D.t4193 G.t1013 S.t3593 S.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1014 S.t3592 G.t1014 D.t4203 S.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1015 S.t3591 G.t1015 D.t4239 S.t357 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1016 D.t4224 G.t1016 S.t3590 S.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1017 S.t3589 G.t1017 D.t4218 S.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1018 S.t3588 G.t1018 D.t4225 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1019 D.t4229 G.t1019 S.t3587 S.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1020 S.t3586 G.t1020 D.t4232 S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1021 D.t4234 G.t1021 S.t3585 S.t198 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1022 S.t3584 G.t1022 D.t4235 S.t176 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1023 D.t4237 G.t1023 S.t3583 S.t139 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1024 S.t3582 G.t1024 D.t4238 S.t538 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1025 D.t4240 G.t1025 S.t3581 S.t270 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1026 D.t4196 G.t1026 S.t3580 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1027 D.t4200 G.t1027 S.t3579 S.t321 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1028 S.t3578 G.t1028 D.t4190 S.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1029 S.t3577 G.t1029 D.t4191 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1030 D.t4195 G.t1030 S.t3576 S.t183 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1031 S.t3575 G.t1031 D.t4197 S.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1032 D.t4199 G.t1032 S.t3574 S.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1033 S.t3573 G.t1033 D.t4201 S.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1034 D.t4202 G.t1034 S.t3572 S.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1035 S.t3571 G.t1035 D.t4204 S.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1036 D.t4205 G.t1036 S.t3570 S.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1037 D.t4207 G.t1037 S.t3569 S.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1038 S.t3568 G.t1038 D.t2378 S.t150 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1039 D.t2447 G.t1039 S.t3567 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1040 S.t3566 G.t1040 D.t2444 S.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1041 S.t3565 G.t1041 D.t2427 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1042 D.t2399 G.t1042 S.t3564 S.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1043 S.t3563 G.t1043 D.t990 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1044 D.t3438 G.t1044 S.t3562 S.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1045 S.t3561 G.t1045 D.t1221 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1046 D.t2358 G.t1046 S.t3560 S.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1047 S.t3559 G.t1047 D.t2303 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1048 D.t2408 G.t1048 S.t3558 S.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1049 S.t3557 G.t1049 D.t2373 S.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1050 S.t3556 G.t1050 D.t2223 S.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1051 S.t3555 G.t1051 D.t2230 S.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1052 S.t3554 G.t1052 D.t2242 S.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1053 D.t2265 G.t1053 S.t3553 S.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1054 S.t3552 G.t1054 D.t3908 S.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1055 D.t4092 G.t1055 S.t3551 S.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1056 D.t4127 G.t1056 S.t3550 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1057 S.t3549 G.t1057 D.t3857 S.t443 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1058 S.t3548 G.t1058 D.t3952 S.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1059 D.t3533 G.t1059 S.t3547 S.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1060 D.t3469 G.t1060 S.t3546 S.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1061 S.t3545 G.t1061 D.t3286 S.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1062 S.t3544 G.t1062 D.t3714 S.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1063 D.t3507 G.t1063 S.t3543 S.t218 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1064 D.t3476 G.t1064 S.t3542 S.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1065 S.t3541 G.t1065 D.t3690 S.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1066 D.t3413 G.t1066 S.t3540 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1067 S.t3539 G.t1067 D.t3934 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1068 S.t3538 G.t1068 D.t3694 S.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1069 D.t3775 G.t1069 S.t3537 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1070 S.t3536 G.t1070 D.t3754 S.t406 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1071 S.t3535 G.t1071 D.t3776 S.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1072 D.t3519 G.t1072 S.t3534 S.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1073 D.t3821 G.t1073 S.t3533 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1074 S.t3532 G.t1074 D.t3801 S.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1075 D.t3874 G.t1075 S.t3531 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1076 S.t3530 G.t1076 D.t4068 S.t538 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1077 D.t3742 G.t1077 S.t3529 S.t139 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1078 S.t3528 G.t1078 D.t4074 S.t443 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1079 D.t3566 G.t1079 S.t3527 S.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1080 D.t3560 G.t1080 S.t3526 S.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1081 D.t3561 G.t1081 S.t3525 S.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1082 D.t3619 G.t1082 S.t3524 S.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1083 D.t3581 G.t1083 S.t3523 S.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1084 S.t3522 G.t1084 D.t3618 S.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1085 D.t3580 G.t1085 S.t3521 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1086 D.t3430 G.t1086 S.t3520 S.t216 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1087 D.t3431 G.t1087 S.t3519 S.t321 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1088 D.t4087 G.t1088 S.t3518 S.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1089 D.t4088 G.t1089 S.t3517 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1090 D.t4044 G.t1090 S.t3516 S.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1091 S.t3515 G.t1091 D.t4086 S.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1092 S.t3514 G.t1092 D.t4043 S.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1093 D.t4085 G.t1093 S.t3513 S.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1094 S.t3512 G.t1094 D.t3265 S.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1095 D.t3266 G.t1095 S.t3511 S.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1096 S.t3510 G.t1096 D.t3796 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1097 S.t3509 G.t1097 D.t3797 S.t406 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1098 D.t3910 G.t1098 S.t3508 S.t198 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1099 S.t3507 G.t1099 D.t3909 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1100 S.t3506 G.t1100 D.t3042 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1101 S.t3505 G.t1101 D.t3160 S.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1102 D.t2827 G.t1102 S.t3504 S.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1103 S.t3503 G.t1103 D.t3746 S.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1104 D.t4451 G.t1104 S.t3502 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1105 S.t3501 G.t1105 D.t2824 S.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1106 D.t3145 G.t1106 S.t3500 S.t183 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1107 D.t4447 G.t1107 S.t3499 S.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1108 S.t3498 G.t1108 D.t1094 S.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1109 D.t2909 G.t1109 S.t3497 S.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1110 S.t3496 G.t1110 D.t4430 S.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1111 D.t2848 G.t1111 S.t3495 S.t388 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1112 S.t3494 G.t1112 D.t3147 S.t538 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1113 D.t2961 G.t1113 S.t3493 S.t270 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1114 S.t3492 G.t1114 D.t4458 S.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1115 D.t4459 G.t1115 S.t3491 S.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1116 D.t2825 G.t1116 S.t3490 S.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1117 D.t3111 G.t1117 S.t3489 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1118 D.t2810 G.t1118 S.t3488 S.t209 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1119 S.t3487 G.t1119 D.t2793 S.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1120 S.t3486 G.t1120 D.t589 S.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1121 S.t3485 G.t1121 D.t2732 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1122 D.t4221 G.t1122 S.t3484 S.t231 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1123 S.t3483 G.t1123 D.t2692 S.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1124 S.t3482 G.t1124 D.t2712 S.t150 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1125 S.t3481 G.t1125 D.t1358 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1126 S.t3480 G.t1126 D.t504 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1127 D.t1674 G.t1127 S.t3479 S.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1128 S.t3478 G.t1128 D.t1570 S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1129 S.t3477 G.t1129 D.t3166 S.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1130 S.t3476 G.t1130 D.t3960 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1131 D.t3692 G.t1131 S.t3475 S.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1132 S.t3474 G.t1132 D.t3264 S.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1133 D.t3518 G.t1133 S.t3473 S.t218 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1134 D.t3727 G.t1134 S.t3472 S.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1135 S.t3471 G.t1135 D.t3521 S.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1136 D.t3838 G.t1136 S.t3470 S.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1137 S.t3469 G.t1137 D.t3523 S.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1138 D.t3700 G.t1138 S.t3468 S.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1139 D.t2675 G.t1139 S.t3467 S.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1140 D.t3187 G.t1140 S.t3466 S.t139 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1141 S.t3465 G.t1141 D.t117 S.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1142 S.t3464 G.t1142 D.t84 S.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1143 D.t76 G.t1143 S.t3463 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1144 D.t72 G.t1144 S.t3462 S.t357 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1145 S.t3461 G.t1145 D.t3183 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1146 S.t3460 G.t1146 D.t1 S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1147 S.t3459 G.t1147 D.t4356 S.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1148 S.t3458 G.t1148 D.t3172 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1149 D.t79 G.t1149 S.t3457 S.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1150 S.t3456 G.t1150 D.t2087 S.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1151 D.t4166 G.t1151 S.t3455 S.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1152 S.t3454 G.t1152 D.t4418 S.t198 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1153 D.t2611 G.t1153 S.t3453 S.t176 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1154 D.t2637 G.t1154 S.t3452 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1155 D.t2655 G.t1155 S.t3451 S.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1156 D.t2613 G.t1156 S.t3450 S.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1157 S.t3449 G.t1157 D.t2643 S.t183 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1158 D.t2660 G.t1158 S.t3448 S.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1159 D.t4427 G.t1159 S.t3447 S.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1160 D.t2624 G.t1160 S.t3446 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1161 D.t4332 G.t1161 S.t3445 S.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1162 D.t4353 G.t1162 S.t3444 S.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1163 S.t3443 G.t1163 D.t4354 S.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1164 S.t3442 G.t1164 D.t2698 S.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1165 D.t3174 G.t1165 S.t3441 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1166 D.t4168 G.t1166 S.t3440 S.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1167 S.t3439 G.t1167 D.t4242 S.t139 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1168 S.t3438 G.t1168 D.t2711 S.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1169 D.t2716 G.t1169 S.t3437 S.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1170 D.t4171 G.t1170 S.t3436 S.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1171 S.t3435 G.t1171 D.t4167 S.t332 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1172 D.t2714 G.t1172 S.t3434 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1173 D.t4172 G.t1173 S.t3433 S.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1174 S.t3432 G.t1174 D.t3108 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1175 S.t3431 G.t1175 D.t4170 S.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1176 S.t3430 G.t1176 D.t4165 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1177 S.t3429 G.t1177 D.t4173 S.t176 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1178 D.t2731 G.t1178 S.t3428 S.t321 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1179 D.t2836 G.t1179 S.t3427 S.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1180 D.t3173 G.t1180 S.t3426 S.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1181 D.t3170 G.t1181 S.t3425 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1182 D.t4174 G.t1182 S.t3424 S.t183 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1183 D.t2339 G.t1183 S.t3423 S.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1184 D.t2619 G.t1184 S.t3422 S.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1185 D.t2676 G.t1185 S.t3421 S.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1186 S.t3420 G.t1186 D.t3176 S.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1187 D.t2603 G.t1187 S.t3419 S.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1188 D.t2654 G.t1188 S.t3418 S.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1189 S.t3417 G.t1189 D.t2632 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1190 D.t2657 G.t1190 S.t3416 S.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1191 D.t2212 G.t1191 S.t3415 S.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1192 D.t2661 G.t1192 S.t3414 S.t209 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1193 S.t3413 G.t1193 D.t1717 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1194 S.t3412 G.t1194 D.t4169 S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1195 S.t3411 G.t1195 D.t2336 S.t139 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1196 S.t3410 G.t1196 D.t2599 S.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1197 D.t2629 G.t1197 S.t3409 S.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1198 S.t3408 G.t1198 D.t2680 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1199 D.t3970 G.t1199 S.t3407 S.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1200 D.t3570 G.t1200 S.t3406 S.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1201 S.t3405 G.t1201 D.t3980 S.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1202 D.t3432 G.t1202 S.t3404 S.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1203 D.t3267 G.t1203 S.t3403 S.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1204 S.t3402 G.t1204 D.t3031 S.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1205 D.t2910 G.t1205 S.t3401 S.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1206 S.t3400 G.t1206 D.t4347 S.t443 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1207 D.t4338 G.t1207 S.t3399 S.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1208 D.t2727 G.t1208 S.t3398 S.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1209 D.t3133 G.t1209 S.t3397 S.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1210 S.t3396 G.t1210 D.t2770 S.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1211 D.t2786 G.t1211 S.t3395 S.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1212 S.t3394 G.t1212 D.t2845 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1213 D.t2899 G.t1213 S.t3393 S.t388 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1214 S.t3392 G.t1214 D.t3025 S.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1215 S.t3391 G.t1215 D.t3120 S.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1216 D.t2951 G.t1216 S.t3390 S.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1217 D.t3023 G.t1217 S.t3389 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1218 S.t3388 G.t1218 D.t2778 S.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1219 D.t2876 G.t1219 S.t3387 S.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1220 D.t2904 G.t1220 S.t3386 S.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1221 D.t2921 G.t1221 S.t3385 S.t216 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1222 S.t3384 G.t1222 D.t3000 S.t79 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1223 D.t3048 G.t1223 S.t3383 S.t176 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1224 D.t3140 G.t1224 S.t3382 S.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1225 D.t2945 G.t1225 S.t3381 S.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1226 S.t3380 G.t1226 D.t2994 S.t270 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1227 D.t3009 G.t1227 S.t3379 S.t321 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1228 S.t3378 G.t1228 D.t3019 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1229 S.t3377 G.t1229 D.t2938 S.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1230 D.t2934 G.t1230 S.t3376 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1231 S.t3375 G.t1231 D.t2959 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1232 D.t4391 G.t1232 S.t3374 S.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1233 D.t2842 G.t1233 S.t3373 S.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1234 D.t2886 G.t1234 S.t3372 S.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1235 D.t3158 G.t1235 S.t3371 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1236 D.t4164 G.t1236 S.t3370 S.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1237 S.t3369 G.t1237 D.t3167 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1238 D.t4335 G.t1238 S.t3368 S.t150 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1239 D.t4340 G.t1239 S.t3367 S.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1240 S.t3366 G.t1240 D.t4398 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1241 D.t4411 G.t1241 S.t3365 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1242 S.t3364 G.t1242 D.t2993 S.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1243 D.t2797 G.t1243 S.t3363 S.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1244 S.t3362 G.t1244 D.t2863 S.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1245 S.t3361 G.t1245 D.t3044 S.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1246 D.t3118 G.t1246 S.t3360 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1247 D.t3165 G.t1247 S.t3359 S.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1248 S.t3358 G.t1248 D.t3106 S.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1249 S.t3357 G.t1249 D.t2800 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1250 D.t3128 G.t1250 S.t3356 S.t388 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1251 D.t2997 G.t1251 S.t3355 S.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1252 D.t2774 G.t1252 S.t3354 S.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1253 D.t2841 G.t1253 S.t3353 S.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1254 S.t3352 G.t1254 D.t2733 S.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1255 D.t3051 G.t1255 S.t3351 S.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1256 S.t3350 G.t1256 D.t2949 S.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1257 D.t3134 G.t1257 S.t3349 S.t209 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1258 D.t2756 G.t1258 S.t3348 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1259 S.t3347 G.t1259 D.t3114 S.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1260 D.t3125 G.t1260 S.t3346 S.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1261 S.t3345 G.t1261 D.t2980 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1262 D.t4392 G.t1262 S.t3344 S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1263 S.t3343 G.t1263 D.t3071 S.t231 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1264 D.t2851 G.t1264 S.t3342 S.t231 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1265 D.t2796 G.t1265 S.t3341 S.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1266 S.t3340 G.t1266 D.t2782 S.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1267 D.t3094 G.t1267 S.t3339 S.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1268 S.t3338 G.t1268 D.t2882 S.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1269 S.t3337 G.t1269 D.t2781 S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1270 S.t3336 G.t1270 D.t2855 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1271 D.t3141 G.t1271 S.t3335 S.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1272 S.t3334 G.t1272 D.t2885 S.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1273 S.t3333 G.t1273 D.t2942 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1274 S.t3332 G.t1274 D.t2780 S.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1275 S.t3331 G.t1275 D.t3150 S.t218 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1276 D.t2868 G.t1276 S.t3330 S.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1277 S.t3329 G.t1277 D.t2977 S.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1278 D.t3138 G.t1278 S.t3328 S.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1279 S.t3327 G.t1279 D.t2831 S.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1280 S.t3326 G.t1280 D.t2888 S.t209 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1281 D.t3063 G.t1281 S.t3325 S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1282 S.t3324 G.t1282 D.t2943 S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1283 S.t3323 G.t1283 D.t2805 S.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1284 S.t3322 G.t1284 D.t3135 S.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1285 S.t3321 G.t1285 D.t2990 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1286 D.t2809 G.t1286 S.t3320 S.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1287 S.t3319 G.t1287 D.t2900 S.t198 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1288 D.t3018 G.t1288 S.t3318 S.t176 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1289 D.t2950 G.t1289 S.t3317 S.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1290 D.t2879 G.t1290 S.t3316 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1291 D.t2872 G.t1291 S.t3315 S.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1292 S.t3314 G.t1292 D.t2772 S.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1293 D.t3157 G.t1293 S.t3313 S.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1294 S.t3312 G.t1294 D.t3045 S.t183 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1295 S.t3311 G.t1295 D.t2871 S.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1296 D.t2835 G.t1296 S.t3310 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1297 D.t2893 G.t1297 S.t3309 S.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1298 D.t2937 G.t1298 S.t3308 S.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1299 S.t3307 G.t1299 D.t3153 S.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1300 D.t3090 G.t1300 S.t3306 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1301 D.t3164 G.t1301 S.t3305 S.t183 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1302 S.t3304 G.t1302 D.t2776 S.t270 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1303 S.t3303 G.t1303 D.t3039 S.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1304 D.t3049 G.t1304 S.t3302 S.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1305 S.t3301 G.t1305 D.t2946 S.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1306 S.t3300 G.t1306 D.t2790 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1307 D.t2957 G.t1307 S.t3299 S.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1308 S.t3298 G.t1308 D.t3002 S.t332 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1309 D.t2898 G.t1309 S.t3297 S.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1310 D.t2965 G.t1310 S.t3296 S.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1311 D.t2866 G.t1311 S.t3295 S.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1312 D.t2777 G.t1312 S.t3294 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1313 S.t3293 G.t1313 D.t2869 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1314 D.t2761 G.t1314 S.t3292 S.t321 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1315 S.t3291 G.t1315 D.t2754 S.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1316 D.t2787 G.t1316 S.t3290 S.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1317 S.t3289 G.t1317 D.t3057 S.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1318 S.t3288 G.t1318 D.t3015 S.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1319 S.t3287 G.t1319 D.t2799 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1320 S.t3286 G.t1320 D.t2865 S.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1321 D.t2917 G.t1321 S.t3285 S.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1322 D.t2861 G.t1322 S.t3284 S.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1323 S.t3283 G.t1323 D.t2783 S.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1324 D.t2901 G.t1324 S.t3282 S.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1325 S.t3281 G.t1325 D.t3041 S.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1326 D.t3115 G.t1326 S.t3280 S.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1327 S.t3279 G.t1327 D.t3052 S.t150 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1328 S.t3278 G.t1328 D.t2766 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1329 D.t2975 G.t1329 S.t3277 S.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1330 S.t3276 G.t1330 D.t2850 S.t139 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1331 S.t3275 G.t1331 D.t2953 S.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1332 S.t3274 G.t1332 D.t3058 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1333 D.t2887 G.t1333 S.t3273 S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1334 S.t3272 G.t1334 D.t3008 S.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1335 D.t2823 G.t1335 S.t3271 S.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1336 S.t3270 G.t1336 D.t3062 S.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1337 S.t3269 G.t1337 D.t3117 S.t216 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1338 S.t3268 G.t1338 D.t2817 S.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1339 D.t3124 G.t1339 S.t3267 S.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1340 D.t3162 G.t1340 S.t3266 S.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1341 S.t3265 G.t1341 D.t2998 S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1342 D.t3037 G.t1342 S.t3264 S.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1343 S.t3263 G.t1343 D.t2974 S.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1344 S.t3262 G.t1344 D.t2987 S.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1345 S.t3261 G.t1345 D.t2874 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1346 D.t2944 G.t1346 S.t3260 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1347 S.t3259 G.t1347 D.t2794 S.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1348 D.t3064 G.t1348 S.t3258 S.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1349 D.t3148 G.t1349 S.t3257 S.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1350 D.t3113 G.t1350 S.t3256 S.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1351 D.t4389 G.t1351 S.t3255 S.t538 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1352 S.t3254 G.t1352 D.t3059 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1353 D.t2819 G.t1353 S.t3253 S.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1354 D.t2895 G.t1354 S.t3252 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1355 S.t3251 G.t1355 D.t3109 S.t79 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1356 S.t3250 G.t1356 D.t2952 S.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1357 D.t2813 G.t1357 S.t3249 S.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1358 D.t2929 G.t1358 S.t3248 S.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1359 D.t2978 G.t1359 S.t3247 S.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1360 S.t3246 G.t1360 D.t2988 S.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1361 S.t3245 G.t1361 D.t2996 S.t270 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1362 S.t3244 G.t1362 D.t2684 S.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1363 S.t3243 G.t1363 D.t2839 S.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1364 D.t2889 G.t1364 S.t3242 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1365 S.t3241 G.t1365 D.t3137 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1366 S.t3240 G.t1366 D.t3050 S.t79 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1367 D.t2981 G.t1367 S.t3239 S.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1368 D.t2982 G.t1368 S.t3238 S.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1369 D.t2859 G.t1369 S.t3237 S.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1370 S.t3236 G.t1370 D.t2969 S.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1371 D.t3020 G.t1371 S.t3235 S.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1372 D.t3053 G.t1372 S.t3234 S.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1373 S.t3233 G.t1373 D.t3073 S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1374 D.t3126 G.t1374 S.t3232 S.t150 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1375 S.t3231 G.t1375 D.t2856 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1376 D.t2925 G.t1376 S.t3230 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1377 S.t3229 G.t1377 D.t3132 S.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1378 D.t2806 G.t1378 S.t3228 S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1379 S.t3227 G.t1379 D.t3055 S.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1380 S.t3226 G.t1380 D.t2811 S.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1381 D.t2878 G.t1381 S.t3225 S.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1382 D.t2864 G.t1382 S.t3224 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1383 S.t3223 G.t1383 D.t2918 S.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1384 S.t3222 G.t1384 D.t2936 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1385 D.t2906 G.t1385 S.t3221 S.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1386 D.t3046 G.t1386 S.t3220 S.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1387 S.t3219 G.t1387 D.t3029 S.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1388 S.t3218 G.t1388 D.t3036 S.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1389 S.t3217 G.t1389 D.t3149 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1390 D.t2971 G.t1390 S.t3216 S.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1391 S.t3215 G.t1391 D.t3047 S.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1392 D.t2837 G.t1392 S.t3214 S.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1393 S.t3213 G.t1393 D.t2822 S.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1394 D.t2939 G.t1394 S.t3212 S.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1395 S.t3211 G.t1395 D.t3122 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1396 S.t3210 G.t1396 D.t3121 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1397 D.t3127 G.t1397 S.t3209 S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1398 S.t3208 G.t1398 D.t3139 S.t231 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1399 S.t3207 G.t1399 D.t4395 S.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1400 D.t2816 G.t1400 S.t3206 S.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1401 S.t3205 G.t1401 D.t3011 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1402 S.t3204 G.t1402 D.t3072 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1403 S.t3203 G.t1403 D.t3092 S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1404 S.t3202 G.t1404 D.t2928 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1405 S.t3201 G.t1405 D.t2966 S.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1406 S.t3200 G.t1406 D.t2986 S.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1407 S.t3199 G.t1407 D.t3060 S.t218 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1408 S.t3198 G.t1408 D.t3078 S.t216 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1409 S.t3197 G.t1409 D.t3080 S.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1410 D.t3101 G.t1410 S.t3196 S.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1411 S.t3195 G.t1411 D.t2915 S.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1412 S.t3194 G.t1412 D.t2807 S.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1413 S.t3193 G.t1413 D.t2847 S.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1414 S.t3192 G.t1414 D.t2843 S.t158 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1415 S.t3191 G.t1415 D.t2884 S.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1416 S.t3190 G.t1416 D.t2897 S.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1417 D.t2931 G.t1417 S.t3189 S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1418 S.t3188 G.t1418 D.t2908 S.t209 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1419 S.t3187 G.t1419 D.t2852 S.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1420 S.t3186 G.t1420 D.t2829 S.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1421 D.t2956 G.t1421 S.t3185 S.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1422 D.t3068 G.t1422 S.t3184 S.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1423 S.t3183 G.t1423 D.t2808 S.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1424 D.t2791 G.t1424 S.t3182 S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1425 D.t2779 G.t1425 S.t3181 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1426 D.t2803 G.t1426 S.t3180 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1427 S.t3179 G.t1427 D.t2960 S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1428 S.t3178 G.t1428 D.t3154 S.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1429 D.t3156 G.t1429 S.t3177 S.t538 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1430 S.t3176 G.t1430 D.t3056 S.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1431 D.t2857 G.t1431 S.t3175 S.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1432 S.t3174 G.t1432 D.t2775 S.t183 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1433 S.t3173 G.t1433 D.t2970 S.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1434 D.t2992 G.t1434 S.t3172 S.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1435 D.t3142 G.t1435 S.t3171 S.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1436 S.t3170 G.t1436 D.t3040 S.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1437 S.t3169 G.t1437 D.t3054 S.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1438 D.t3061 G.t1438 S.t3168 S.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1439 D.t3066 G.t1439 S.t3167 S.t183 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1440 S.t3166 G.t1440 D.t3084 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1441 D.t3086 G.t1441 S.t3165 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1442 S.t3164 G.t1442 D.t3103 S.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1443 D.t3035 G.t1443 S.t3163 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1444 D.t2941 G.t1444 S.t3162 S.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1445 S.t3161 G.t1445 D.t2948 S.t176 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1446 D.t2983 G.t1446 S.t3160 S.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1447 D.t2989 G.t1447 S.t3159 S.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1448 S.t3158 G.t1448 D.t3005 S.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1449 S.t3157 G.t1449 D.t3016 S.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1450 D.t3032 G.t1450 S.t3156 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1451 S.t3155 G.t1451 D.t2919 S.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1452 D.t2846 G.t1452 S.t3154 S.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1453 D.t2862 G.t1453 S.t3153 S.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1454 D.t2870 G.t1454 S.t3152 S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1455 S.t3151 G.t1455 D.t2883 S.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1456 D.t2891 G.t1456 S.t3150 S.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1457 S.t3149 G.t1457 D.t3096 S.t158 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1458 D.t3095 G.t1458 S.t3148 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1459 S.t3147 G.t1459 D.t2854 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1460 D.t2792 G.t1460 S.t3146 S.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1461 S.t3145 G.t1461 D.t2795 S.t150 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1462 D.t2798 G.t1462 S.t3144 S.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1463 D.t3030 G.t1463 S.t3143 S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1464 S.t3142 G.t1464 D.t2826 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1465 D.t2832 G.t1465 S.t3141 S.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1466 S.t3140 G.t1466 D.t2840 S.t139 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1467 S.t3139 G.t1467 D.t2769 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1468 S.t3138 G.t1468 D.t2844 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1469 S.t3137 G.t1469 D.t2873 S.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1470 S.t3136 G.t1470 D.t2785 S.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1471 S.t3135 G.t1471 D.t3003 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1472 D.t3010 G.t1472 S.t3134 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1473 D.t2815 G.t1473 S.t3133 S.t79 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1474 S.t3132 G.t1474 D.t2812 S.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1475 S.t3131 G.t1475 D.t2767 S.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1476 S.t3130 G.t1476 D.t4387 S.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1477 D.t4333 G.t1477 S.t3129 S.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1478 S.t3128 G.t1478 D.t2905 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1479 S.t3127 G.t1479 D.t3065 S.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1480 S.t3126 G.t1480 D.t2890 S.t158 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1481 S.t3125 G.t1481 D.t3143 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1482 S.t3124 G.t1482 D.t3152 S.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1483 S.t3123 G.t1483 D.t4328 S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1484 S.t3122 G.t1484 D.t4163 S.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1485 S.t3121 G.t1485 D.t4355 S.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1486 D.t4410 G.t1486 S.t3120 S.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1487 S.t3119 G.t1487 D.t4386 S.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1488 S.t3118 G.t1488 D.t4344 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1489 D.t4293 G.t1489 S.t3117 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1490 S.t3116 G.t1490 D.t4334 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1491 S.t3115 G.t1491 D.t1207 S.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1492 S.t3114 G.t1492 D.t3151 S.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1493 S.t3113 G.t1493 D.t3155 S.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1494 D.t3161 G.t1494 S.t3112 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1495 S.t3111 G.t1495 D.t2912 S.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1496 D.t3079 G.t1496 S.t3110 S.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1497 S.t3109 G.t1497 D.t3082 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1498 D.t1185 G.t1498 S.t3108 S.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1499 S.t3107 G.t1499 D.t3146 S.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1500 S.t3106 G.t1500 D.t3110 S.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1501 S.t3105 G.t1501 D.t3119 S.t79 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1502 S.t3104 G.t1502 D.t3123 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1503 D.t3129 G.t1503 S.t3103 S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1504 D.t3131 G.t1504 S.t3102 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1505 D.t3136 G.t1505 S.t3101 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1506 S.t3100 G.t1506 D.t3144 S.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1507 S.t3099 G.t1507 D.t3105 S.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1508 S.t3098 G.t1508 D.t3087 S.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1509 S.t3097 G.t1509 D.t3089 S.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1510 S.t3096 G.t1510 D.t3091 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1511 D.t3093 G.t1511 S.t3095 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1512 S.t3094 G.t1512 D.t3097 S.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1513 S.t3093 G.t1513 D.t3100 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1514 S.t3092 G.t1514 D.t3102 S.t79 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1515 S.t3091 G.t1515 D.t3085 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1516 D.t3001 G.t1516 S.t3090 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1517 S.t3089 G.t1517 D.t3004 S.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1518 S.t3088 G.t1518 D.t3007 S.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1519 D.t3013 G.t1519 S.t3087 S.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1520 S.t3086 G.t1520 D.t3027 S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1521 D.t3038 G.t1521 S.t3085 S.t231 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1522 D.t3083 G.t1522 S.t3084 S.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1523 S.t3083 G.t1523 D.t2991 S.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1524 S.t3082 G.t1524 D.t2920 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1525 D.t2924 G.t1525 S.t3081 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1526 D.t2935 G.t1526 S.t3080 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1527 S.t3079 G.t1527 D.t2955 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1528 D.t2964 G.t1528 S.t3078 S.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1529 D.t2968 G.t1529 S.t3077 S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1530 S.t3076 G.t1530 D.t2973 S.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1531 S.t3075 G.t1531 D.t2916 S.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1532 S.t3074 G.t1532 D.t2768 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1533 S.t3073 G.t1533 D.t2788 S.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1534 D.t2804 G.t1534 S.t3072 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1535 S.t3071 G.t1535 D.t2828 S.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1536 D.t2853 G.t1536 S.t3070 S.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1537 S.t3069 G.t1537 D.t2894 S.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1538 S.t3068 G.t1538 D.t2914 S.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1539 S.t3067 G.t1539 D.t3529 S.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1540 D.t1497 G.t1540 S.t3066 S.t443 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1541 S.t3065 G.t1541 D.t1496 S.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1542 S.t3064 G.t1542 D.t1495 S.t209 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1543 S.t3063 G.t1543 D.t1494 S.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1544 S.t3062 G.t1544 D.t1668 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1545 S.t3061 G.t1545 D.t1667 S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1546 D.t1666 G.t1546 S.t3060 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1547 D.t1665 G.t1547 S.t3059 S.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1548 S.t3058 G.t1548 D.t1664 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1549 S.t3057 G.t1549 D.t1663 S.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1550 D.t1662 G.t1550 S.t3056 S.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1551 D.t1661 G.t1551 S.t3055 S.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1552 D.t1733 G.t1552 S.t3054 S.t443 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1553 S.t3053 G.t1553 D.t1732 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1554 D.t1731 G.t1554 S.t3052 S.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1555 S.t3051 G.t1555 D.t1730 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1556 S.t3050 G.t1556 D.t1729 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1557 S.t3049 G.t1557 D.t1728 S.t538 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1558 S.t3048 G.t1558 D.t1727 S.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1559 S.t3047 G.t1559 D.t1726 S.t218 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1560 D.t562 G.t1560 S.t3046 S.t79 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1561 S.t3045 G.t1561 D.t561 S.t218 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1562 S.t3044 G.t1562 D.t560 S.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1563 D.t559 G.t1563 S.t3043 S.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1564 S.t3042 G.t1564 D.t558 S.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1565 S.t3041 G.t1565 D.t557 S.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1566 S.t3040 G.t1566 D.t556 S.t183 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1567 D.t555 G.t1567 S.t3039 S.t139 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1568 S.t3038 G.t1568 D.t550 S.t158 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1569 S.t3037 G.t1569 D.t549 S.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1570 S.t3036 G.t1570 D.t548 S.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1571 S.t3035 G.t1571 D.t547 S.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1572 D.t546 G.t1572 S.t3034 S.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1573 D.t545 G.t1573 S.t3033 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1574 S.t3032 G.t1574 D.t544 S.t209 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1575 S.t3031 G.t1575 D.t543 S.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1576 D.t583 G.t1576 S.t3030 S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1577 S.t3029 G.t1577 D.t582 S.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1578 S.t3028 G.t1578 D.t581 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1579 D.t580 G.t1579 S.t3027 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1580 S.t3026 G.t1580 D.t579 S.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1581 D.t578 G.t1581 S.t3025 S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1582 D.t577 G.t1582 S.t3024 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1583 D.t576 G.t1583 S.t3023 S.t406 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1584 D.t725 G.t1584 S.t3022 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1585 S.t3021 G.t1585 D.t724 S.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1586 D.t723 G.t1586 S.t3020 S.t198 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1587 D.t722 G.t1587 S.t3019 S.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1588 S.t3018 G.t1588 D.t721 S.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1589 S.t3017 G.t1589 D.t720 S.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1590 D.t719 G.t1590 S.t3016 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1591 D.t718 G.t1591 S.t3015 S.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1592 S.t3014 G.t1592 D.t1391 S.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1593 S.t3013 G.t1593 D.t1390 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1594 D.t1389 G.t1594 S.t3012 S.t150 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1595 S.t3011 G.t1595 D.t1388 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1596 D.t1387 G.t1596 S.t3010 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1597 S.t3009 G.t1597 D.t1386 S.t176 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1598 D.t1385 G.t1598 S.t3008 S.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1599 S.t3007 G.t1599 D.t1599 S.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1600 D.t1598 G.t1600 S.t3006 S.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1601 D.t1597 G.t1601 S.t3005 S.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1602 D.t1596 G.t1602 S.t3004 S.t332 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1603 D.t1595 G.t1603 S.t3003 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1604 S.t3002 G.t1604 D.t1594 S.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1605 D.t1593 G.t1605 S.t3001 S.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1606 D.t1369 G.t1606 S.t3000 S.t231 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1607 D.t1368 G.t1607 S.t2999 S.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1608 D.t1367 G.t1608 S.t2998 S.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1609 S.t2997 G.t1609 D.t1366 S.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1610 D.t1365 G.t1610 S.t2996 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1611 S.t2995 G.t1611 D.t1364 S.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1612 S.t2994 G.t1612 D.t1363 S.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1613 D.t1645 G.t1613 S.t2993 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1614 D.t1644 G.t1614 S.t2992 S.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1615 D.t1643 G.t1615 S.t2991 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1616 S.t2990 G.t1616 D.t1642 S.t158 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1617 D.t1641 G.t1617 S.t2989 S.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1618 D.t1640 G.t1618 S.t2988 S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1619 S.t2987 G.t1619 D.t740 S.t388 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1620 D.t739 G.t1620 S.t2986 S.t218 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1621 D.t738 G.t1621 S.t2985 S.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1622 S.t2984 G.t1622 D.t737 S.t150 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1623 S.t2983 G.t1623 D.t736 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1624 D.t735 G.t1624 S.t2982 S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1625 S.t2981 G.t1625 D.t680 S.t209 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1626 D.t679 G.t1626 S.t2980 S.t209 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1627 S.t2979 G.t1627 D.t678 S.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1628 S.t2978 G.t1628 D.t677 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1629 S.t2977 G.t1629 D.t676 S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1630 S.t2976 G.t1630 D.t675 S.t357 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1631 S.t2975 G.t1631 D.t279 S.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1632 D.t278 G.t1632 S.t2974 S.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1633 D.t277 G.t1633 S.t2973 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1634 S.t2972 G.t1634 D.t276 S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1635 D.t275 G.t1635 S.t2971 S.t79 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1636 S.t2970 G.t1636 D.t274 S.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1637 D.t1397 G.t1637 S.t2969 S.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1638 D.t1396 G.t1638 S.t2968 S.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1639 S.t2967 G.t1639 D.t1395 S.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1640 S.t2966 G.t1640 D.t1394 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1641 S.t2965 G.t1641 D.t1393 S.t321 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1642 D.t1392 G.t1642 S.t2964 S.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1643 D.t1918 G.t1643 S.t2963 S.t79 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1644 D.t1917 G.t1644 S.t2962 S.t216 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1645 S.t2961 G.t1645 D.t1916 S.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1646 S.t2960 G.t1646 D.t1915 S.t218 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1647 S.t2959 G.t1647 D.t1914 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1648 D.t1913 G.t1648 S.t2958 S.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1649 S.t2957 G.t1649 D.t405 S.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1650 S.t2956 G.t1650 D.t404 S.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1651 D.t403 G.t1651 S.t2955 S.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1652 S.t2954 G.t1652 D.t402 S.t183 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1653 S.t2953 G.t1653 D.t401 S.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1654 D.t400 G.t1654 S.t2952 S.t139 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1655 D.t1616 G.t1655 S.t2951 S.t406 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1656 D.t1615 G.t1656 S.t2950 S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1657 D.t1614 G.t1657 S.t2949 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1658 D.t1613 G.t1658 S.t2948 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1659 D.t1612 G.t1659 S.t2947 S.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1660 S.t2946 G.t1660 D.t1611 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1661 D.t805 G.t1661 S.t2945 S.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1662 S.t2944 G.t1662 D.t804 S.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1663 S.t2943 G.t1663 D.t803 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1664 D.t802 G.t1664 S.t2942 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1665 D.t801 G.t1665 S.t2941 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1666 D.t800 G.t1666 S.t2940 S.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1667 S.t2939 G.t1667 D.t2572 S.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1668 S.t2938 G.t1668 D.t2571 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1669 D.t2570 G.t1669 S.t2937 S.t270 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1670 D.t2569 G.t1670 S.t2936 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1671 S.t2935 G.t1671 D.t2568 S.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1672 S.t2934 G.t1672 D.t2567 S.t79 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1673 D.t209 G.t1673 S.t2933 S.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1674 D.t208 G.t1674 S.t2932 S.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1675 S.t2931 G.t1675 D.t207 S.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1676 D.t206 G.t1676 S.t2930 S.t332 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1677 S.t2929 G.t1677 D.t205 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1678 D.t204 G.t1678 S.t2928 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1679 S.t2927 G.t1679 D.t2330 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1680 S.t2926 G.t1680 D.t2329 S.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1681 D.t2328 G.t1681 S.t2925 S.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1682 D.t2327 G.t1682 S.t2924 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1683 S.t2923 G.t1683 D.t2326 S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1684 D.t2325 G.t1684 S.t2922 S.t150 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1685 S.t2921 G.t1685 D.t1930 S.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1686 D.t1929 G.t1686 S.t2920 S.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1687 S.t2919 G.t1687 D.t1928 S.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1688 D.t1927 G.t1688 S.t2918 S.t198 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1689 D.t1926 G.t1689 S.t2917 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1690 D.t1925 G.t1690 S.t2916 S.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1691 D.t1909 G.t1691 S.t2915 S.t216 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1692 D.t1908 G.t1692 S.t2914 S.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1693 D.t1907 G.t1693 S.t2913 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1694 D.t1906 G.t1694 S.t2912 S.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1695 D.t1905 G.t1695 S.t2911 S.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1696 D.t1904 G.t1696 S.t2910 S.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1697 D.t1568 G.t1697 S.t2909 S.t218 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1698 S.t2908 G.t1698 D.t1567 S.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1699 D.t1566 G.t1699 S.t2907 S.t443 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1700 D.t1565 G.t1700 S.t2906 S.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1701 D.t1564 G.t1701 S.t2905 S.t158 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1702 D.t2522 G.t1702 S.t2904 S.t270 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1703 D.t2521 G.t1703 S.t2903 S.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1704 D.t2520 G.t1704 S.t2902 S.t321 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1705 D.t2519 G.t1705 S.t2901 S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1706 S.t2900 G.t1706 D.t2518 S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1707 D.t846 G.t1707 S.t2899 S.t209 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1708 D.t845 G.t1708 S.t2898 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1709 S.t2897 G.t1709 D.t844 S.t388 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1710 S.t2896 G.t1710 D.t843 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1711 S.t2895 G.t1711 D.t842 S.t357 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1712 D.t921 G.t1712 S.t2894 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1713 D.t920 G.t1713 S.t2893 S.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1714 S.t2892 G.t1714 D.t919 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1715 D.t918 G.t1715 S.t2891 S.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1716 D.t917 G.t1716 S.t2890 S.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1717 D.t891 G.t1717 S.t2889 S.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1718 D.t890 G.t1718 S.t2888 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1719 S.t2887 G.t1719 D.t889 S.t538 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1720 D.t888 G.t1720 S.t2886 S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1721 D.t887 G.t1721 S.t2885 S.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1722 S.t2884 G.t1722 D.t826 S.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1723 D.t825 G.t1723 S.t2883 S.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1724 D.t824 G.t1724 S.t2882 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1725 D.t823 G.t1725 S.t2881 S.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1726 S.t2880 G.t1726 D.t822 S.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1727 S.t2879 G.t1727 D.t1347 S.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1728 D.t1346 G.t1728 S.t2878 S.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1729 D.t1345 G.t1729 S.t2877 S.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1730 D.t1344 G.t1730 S.t2876 S.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1731 S.t2875 G.t1731 D.t1343 S.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1732 S.t2874 G.t1732 D.t1330 S.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1733 S.t2873 G.t1733 D.t1329 S.t321 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1734 D.t1328 G.t1734 S.t2872 S.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1735 D.t1327 G.t1735 S.t2871 S.t139 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1736 D.t1326 G.t1736 S.t2870 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1737 D.t455 G.t1737 S.t2869 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1738 D.t454 G.t1738 S.t2868 S.t176 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1739 D.t453 G.t1739 S.t2867 S.t79 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1740 S.t2866 G.t1740 D.t452 S.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1741 D.t451 G.t1741 S.t2865 S.t216 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1742 S.t2864 G.t1742 D.t693 S.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1743 S.t2863 G.t1743 D.t692 S.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1744 D.t691 G.t1744 S.t2862 S.t406 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1745 D.t690 G.t1745 S.t2861 S.t406 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1746 D.t689 G.t1746 S.t2860 S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1747 D.t730 G.t1747 S.t2859 S.t198 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1748 S.t2858 G.t1748 D.t729 S.t176 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1749 S.t2857 G.t1749 D.t728 S.t150 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1750 D.t727 G.t1750 S.t2856 S.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1751 S.t2855 G.t1751 D.t726 S.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1752 D.t395 G.t1752 S.t2854 S.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1753 S.t2853 G.t1753 D.t394 S.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1754 D.t393 G.t1754 S.t2852 S.t332 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1755 D.t392 G.t1755 S.t2851 S.t158 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1756 D.t391 G.t1756 S.t2850 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1757 D.t410 G.t1757 S.t2849 S.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1758 D.t409 G.t1758 S.t2848 S.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1759 D.t408 G.t1759 S.t2847 S.t150 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1760 D.t407 G.t1760 S.t2846 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1761 D.t406 G.t1761 S.t2845 S.t270 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1762 S.t2844 G.t1762 D.t948 S.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1763 S.t2843 G.t1763 D.t947 S.t176 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1764 D.t946 G.t1764 S.t2842 S.t198 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1765 D.t945 G.t1765 S.t2841 S.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1766 D.t944 G.t1766 S.t2840 S.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1767 D.t931 G.t1767 S.t2839 S.t209 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1768 D.t930 G.t1768 S.t2838 S.t332 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1769 S.t2837 G.t1769 D.t929 S.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1770 D.t928 G.t1770 S.t2836 S.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1771 D.t927 G.t1771 S.t2835 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1772 D.t953 G.t1772 S.t2834 S.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1773 D.t952 G.t1773 S.t2833 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1774 S.t2832 G.t1774 D.t951 S.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1775 D.t950 G.t1775 S.t2831 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1776 S.t2830 G.t1776 D.t949 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1777 S.t2829 G.t1777 D.t943 S.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1778 D.t942 G.t1778 S.t2828 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1779 D.t941 G.t1779 S.t2827 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1780 D.t940 G.t1780 S.t2826 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1781 D.t939 G.t1781 S.t2825 S.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1782 S.t2824 G.t1782 D.t936 S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1783 D.t935 G.t1783 S.t2823 S.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1784 S.t2822 G.t1784 D.t934 S.t158 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1785 D.t933 G.t1785 S.t2821 S.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1786 D.t932 G.t1786 S.t2820 S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1787 S.t2819 G.t1787 D.t916 S.t388 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1788 D.t915 G.t1788 S.t2818 S.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1789 D.t914 G.t1789 S.t2817 S.t218 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1790 D.t913 G.t1790 S.t2816 S.t218 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1791 D.t912 G.t1791 S.t2815 S.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1792 S.t2814 G.t1792 D.t906 S.t79 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1793 S.t2813 G.t1793 D.t905 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1794 D.t904 G.t1794 S.t2812 S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1795 D.t903 G.t1795 S.t2811 S.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1796 D.t902 G.t1796 S.t2810 S.t158 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1797 D.t810 G.t1797 S.t2809 S.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1798 D.t809 G.t1798 S.t2808 S.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1799 S.t2807 G.t1799 D.t808 S.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1800 D.t807 G.t1800 S.t2806 S.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1801 D.t806 G.t1801 S.t2805 S.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1802 S.t2804 G.t1802 D.t364 S.t139 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1803 S.t2803 G.t1803 D.t363 S.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1804 D.t362 G.t1804 S.t2802 S.t209 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1805 S.t2801 G.t1805 D.t361 S.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1806 S.t2800 G.t1806 D.t360 S.t357 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1807 D.t242 G.t1807 S.t2799 S.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1808 D.t241 G.t1808 S.t2798 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1809 S.t2797 G.t1809 D.t240 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1810 D.t239 G.t1810 S.t2796 S.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1811 S.t2795 G.t1811 D.t238 S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1812 D.t633 G.t1812 S.t2794 S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1813 D.t632 G.t1813 S.t2793 S.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1814 D.t631 G.t1814 S.t2792 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1815 D.t630 G.t1815 S.t2791 S.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1816 D.t629 G.t1816 S.t2790 S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1817 S.t2789 G.t1817 D.t1725 S.t321 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1818 D.t1724 G.t1818 S.t2788 S.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1819 D.t1723 G.t1819 S.t2787 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1820 S.t2786 G.t1820 D.t1722 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1821 S.t2785 G.t1821 D.t1721 S.t332 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1822 D.t1528 G.t1822 S.t2784 S.t216 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1823 S.t2783 G.t1823 D.t1527 S.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1824 D.t1526 G.t1824 S.t2782 S.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1825 S.t2781 G.t1825 D.t1525 S.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1826 S.t2780 G.t1826 D.t1524 S.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1827 D.t509 G.t1827 S.t2779 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1828 S.t2778 G.t1828 D.t508 S.t198 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1829 D.t507 G.t1829 S.t2777 S.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1830 D.t506 G.t1830 S.t2776 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1831 S.t2775 G.t1831 D.t505 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1832 S.t2774 G.t1832 D.t537 S.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1833 D.t536 G.t1833 S.t2773 S.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1834 D.t535 G.t1834 S.t2772 S.t176 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1835 D.t534 G.t1835 S.t2771 S.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1836 S.t2770 G.t1836 D.t533 S.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1837 S.t2769 G.t1837 D.t572 S.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1838 D.t571 G.t1838 S.t2768 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1839 S.t2767 G.t1839 D.t570 S.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1840 D.t569 G.t1840 S.t2766 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1841 S.t2765 G.t1841 D.t568 S.t176 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1842 D.t650 G.t1842 S.t2764 S.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1843 D.t649 G.t1843 S.t2763 S.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1844 D.t648 G.t1844 S.t2762 S.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1845 S.t2761 G.t1845 D.t647 S.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1846 S.t2760 G.t1846 D.t646 S.t443 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1847 S.t2759 G.t1847 D.t608 S.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1848 S.t2758 G.t1848 D.t607 S.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1849 S.t2757 G.t1849 D.t606 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1850 D.t605 G.t1850 S.t2756 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1851 D.t667 G.t1851 S.t2755 S.t158 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1852 D.t666 G.t1852 S.t2754 S.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1853 D.t665 G.t1853 S.t2753 S.t332 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1854 S.t2752 G.t1854 D.t664 S.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1855 S.t2751 G.t1855 D.t1484 S.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1856 D.t1483 G.t1856 S.t2750 S.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1857 D.t1482 G.t1857 S.t2749 S.t388 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1858 D.t1481 G.t1858 S.t2748 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1859 S.t2747 G.t1859 D.t1468 S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1860 S.t2746 G.t1860 D.t1467 S.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1861 D.t1466 G.t1861 S.t2745 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1862 S.t2744 G.t1862 D.t1465 S.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1863 D.t1452 G.t1863 S.t2743 S.t198 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1864 S.t2742 G.t1864 D.t1451 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1865 D.t1450 G.t1865 S.t2741 S.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1866 S.t2740 G.t1866 D.t1449 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1867 S.t2739 G.t1867 D.t1436 S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1868 D.t1435 G.t1868 S.t2738 S.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1869 D.t1434 G.t1869 S.t2737 S.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1870 D.t1433 G.t1870 S.t2736 S.t216 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1871 D.t1420 G.t1871 S.t2735 S.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1872 S.t2734 G.t1872 D.t1419 S.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1873 S.t2733 G.t1873 D.t1418 S.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1874 S.t2732 G.t1874 D.t1417 S.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1875 D.t1404 G.t1875 S.t2731 S.t443 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1876 D.t1403 G.t1876 S.t2730 S.t321 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1877 D.t1402 G.t1877 S.t2729 S.t158 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1878 D.t1401 G.t1878 S.t2728 S.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1879 D.t3516 G.t1879 S.t2727 S.t270 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1880 D.t3515 G.t1880 S.t2726 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1881 S.t2725 G.t1881 D.t3514 S.t216 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1882 D.t3513 G.t1882 S.t2724 S.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1883 S.t2723 G.t1883 D.t3396 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1884 S.t2722 G.t1884 D.t3395 S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1885 D.t3394 G.t1885 S.t2721 S.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1886 D.t3393 G.t1886 S.t2720 S.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1887 D.t3243 G.t1887 S.t2719 S.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1888 S.t2718 G.t1888 D.t3242 S.t406 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1889 D.t3241 G.t1889 S.t2717 S.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1890 D.t3240 G.t1890 S.t2716 S.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1891 S.t2715 G.t1891 D.t3400 S.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1892 S.t2714 G.t1892 D.t3399 S.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1893 S.t2713 G.t1893 D.t3398 S.t198 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1894 D.t3397 G.t1894 S.t2712 S.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1895 S.t2711 G.t1895 D.t3315 S.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1896 D.t3314 G.t1896 S.t2710 S.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1897 S.t2709 G.t1897 D.t3313 S.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1898 D.t3312 G.t1898 S.t2708 S.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1899 D.t3924 G.t1899 S.t2707 S.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1900 S.t2706 G.t1900 D.t3923 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1901 D.t3922 G.t1901 S.t2705 S.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1902 D.t3921 G.t1902 S.t2704 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1903 D.t3547 G.t1903 S.t2703 S.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1904 D.t3546 G.t1904 S.t2702 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1905 S.t2701 G.t1905 D.t3545 S.t270 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1906 D.t3544 G.t1906 S.t2700 S.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1907 D.t3404 G.t1907 S.t2699 S.t176 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1908 S.t2698 G.t1908 D.t3403 S.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1909 D.t3402 G.t1909 S.t2697 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1910 S.t2696 G.t1910 D.t3401 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1911 D.t3360 G.t1911 S.t2695 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1912 D.t3359 G.t1912 S.t2694 S.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1913 S.t2693 G.t1913 D.t3358 S.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1914 D.t3357 G.t1914 S.t2692 S.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1915 S.t2691 G.t1915 D.t3984 S.t150 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1916 S.t2690 G.t1916 D.t3983 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1917 D.t3982 G.t1917 S.t2689 S.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1918 D.t3981 G.t1918 S.t2688 S.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1919 S.t2687 G.t1919 D.t3480 S.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1920 D.t3479 G.t1920 S.t2686 S.t158 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1921 S.t2685 G.t1921 D.t3478 S.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1922 S.t2684 G.t1922 D.t3477 S.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1923 S.t2683 G.t1923 D.t3610 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1924 D.t3609 G.t1924 S.t2682 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1925 S.t2681 G.t1925 D.t3608 S.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1926 D.t3607 G.t1926 S.t2680 S.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1927 D.t4049 G.t1927 S.t2679 S.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1928 D.t4048 G.t1928 S.t2678 S.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1929 D.t4047 G.t1929 S.t2677 S.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1930 D.t4046 G.t1930 S.t2676 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1931 S.t2675 G.t1931 D.t3671 S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1932 S.t2674 G.t1932 D.t3670 S.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1933 S.t2673 G.t1933 D.t3669 S.t443 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1934 D.t3668 G.t1934 S.t2672 S.t209 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1935 S.t2671 G.t1935 D.t4053 S.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1936 D.t4052 G.t1936 S.t2670 S.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1937 D.t4051 G.t1937 S.t2669 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1938 S.t2668 G.t1938 D.t4050 S.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1939 D.t3683 G.t1939 S.t2667 S.t357 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1940 S.t2666 G.t1940 D.t3682 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1941 S.t2665 G.t1941 D.t3681 S.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1942 S.t2664 G.t1942 D.t3680 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1943 S.t2663 G.t1943 D.t4142 S.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1944 D.t4141 G.t1944 S.t2662 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1945 S.t2661 G.t1945 D.t4140 S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1946 S.t2660 G.t1946 D.t4139 S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1947 D.t3484 G.t1947 S.t2659 S.t218 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1948 D.t3483 G.t1948 S.t2658 S.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1949 S.t2657 G.t1949 D.t3482 S.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1950 D.t3481 G.t1950 S.t2656 S.t216 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1951 S.t2655 G.t1951 D.t3364 S.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1952 S.t2654 G.t1952 D.t3363 S.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1953 D.t3362 G.t1953 S.t2653 S.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1954 S.t2652 G.t1954 D.t3361 S.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1955 D.t4147 G.t1955 S.t2651 S.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1956 S.t2650 G.t1956 D.t4146 S.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1957 D.t4145 G.t1957 S.t2649 S.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1958 S.t2648 G.t1958 D.t4144 S.t139 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1959 D.t3303 G.t1959 S.t2647 S.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1960 S.t2646 G.t1960 D.t3302 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1961 S.t2645 G.t1961 D.t3301 S.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1962 S.t2644 G.t1962 D.t3300 S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1963 S.t2643 G.t1963 D.t4151 S.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1964 D.t4150 G.t1964 S.t2642 S.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1965 S.t2641 G.t1965 D.t4149 S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1966 S.t2640 G.t1966 D.t4148 S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1967 S.t2639 G.t1967 D.t3679 S.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1968 S.t2638 G.t1968 D.t3678 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1969 D.t3677 G.t1969 S.t2637 S.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1970 S.t2636 G.t1970 D.t3676 S.t406 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1971 S.t2635 G.t1971 D.t3380 S.t198 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1972 D.t3379 G.t1972 S.t2634 S.t176 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1973 S.t2633 G.t1973 D.t3378 S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1974 D.t3377 G.t1974 S.t2632 S.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1975 D.t3408 G.t1975 S.t2631 S.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1976 D.t3407 G.t1976 S.t2630 S.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1977 S.t2629 G.t1977 D.t3406 S.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1978 S.t2628 G.t1978 D.t3405 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1979 D.t3614 G.t1979 S.t2627 S.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1980 S.t2626 G.t1980 D.t3613 S.t332 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1981 S.t2625 G.t1981 D.t3612 S.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1982 S.t2624 G.t1982 D.t3611 S.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1983 D.t3239 G.t1983 S.t2623 S.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1984 S.t2622 G.t1984 D.t3238 S.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1985 S.t2621 G.t1985 D.t3237 S.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1986 D.t3236 G.t1986 S.t2620 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1987 D.t3368 G.t1987 S.t2619 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1988 S.t2618 G.t1988 D.t3367 S.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1989 S.t2617 G.t1989 D.t3366 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1990 S.t2616 G.t1990 D.t3365 S.t198 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1991 S.t2615 G.t1991 D.t3384 S.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1992 S.t2614 G.t1992 D.t3383 S.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1993 D.t3382 G.t1993 S.t2613 S.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1994 S.t2612 G.t1994 D.t3381 S.t332 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1995 S.t2611 G.t1995 D.t3928 S.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1996 D.t3927 G.t1996 S.t2610 S.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1997 D.t3926 G.t1997 S.t2609 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1998 S.t2608 G.t1998 D.t3925 S.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1999 S.t2607 G.t1999 D.t3307 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2000 S.t2606 G.t2000 D.t3306 S.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2001 D.t3305 G.t2001 S.t2605 S.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2002 D.t3304 G.t2002 S.t2604 S.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2003 S.t2603 G.t2003 D.t3675 S.t443 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2004 D.t3674 G.t2004 S.t2602 S.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2005 S.t2601 G.t2005 D.t3673 S.t270 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2006 S.t2600 G.t2006 D.t3672 S.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2007 S.t2599 G.t2007 D.t3865 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2008 D.t3864 G.t2008 S.t2598 S.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2009 D.t3863 G.t2009 S.t2597 S.t388 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2010 D.t3862 G.t2010 S.t2596 S.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2011 S.t2595 G.t2011 D.t3462 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2012 S.t2594 G.t2012 D.t3461 S.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2013 S.t2593 G.t2013 D.t3460 S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2014 S.t2592 G.t2014 D.t3459 S.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2015 D.t3687 G.t2015 S.t2591 S.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2016 D.t3686 G.t2016 S.t2590 S.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2017 D.t3685 G.t2017 S.t2589 S.t357 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2018 S.t2588 G.t2018 D.t3684 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2019 S.t2587 G.t2019 D.t3388 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2020 D.t3387 G.t2020 S.t2586 S.t216 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2021 S.t2585 G.t2021 D.t3386 S.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2022 S.t2584 G.t2022 D.t3385 S.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2023 D.t3392 G.t2023 S.t2583 S.t270 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2024 D.t3391 G.t2024 S.t2582 S.t321 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2025 S.t2581 G.t2025 D.t3390 S.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2026 D.t3389 G.t2026 S.t2580 S.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2027 S.t2579 G.t2027 D.t3372 S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2028 D.t3371 G.t2028 S.t2578 S.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2029 S.t2577 G.t2029 D.t3370 S.t216 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2030 D.t3369 G.t2030 S.t2576 S.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2031 S.t2575 G.t2031 D.t3311 S.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2032 S.t2574 G.t2032 D.t3310 S.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2033 D.t3309 G.t2033 S.t2573 S.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2034 D.t3308 G.t2034 S.t2572 S.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2035 S.t2571 G.t2035 D.t3731 S.t158 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2036 D.t3730 G.t2036 S.t2570 S.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2037 D.t3729 G.t2037 S.t2569 S.t150 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2038 S.t2568 G.t2038 D.t3728 S.t406 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2039 D.t3718 G.t2039 S.t2567 S.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2040 D.t3717 G.t2040 S.t2566 S.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2041 S.t2565 G.t2041 D.t3716 S.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2042 S.t2564 G.t2042 D.t3715 S.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2043 S.t2563 G.t2043 D.t3780 S.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2044 D.t3779 G.t2044 S.t2562 S.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2045 D.t3778 G.t2045 S.t2561 S.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2046 S.t2560 G.t2046 D.t3777 S.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2047 D.t3735 G.t2047 S.t2559 S.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2048 D.t3734 G.t2048 S.t2558 S.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2049 S.t2557 G.t2049 D.t3733 S.t270 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2050 S.t2556 G.t2050 D.t3732 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2051 D.t3722 G.t2051 S.t2555 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2052 S.t2554 G.t2052 D.t3721 S.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2053 S.t2553 G.t2053 D.t3720 S.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2054 S.t2552 G.t2054 D.t3719 S.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2055 D.t3784 G.t2055 S.t2551 S.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2056 D.t3783 G.t2056 S.t2550 S.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2057 S.t2549 G.t2057 D.t3782 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2058 S.t2548 G.t2058 D.t3781 S.t231 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2059 S.t2547 G.t2059 D.t3938 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2060 D.t3937 G.t2060 S.t2546 S.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2061 S.t2545 G.t2061 D.t3936 S.t150 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2062 S.t2544 G.t2062 D.t3935 S.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2063 S.t2543 G.t2063 D.t3551 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2064 S.t2542 G.t2064 D.t3550 S.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2065 S.t2541 G.t2065 D.t3549 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2066 D.t3548 G.t2066 S.t2540 S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2067 S.t2539 G.t2067 D.t3420 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2068 S.t2538 G.t2068 D.t3419 S.t357 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2069 S.t2537 G.t2069 D.t3418 S.t216 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2070 S.t2536 G.t2070 D.t3417 S.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2071 D.t3816 G.t2071 S.t2535 S.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2072 S.t2534 G.t2072 D.t3815 S.t270 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2073 S.t2533 G.t2073 D.t3814 S.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2074 S.t2532 G.t2074 D.t3813 S.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2075 D.t3946 G.t2075 S.t2531 S.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2076 D.t3945 G.t2076 S.t2530 S.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2077 D.t3944 G.t2077 S.t2529 S.t357 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2078 S.t2528 G.t2078 D.t3943 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2079 S.t2527 G.t2079 D.t3833 S.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2080 D.t3832 G.t2080 S.t2526 S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2081 S.t2525 G.t2081 D.t3831 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2082 S.t2524 G.t2082 D.t3830 S.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2083 S.t2523 G.t2083 D.t3820 S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2084 S.t2522 G.t2084 D.t3819 S.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2085 S.t2521 G.t2085 D.t3818 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2086 D.t3817 G.t2086 S.t2520 S.t538 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2087 S.t2519 G.t2087 D.t3559 S.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2088 S.t2518 G.t2088 D.t3558 S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2089 S.t2517 G.t2089 D.t3557 S.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2090 S.t2516 G.t2090 D.t3556 S.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2091 S.t2515 G.t2091 D.t3951 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2092 S.t2514 G.t2092 D.t3950 S.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2093 D.t3949 G.t2093 S.t2513 S.t183 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2094 S.t2512 G.t2094 D.t3948 S.t139 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2095 D.t3698 G.t2095 S.t2511 S.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2096 S.t2510 G.t2096 D.t3697 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2097 D.t3696 G.t2097 S.t2509 S.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2098 D.t3695 G.t2098 S.t2508 S.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2099 S.t2507 G.t2099 D.t3426 S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2100 S.t2506 G.t2100 D.t3425 S.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2101 D.t3424 G.t2101 S.t2505 S.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2102 S.t2504 G.t2102 D.t3423 S.t79 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2103 D.t3873 G.t2103 S.t2503 S.t150 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2104 D.t3872 G.t2104 S.t2502 S.t176 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2105 S.t2501 G.t2105 D.t3871 S.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2106 S.t2500 G.t2106 D.t3870 S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2107 S.t2499 G.t2107 D.t3883 S.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2108 S.t2498 G.t2108 D.t3882 S.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2109 S.t2497 G.t2109 D.t3881 S.t332 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2110 S.t2496 G.t2110 D.t3880 S.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2111 D.t3348 G.t2111 S.t2495 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2112 D.t3347 G.t2112 S.t2494 S.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2113 S.t2493 G.t2113 D.t3346 S.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2114 S.t2492 G.t2114 D.t3345 S.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2115 D.t3976 G.t2115 S.t2491 S.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2116 S.t2490 G.t2116 D.t3975 S.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2117 S.t2489 G.t2117 D.t3974 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2118 S.t2488 G.t2118 D.t3973 S.t198 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2119 D.t3437 G.t2119 S.t2487 S.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2120 S.t2486 G.t2120 D.t3436 S.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2121 D.t3435 G.t2121 S.t2485 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2122 D.t3434 G.t2122 S.t2484 S.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2123 D.t3258 G.t2123 S.t2483 S.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2124 S.t2482 G.t2124 D.t3257 S.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2125 S.t2481 G.t2125 D.t3256 S.t231 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2126 D.t3255 G.t2126 S.t2480 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2127 S.t2479 G.t2127 D.t3341 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2128 D.t3340 G.t2128 S.t2478 S.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2129 D.t3339 G.t2129 S.t2477 S.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2130 D.t3338 G.t2130 S.t2476 S.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2131 S.t2475 G.t2131 D.t3850 S.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2132 D.t3849 G.t2132 S.t2474 S.t388 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2133 D.t3848 G.t2133 S.t2473 S.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2134 D.t3847 G.t2134 S.t2472 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2135 D.t3667 G.t2135 S.t2471 S.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2136 D.t3666 G.t2136 S.t2470 S.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2137 S.t2469 G.t2137 D.t3665 S.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2138 D.t3664 G.t2138 S.t2468 S.t406 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2139 S.t2467 G.t2139 D.t1774 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2140 D.t1773 G.t2140 S.t2466 S.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2141 S.t2465 G.t2141 D.t1772 S.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2142 D.t1771 G.t2142 S.t2464 S.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2143 S.t2463 G.t2143 D.t659 S.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2144 D.t658 G.t2144 S.t2462 S.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2145 S.t2461 G.t2145 D.t657 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2146 S.t2460 G.t2146 D.t656 S.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2147 D.t2592 G.t2147 S.t2459 S.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2148 S.t2458 G.t2148 D.t2591 S.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2149 S.t2457 G.t2149 D.t2590 S.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2150 S.t2456 G.t2150 D.t2589 S.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2151 S.t2455 G.t2151 D.t554 S.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2152 S.t2454 G.t2152 D.t553 S.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2153 S.t2453 G.t2153 D.t552 S.t158 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2154 S.t2452 G.t2154 D.t551 S.t216 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2155 S.t2451 G.t2155 D.t1903 S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2156 S.t2450 G.t2156 D.t1902 S.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2157 D.t1901 G.t2157 S.t2449 S.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2158 D.t1900 G.t2158 S.t2448 S.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2159 D.t1898 G.t2159 S.t2447 S.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2160 D.t1897 G.t2160 S.t2446 S.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2161 S.t2445 G.t2161 D.t1896 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2162 D.t1895 G.t2162 S.t2444 S.t183 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2163 D.t1873 G.t2163 S.t2443 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2164 D.t1872 G.t2164 S.t2442 S.t150 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2165 S.t2441 G.t2165 D.t1871 S.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2166 D.t1870 G.t2166 S.t2440 S.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2167 S.t2439 G.t2167 D.t1865 S.t209 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2168 D.t1864 G.t2168 S.t2438 S.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2169 S.t2437 G.t2169 D.t1863 S.t79 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2170 S.t2436 G.t2170 D.t1862 S.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2171 S.t2435 G.t2171 D.t1857 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2172 D.t1856 G.t2172 S.t2434 S.t538 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2173 S.t2433 G.t2173 D.t1855 S.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2174 D.t1854 G.t2174 S.t2432 S.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2175 D.t1820 G.t2175 S.t2431 S.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2176 D.t1819 G.t2176 S.t2430 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2177 S.t2429 G.t2177 D.t1818 S.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2178 D.t1817 G.t2178 S.t2428 S.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2179 D.t1812 G.t2179 S.t2427 S.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2180 S.t2426 G.t2180 D.t1811 S.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2181 S.t2425 G.t2181 D.t1810 S.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2182 S.t2424 G.t2182 D.t1809 S.t231 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2183 S.t2423 G.t2183 D.t1803 S.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2184 D.t1802 G.t2184 S.t2422 S.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2185 D.t1801 G.t2185 S.t2421 S.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2186 S.t2420 G.t2186 D.t1800 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2187 D.t1540 G.t2187 S.t2419 S.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2188 D.t1539 G.t2188 S.t2418 S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2189 S.t2417 G.t2189 D.t1538 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2190 S.t2416 G.t2190 D.t1537 S.t357 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2191 S.t2415 G.t2191 D.t1554 S.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2192 S.t2414 G.t2192 D.t1553 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2193 D.t1552 G.t2193 S.t2413 S.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2194 S.t2412 G.t2194 D.t1551 S.t216 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2195 S.t2411 G.t2195 D.t640 S.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2196 S.t2410 G.t2196 D.t639 S.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2197 S.t2409 G.t2197 D.t638 S.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2198 D.t637 G.t2198 S.t2408 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2199 D.t383 G.t2199 S.t2407 S.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2200 D.t382 G.t2200 S.t2406 S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2201 S.t2405 G.t2201 D.t381 S.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2202 S.t2404 G.t2202 D.t380 S.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2203 D.t4072 G.t2203 S.t2403 S.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2204 S.t2402 G.t2204 D.t4071 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2205 S.t2401 G.t2205 D.t4070 S.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2206 D.t4069 G.t2206 S.t2400 S.t538 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2207 D.t3647 G.t2207 S.t2399 S.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2208 D.t3646 G.t2208 S.t2398 S.t443 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2209 D.t3645 G.t2209 S.t2397 S.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2210 D.t3644 G.t2210 S.t2396 S.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2211 S.t2395 G.t2211 D.t3630 S.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2212 S.t2394 G.t2212 D.t3629 S.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2213 S.t2393 G.t2213 D.t3628 S.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2214 S.t2392 G.t2214 D.t3627 S.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2215 D.t203 G.t2215 S.t2391 S.t183 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2216 S.t2390 G.t2216 D.t202 S.t158 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2217 S.t2389 G.t2217 D.t201 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2218 S.t2388 G.t2218 D.t200 S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2219 D.t214 G.t2219 S.t2387 S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2220 D.t213 G.t2220 S.t2386 S.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2221 S.t2385 G.t2221 D.t212 S.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2222 S.t2384 G.t2222 D.t211 S.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2223 D.t2150 G.t2223 S.t2383 S.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2224 D.t2149 G.t2224 S.t2382 S.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2225 D.t2148 G.t2225 S.t2381 S.t231 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2226 D.t2147 G.t2226 S.t2380 S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2227 S.t2379 G.t2227 D.t1290 S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2228 D.t1289 G.t2228 S.t2378 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2229 S.t2377 G.t2229 D.t1288 S.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2230 D.t1287 G.t2230 S.t2376 S.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2231 D.t1272 G.t2231 S.t2375 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2232 S.t2374 G.t2232 D.t1271 S.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2233 S.t2373 G.t2233 D.t1270 S.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2234 D.t1269 G.t2234 S.t2372 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2235 D.t1250 G.t2235 S.t2371 S.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2236 D.t1249 G.t2236 S.t2370 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2237 S.t2369 G.t2237 D.t1248 S.t209 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2238 D.t1247 G.t2238 S.t2368 S.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2239 S.t2367 G.t2239 D.t1206 S.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2240 S.t2366 G.t2240 D.t1205 S.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2241 D.t1204 G.t2241 S.t2365 S.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2242 D.t1203 G.t2242 S.t2364 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2243 D.t1177 G.t2243 S.t2363 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2244 D.t1176 G.t2244 S.t2362 S.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2245 D.t1175 G.t2245 S.t2361 S.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2246 D.t1174 G.t2246 S.t2360 S.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2247 D.t974 G.t2247 S.t2359 S.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2248 D.t973 G.t2248 S.t2358 S.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2249 D.t972 G.t2249 S.t2357 S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2250 S.t2356 G.t2250 D.t971 S.t218 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2251 D.t967 G.t2251 S.t2355 S.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2252 D.t966 G.t2252 S.t2354 S.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2253 S.t2353 G.t2253 D.t965 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2254 S.t2352 G.t2254 D.t964 S.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2255 D.t832 G.t2255 S.t2351 S.t406 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2256 S.t2350 G.t2256 D.t831 S.t183 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2257 D.t830 G.t2257 S.t2349 S.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2258 S.t2348 G.t2258 D.t829 S.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2259 D.t473 G.t2259 S.t2347 S.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2260 D.t472 G.t2260 S.t2346 S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2261 S.t2345 G.t2261 D.t471 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2262 S.t2344 G.t2262 D.t470 S.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2263 D.t1310 G.t2263 S.t2343 S.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2264 D.t1309 G.t2264 S.t2342 S.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2265 D.t1308 G.t2265 S.t2341 S.t79 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2266 S.t2340 G.t2266 D.t1307 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2267 S.t2339 G.t2267 D.t1998 S.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2268 S.t2338 G.t2268 D.t1997 S.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2269 D.t1996 G.t2269 S.t2337 S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2270 S.t2336 G.t2270 D.t1995 S.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2271 S.t2335 G.t2271 D.t1604 S.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2272 D.t1603 G.t2272 S.t2334 S.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2273 D.t1602 G.t2273 S.t2333 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2274 S.t2332 G.t2274 D.t1601 S.t321 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2275 S.t2331 G.t2275 D.t1123 S.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2276 D.t1122 G.t2276 S.t2330 S.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2277 D.t1121 G.t2277 S.t2329 S.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2278 D.t1120 G.t2278 S.t2328 S.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2279 S.t2327 G.t2279 D.t336 S.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2280 D.t335 G.t2280 S.t2326 S.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2281 S.t2325 G.t2281 D.t334 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2282 D.t333 G.t2282 S.t2324 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2283 D.t252 G.t2283 S.t2323 S.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2284 D.t251 G.t2284 S.t2322 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2285 D.t250 G.t2285 S.t2321 S.t406 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2286 D.t249 G.t2286 S.t2320 S.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2287 D.t3956 G.t2287 S.t2319 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2288 D.t3955 G.t2288 S.t2318 S.t357 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2289 S.t2317 G.t2289 D.t3954 S.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2290 D.t3953 G.t2290 S.t2316 S.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2291 D.t3250 G.t2291 S.t2315 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2292 S.t2314 G.t2292 D.t3249 S.t388 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2293 D.t3248 G.t2293 S.t2313 S.t538 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2294 S.t2312 G.t2294 D.t3247 S.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2295 S.t2311 G.t2295 D.t3600 S.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2296 S.t2310 G.t2296 D.t3599 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2297 D.t3598 G.t2297 S.t2309 S.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2298 S.t2308 G.t2298 D.t3597 S.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2299 S.t2307 G.t2299 D.t3280 S.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2300 S.t2306 G.t2300 D.t3279 S.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2301 D.t3278 G.t2301 S.t2305 S.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2302 S.t2304 G.t2302 D.t3277 S.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2303 D.t3593 G.t2303 S.t2303 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2304 D.t3592 G.t2304 S.t2302 S.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2305 S.t2301 G.t2305 D.t3591 S.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2306 S.t2300 G.t2306 D.t3590 S.t231 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2307 D.t3651 G.t2307 S.t2299 S.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2308 D.t3650 G.t2308 S.t2298 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2309 S.t2297 G.t2309 D.t3649 S.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2310 D.t3648 G.t2310 S.t2296 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2311 S.t2295 G.t2311 D.t1493 S.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2312 S.t2294 G.t2312 D.t1492 S.t538 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2313 S.t2293 G.t2313 D.t1491 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2314 D.t1490 G.t2314 S.t2292 S.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2315 S.t2291 G.t2315 D.t1489 S.t357 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2316 D.t1488 G.t2316 S.t2290 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2317 D.t1487 G.t2317 S.t2289 S.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2318 D.t1486 G.t2318 S.t2288 S.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2319 S.t2287 G.t2319 D.t1477 S.t216 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2320 D.t1476 G.t2320 S.t2286 S.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2321 D.t1475 G.t2321 S.t2285 S.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2322 S.t2284 G.t2322 D.t1474 S.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2323 D.t1473 G.t2323 S.t2283 S.t158 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2324 S.t2282 G.t2324 D.t1472 S.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2325 D.t1471 G.t2325 S.t2281 S.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2326 D.t1470 G.t2326 S.t2280 S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2327 S.t2279 G.t2327 D.t1461 S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2328 S.t2278 G.t2328 D.t1460 S.t357 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2329 D.t1459 G.t2329 S.t2277 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2330 S.t2276 G.t2330 D.t1458 S.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2331 S.t2275 G.t2331 D.t1457 S.t388 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2332 D.t1456 G.t2332 S.t2274 S.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2333 S.t2273 G.t2333 D.t1455 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2334 S.t2272 G.t2334 D.t1454 S.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2335 S.t2271 G.t2335 D.t1445 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2336 D.t1444 G.t2336 S.t2270 S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2337 D.t1443 G.t2337 S.t2269 S.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2338 D.t1442 G.t2338 S.t2268 S.t198 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2339 D.t1441 G.t2339 S.t2267 S.t538 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2340 S.t2266 G.t2340 D.t1440 S.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2341 D.t1439 G.t2341 S.t2265 S.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2342 S.t2264 G.t2342 D.t1438 S.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2343 D.t1429 G.t2343 S.t2263 S.t443 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2344 S.t2262 G.t2344 D.t1428 S.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2345 D.t1427 G.t2345 S.t2261 S.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2346 S.t2260 G.t2346 D.t1426 S.t231 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2347 S.t2259 G.t2347 D.t1425 S.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2348 S.t2258 G.t2348 D.t1424 S.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2349 S.t2257 G.t2349 D.t1423 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2350 D.t1422 G.t2350 S.t2256 S.t139 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2351 D.t1413 G.t2351 S.t2255 S.t270 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2352 D.t1412 G.t2352 S.t2254 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2353 S.t2253 G.t2353 D.t1411 S.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2354 D.t1410 G.t2354 S.t2252 S.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2355 S.t2251 G.t2355 D.t1409 S.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2356 S.t2250 G.t2356 D.t1408 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2357 D.t1407 G.t2357 S.t2249 S.t332 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2358 D.t1406 G.t2358 S.t2248 S.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2359 S.t2247 G.t2359 D.t481 S.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2360 D.t480 G.t2360 S.t2246 S.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2361 D.t479 G.t2361 S.t2245 S.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2362 D.t478 G.t2362 S.t2244 S.t231 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2363 D.t464 G.t2363 S.t2243 S.t406 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2364 S.t2242 G.t2364 D.t463 S.t321 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2365 D.t462 G.t2365 S.t2241 S.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2366 D.t461 G.t2366 S.t2240 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2367 S.t2239 G.t2367 D.t593 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2368 S.t2238 G.t2368 D.t592 S.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2369 D.t591 G.t2369 S.t2237 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2370 D.t590 G.t2370 S.t2236 S.t357 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2371 D.t1629 G.t2371 S.t2235 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2372 S.t2234 G.t2372 D.t1628 S.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2373 S.t2233 G.t2373 D.t1627 S.t388 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2374 D.t1626 G.t2374 S.t2232 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2375 S.t2231 G.t2375 D.t620 S.t209 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2376 D.t619 G.t2376 S.t2230 S.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2377 D.t618 G.t2377 S.t2229 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2378 S.t2228 G.t2378 D.t617 S.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2379 D.t999 G.t2379 S.t2227 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2380 S.t2226 G.t2380 D.t998 S.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2381 D.t997 G.t2381 S.t2225 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2382 D.t996 G.t2382 S.t2224 S.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2383 D.t432 G.t2383 S.t2223 S.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2384 S.t2222 G.t2384 D.t431 S.t231 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2385 D.t430 G.t2385 S.t2221 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2386 D.t429 G.t2386 S.t2220 S.t443 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2387 D.t2552 G.t2387 S.t2219 S.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2388 S.t2218 G.t2388 D.t2551 S.t538 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2389 D.t2550 G.t2389 S.t2217 S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2390 D.t2549 G.t2390 S.t2216 S.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2391 S.t2215 G.t2391 D.t3192 S.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2392 D.t3191 G.t2392 S.t2214 S.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2393 S.t2213 G.t2393 D.t3190 S.t218 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2394 S.t2212 G.t2394 D.t3189 S.t388 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2395 D.t1738 G.t2395 S.t2211 S.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2396 D.t1737 G.t2396 S.t2210 S.t406 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2397 D.t1736 G.t2397 S.t2209 S.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2398 S.t2208 G.t2398 D.t1735 S.t183 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2399 S.t2207 G.t2399 D.t2003 S.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2400 D.t2002 G.t2400 S.t2206 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2401 D.t2001 G.t2401 S.t2205 S.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2402 D.t2000 G.t2402 S.t2204 S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2403 D.t1879 G.t2403 S.t2203 S.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2404 S.t2202 G.t2404 D.t1878 S.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2405 S.t2201 G.t2405 D.t1877 S.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2406 S.t2200 G.t2406 D.t1876 S.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2407 S.t2199 G.t2407 D.t1650 S.t357 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2408 S.t2198 G.t2408 D.t1649 S.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2409 D.t1648 G.t2409 S.t2197 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2410 S.t2196 G.t2410 D.t1647 S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2411 D.t1574 G.t2411 S.t2195 S.t79 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2412 S.t2194 G.t2412 D.t1573 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2413 S.t2193 G.t2413 D.t1572 S.t538 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2414 D.t1571 G.t2414 S.t2192 S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2415 D.t787 G.t2415 S.t2191 S.t198 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2416 S.t2190 G.t2416 D.t786 S.t176 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2417 D.t785 G.t2417 S.t2189 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2418 D.t784 G.t2418 S.t2188 S.t321 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2419 S.t2187 G.t2419 D.t783 S.t321 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2420 S.t2186 G.t2420 D.t782 S.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2421 S.t2185 G.t2421 D.t781 S.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2422 S.t2184 G.t2422 D.t780 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2423 S.t2183 G.t2423 D.t744 S.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2424 S.t2182 G.t2424 D.t743 S.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2425 D.t742 G.t2425 S.t2181 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2426 D.t741 G.t2426 S.t2180 S.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2427 S.t2179 G.t2427 D.t343 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2428 S.t2178 G.t2428 D.t342 S.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2429 S.t2177 G.t2429 D.t341 S.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2430 S.t2176 G.t2430 D.t340 S.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2431 D.t911 G.t2431 S.t2175 S.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2432 S.t2174 G.t2432 D.t910 S.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2433 S.t2173 G.t2433 D.t909 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2434 D.t908 G.t2434 S.t2172 S.t332 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2435 D.t886 G.t2435 S.t2171 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2436 S.t2170 G.t2436 D.t885 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2437 S.t2169 G.t2437 D.t884 S.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2438 S.t2168 G.t2438 D.t883 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2439 S.t2167 G.t2439 D.t1243 S.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2440 D.t1242 G.t2440 S.t2166 S.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2441 S.t2165 G.t2441 D.t1241 S.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2442 S.t2164 G.t2442 D.t1240 S.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2443 S.t2163 G.t2443 D.t1220 S.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2444 S.t2162 G.t2444 D.t1219 S.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2445 S.t2161 G.t2445 D.t1218 S.t388 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2446 D.t1217 G.t2446 S.t2160 S.t538 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2447 S.t2159 G.t2447 D.t926 S.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2448 S.t2158 G.t2448 D.t925 S.t321 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2449 S.t2157 G.t2449 D.t924 S.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2450 D.t923 G.t2450 S.t2156 S.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2451 S.t2155 G.t2451 D.t899 S.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2452 D.t898 G.t2452 S.t2154 S.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2453 S.t2153 G.t2453 D.t897 S.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2454 S.t2152 G.t2454 D.t896 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2455 D.t873 G.t2455 S.t2151 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2456 S.t2150 G.t2456 D.t872 S.t406 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2457 S.t2149 G.t2457 D.t871 S.t231 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2458 D.t870 G.t2458 S.t2148 S.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2459 S.t2147 G.t2459 D.t866 S.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2460 D.t865 G.t2460 S.t2146 S.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2461 S.t2145 G.t2461 D.t864 S.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2462 D.t863 G.t2462 S.t2144 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2463 S.t2143 G.t2463 D.t851 S.t538 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2464 D.t850 G.t2464 S.t2142 S.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2465 S.t2141 G.t2465 D.t849 S.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2466 S.t2140 G.t2466 D.t848 S.t443 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2467 D.t818 G.t2467 S.t2139 S.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2468 D.t817 G.t2468 S.t2138 S.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2469 D.t816 G.t2469 S.t2137 S.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2470 D.t815 G.t2470 S.t2136 S.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2471 S.t2135 G.t2471 D.t390 S.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2472 D.t389 G.t2472 S.t2134 S.t443 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2473 S.t2133 G.t2473 D.t388 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2474 D.t387 G.t2474 S.t2132 S.t158 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2475 D.t3376 G.t2475 S.t2131 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2476 S.t2130 G.t2476 D.t3375 S.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2477 S.t2129 G.t2477 D.t3374 S.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2478 D.t3373 G.t2478 S.t2128 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2479 S.t2127 G.t2479 D.t3543 S.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2480 D.t3542 G.t2480 S.t2126 S.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2481 D.t3541 G.t2481 S.t2125 S.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2482 S.t2124 G.t2482 D.t3540 S.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2483 S.t2123 G.t2483 D.t3412 S.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2484 S.t2122 G.t2484 D.t3411 S.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2485 D.t3410 G.t2485 S.t2121 S.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2486 S.t2120 G.t2486 D.t3409 S.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2487 S.t2119 G.t2487 D.t3491 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2488 D.t3490 G.t2488 S.t2118 S.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2489 D.t3489 G.t2489 S.t2117 S.t198 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2490 D.t3488 G.t2490 S.t2116 S.t218 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2491 D.t2517 G.t2491 S.t2115 S.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2492 S.t2114 G.t2492 D.t2516 S.t406 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2493 D.t2515 G.t2493 S.t2113 S.t443 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2494 S.t2112 G.t2494 D.t2514 S.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2495 D.t2296 G.t2495 S.t2111 S.t183 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2496 S.t2110 G.t2496 D.t2295 S.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2497 S.t2109 G.t2497 D.t2294 S.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2498 S.t2108 G.t2498 D.t2293 S.t332 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2499 D.t3182 G.t2499 S.t2107 S.t388 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2500 S.t2106 G.t2500 D.t3181 S.t538 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2501 D.t3180 G.t2501 S.t2105 S.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2502 D.t3179 G.t2502 S.t2104 S.t270 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2503 D.t1715 G.t2503 S.t2103 S.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2504 D.t1714 G.t2504 S.t2102 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2505 D.t1713 G.t2505 S.t2101 S.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2506 S.t2100 G.t2506 D.t813 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2507 S.t2099 G.t2507 D.t812 S.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2508 D.t811 G.t2508 S.t2098 S.t209 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2509 D.t1924 G.t2509 S.t2097 S.t332 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2510 D.t1923 G.t2510 S.t2096 S.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2511 S.t2095 G.t2511 D.t1922 S.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2512 S.t2094 G.t2512 D.t1921 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2513 D.t1920 G.t2513 S.t2093 S.t231 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2514 S.t2092 G.t2514 D.t1919 S.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2515 D.t1894 G.t2515 S.t2091 S.t231 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2516 S.t2090 G.t2516 D.t1893 S.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2517 D.t1892 G.t2517 S.t2089 S.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2518 S.t2088 G.t2518 D.t600 S.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2519 S.t2087 G.t2519 D.t599 S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2520 D.t598 G.t2520 S.t2086 S.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2521 S.t2085 G.t2521 D.t458 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2522 D.t457 G.t2522 S.t2084 S.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2523 S.t2083 G.t2523 D.t456 S.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2524 D.t442 G.t2524 S.t2082 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2525 D.t441 G.t2525 S.t2081 S.t218 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2526 S.t2080 G.t2526 D.t440 S.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2527 D.t869 G.t2527 S.t2079 S.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2528 S.t2078 G.t2528 D.t868 S.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2529 D.t867 G.t2529 S.t2077 S.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2530 S.t2076 G.t2530 D.t1260 S.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2531 S.t2075 G.t2531 D.t1259 S.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2532 S.t2074 G.t2532 D.t1258 S.t406 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2533 D.t1235 G.t2533 S.t2073 S.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2534 S.t2072 G.t2534 D.t1234 S.t209 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2535 D.t1233 G.t2535 S.t2071 S.t183 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2536 D.t1229 G.t2536 S.t2070 S.t139 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2537 S.t2069 G.t2537 D.t1228 S.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2538 D.t1227 G.t2538 S.t2068 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2539 D.t1189 G.t2539 S.t2067 S.t357 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2540 S.t2066 G.t2540 D.t1188 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2541 S.t2065 G.t2541 D.t1187 S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2542 D.t199 G.t2542 S.t2064 S.t357 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2543 D.t198 G.t2543 S.t2063 S.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2544 S.t2062 G.t2544 D.t197 S.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2545 D.t2513 G.t2545 S.t2061 S.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2546 D.t2512 G.t2546 S.t2060 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2547 S.t2059 G.t2547 D.t2511 S.t198 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2548 D.t2510 G.t2548 S.t2058 S.t176 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2549 D.t2509 G.t2549 S.t2057 S.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2550 S.t2056 G.t2550 D.t2508 S.t443 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2551 D.t2507 G.t2551 S.t2055 S.t321 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2552 S.t2054 G.t2552 D.t2506 S.t218 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2553 D.t2505 G.t2553 S.t2053 S.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2554 S.t2052 G.t2554 D.t2504 S.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2555 D.t2503 G.t2555 S.t2051 S.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2556 D.t2502 G.t2556 S.t2050 S.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2557 D.t2501 G.t2557 S.t2049 S.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2558 S.t2048 G.t2558 D.t2500 S.t183 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2559 D.t2499 G.t2559 S.t2047 S.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2560 D.t2498 G.t2560 S.t2046 S.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2561 S.t2045 G.t2561 D.t2497 S.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2562 S.t2044 G.t2562 D.t2496 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2563 D.t2495 G.t2563 S.t2043 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2564 S.t2042 G.t2564 D.t2494 S.t139 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2565 S.t2041 G.t2565 D.t2493 S.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2566 S.t2040 G.t2566 D.t2492 S.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2567 D.t2491 G.t2567 S.t2039 S.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2568 S.t2038 G.t2568 D.t2490 S.t332 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2569 D.t2489 G.t2569 S.t2037 S.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2570 S.t2036 G.t2570 D.t2488 S.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2571 D.t2487 G.t2571 S.t2035 S.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2572 S.t2034 G.t2572 D.t2486 S.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2573 S.t2033 G.t2573 D.t2485 S.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2574 S.t2032 G.t2574 D.t2484 S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2575 S.t2031 G.t2575 D.t2483 S.t176 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2576 S.t2030 G.t2576 D.t2482 S.t538 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2577 D.t2481 G.t2577 S.t2029 S.t321 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2578 D.t2480 G.t2578 S.t2028 S.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2579 S.t2027 G.t2579 D.t2479 S.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2580 S.t2026 G.t2580 D.t2478 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2581 D.t2477 G.t2581 S.t2025 S.t183 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2582 S.t2024 G.t2582 D.t2476 S.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2583 D.t2475 G.t2583 S.t2023 S.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2584 S.t2022 G.t2584 D.t2474 S.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2585 S.t2021 G.t2585 D.t2473 S.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2586 D.t2472 G.t2586 S.t2020 S.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2587 D.t2471 G.t2587 S.t2019 S.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2588 S.t2018 G.t2588 D.t2470 S.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2589 S.t2017 G.t2589 D.t2469 S.t150 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2590 D.t2468 G.t2590 S.t2016 S.t209 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2591 S.t2015 G.t2591 D.t2467 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2592 S.t2014 G.t2592 D.t2466 S.t139 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2593 S.t2013 G.t2593 D.t2465 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2594 D.t2464 G.t2594 S.t2012 S.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2595 S.t2011 G.t2595 D.t2463 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2596 S.t2010 G.t2596 D.t2462 S.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2597 D.t2461 G.t2597 S.t2009 S.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2598 D.t2460 G.t2598 S.t2008 S.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2599 S.t2007 G.t2599 D.t2459 S.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2600 S.t2006 G.t2600 D.t2458 S.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2601 S.t2005 G.t2601 D.t2457 S.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2602 S.t2004 G.t2602 D.t696 S.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2603 D.t695 G.t2603 S.t2003 S.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2604 S.t2002 G.t2604 D.t694 S.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2605 D.t2385 G.t2605 S.t2001 S.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2606 D.t2384 G.t2606 S.t2000 S.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2607 S.t1999 G.t2607 D.t2383 S.t443 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2608 D.t1351 G.t2608 S.t1998 S.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2609 D.t1350 G.t2609 S.t1997 S.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2610 S.t1996 G.t2610 D.t1349 S.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2611 D.t1654 G.t2611 S.t1995 S.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2612 D.t1653 G.t2612 S.t1994 S.t218 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2613 S.t1993 G.t2613 D.t1652 S.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2614 D.t2143 G.t2614 S.t1992 S.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2615 D.t2142 G.t2615 S.t1991 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2616 D.t2141 G.t2616 S.t1990 S.t388 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2617 S.t1989 G.t2617 D.t1808 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2618 S.t1988 G.t2618 D.t1807 S.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2619 D.t1806 G.t2619 S.t1987 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2620 S.t1986 G.t2620 D.t1832 S.t406 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2621 S.t1985 G.t2621 D.t1831 S.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2622 D.t1830 G.t2622 S.t1984 S.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2623 S.t1983 G.t2623 D.t2037 S.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2624 D.t2036 G.t2624 S.t1982 S.t139 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2625 S.t1981 G.t2625 D.t2035 S.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2626 D.t1849 G.t2626 S.t1980 S.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2627 D.t1848 G.t2627 S.t1979 S.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2628 D.t1847 G.t2628 S.t1978 S.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2629 D.t1842 G.t2629 S.t1977 S.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2630 S.t1976 G.t2630 D.t1841 S.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2631 D.t1840 G.t2631 S.t1975 S.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2632 D.t1835 G.t2632 S.t1974 S.t216 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2633 D.t1834 G.t2633 S.t1973 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2634 D.t1833 G.t2634 S.t1972 S.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2635 S.t1971 G.t2635 D.t1827 S.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2636 D.t1826 G.t2636 S.t1970 S.t321 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2637 D.t1825 G.t2637 S.t1969 S.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2638 S.t1968 G.t2638 D.t1480 S.t270 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2639 D.t1479 G.t2639 S.t1967 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2640 S.t1966 G.t2640 D.t1478 S.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2641 D.t1464 G.t2641 S.t1965 S.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2642 D.t1463 G.t2642 S.t1964 S.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2643 S.t1963 G.t2643 D.t1462 S.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2644 D.t1448 G.t2644 S.t1962 S.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2645 S.t1961 G.t2645 D.t1447 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2646 S.t1960 G.t2646 D.t1446 S.t406 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2647 S.t1959 G.t2647 D.t1432 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2648 D.t1431 G.t2648 S.t1958 S.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2649 S.t1957 G.t2649 D.t1430 S.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2650 D.t1416 G.t2650 S.t1956 S.t183 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2651 D.t1415 G.t2651 S.t1955 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2652 S.t1954 G.t2652 D.t1414 S.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2653 D.t1400 G.t2653 S.t1953 S.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2654 S.t1952 G.t2654 D.t1399 S.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2655 D.t1398 G.t2655 S.t1951 S.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2656 S.t1950 G.t2656 D.t1333 S.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2657 D.t1332 G.t2657 S.t1949 S.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2658 D.t1331 G.t2658 S.t1948 S.t388 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2659 D.t1303 G.t2659 S.t1947 S.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2660 D.t1302 G.t2660 S.t1946 S.t270 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2661 S.t1945 G.t2661 D.t1301 S.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2662 D.t994 G.t2662 S.t1944 S.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2663 D.t993 G.t2663 S.t1943 S.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2664 D.t992 G.t2664 S.t1942 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2665 D.t379 G.t2665 S.t1941 S.t209 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2666 D.t378 G.t2666 S.t1940 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2667 S.t1939 G.t2667 D.t377 S.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2668 S.t1938 G.t2668 D.t526 S.t538 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2669 S.t1937 G.t2669 D.t525 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2670 D.t524 G.t2670 S.t1936 S.t231 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2671 S.t1935 G.t2671 D.t894 S.t150 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2672 S.t1934 G.t2672 D.t893 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2673 D.t892 G.t2673 S.t1933 S.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2674 S.t1932 G.t2674 D.t636 S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2675 D.t635 G.t2675 S.t1931 S.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2676 D.t634 G.t2676 S.t1930 S.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2677 S.t1929 G.t2677 D.t963 S.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2678 S.t1928 G.t2678 D.t962 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2679 D.t961 G.t2679 S.t1927 S.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2680 D.t374 G.t2680 S.t1926 S.t218 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2681 S.t1925 G.t2681 D.t373 S.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2682 D.t372 G.t2682 S.t1924 S.t388 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2683 D.t688 G.t2683 S.t1923 S.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2684 S.t1922 G.t2684 D.t687 S.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2685 D.t686 G.t2685 S.t1921 S.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2686 D.t435 G.t2686 S.t1920 S.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2687 D.t434 G.t2687 S.t1919 S.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2688 S.t1918 G.t2688 D.t433 S.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2689 D.t3846 G.t2689 S.t1917 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2690 D.t3845 G.t2690 S.t1916 S.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2691 D.t3844 G.t2691 S.t1915 S.t357 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2692 S.t1914 G.t2692 D.t3824 S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2693 S.t1913 G.t2693 D.t3823 S.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2694 S.t1912 G.t2694 D.t3822 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2695 S.t1911 G.t2695 D.t3877 S.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2696 S.t1910 G.t2696 D.t3876 S.t198 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2697 D.t3875 G.t2697 S.t1909 S.t176 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2698 D.t3886 G.t2698 S.t1908 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2699 D.t3885 G.t2699 S.t1907 S.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2700 D.t3884 G.t2700 S.t1906 S.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2701 S.t1905 G.t2701 D.t3554 S.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2702 D.t3553 G.t2702 S.t1904 S.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2703 S.t1903 G.t2703 D.t3552 S.t183 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2704 D.t3528 G.t2704 S.t1902 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2705 D.t3527 G.t2705 S.t1901 S.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2706 D.t3526 G.t2706 S.t1900 S.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2707 D.t3842 G.t2707 S.t1899 S.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2708 S.t1898 G.t2708 D.t3841 S.t270 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2709 S.t1897 G.t2709 D.t3840 S.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2710 D.t3804 G.t2710 S.t1896 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2711 S.t1895 G.t2711 D.t3803 S.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2712 D.t3802 G.t2712 S.t1894 S.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2713 S.t1893 G.t2713 D.t3807 S.t139 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2714 S.t1892 G.t2714 D.t3806 S.t332 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2715 D.t3805 G.t2715 S.t1891 S.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2716 D.t232 G.t2716 S.t1890 S.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2717 D.t231 G.t2717 S.t1889 S.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2718 D.t230 G.t2718 S.t1888 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2719 S.t1887 G.t2719 D.t229 S.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2720 D.t228 G.t2720 S.t1886 S.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2721 S.t1885 G.t2721 D.t227 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2722 S.t1884 G.t2722 D.t225 S.t176 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2723 S.t1883 G.t2723 D.t224 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2724 D.t223 G.t2724 S.t1882 S.t321 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2725 D.t218 G.t2725 S.t1881 S.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2726 S.t1880 G.t2726 D.t217 S.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2727 D.t216 G.t2727 S.t1879 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2728 S.t1878 G.t2728 D.t282 S.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2729 D.t281 G.t2729 S.t1877 S.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2730 S.t1876 G.t2730 D.t280 S.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2731 S.t1875 G.t2731 D.t23 S.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2732 D.t22 G.t2732 S.t1874 S.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2733 D.t21 G.t2733 S.t1873 S.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2734 S.t1872 G.t2734 D.t1112 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2735 D.t1111 G.t2735 S.t1871 S.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2736 S.t1870 G.t2736 D.t1110 S.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2737 S.t1869 G.t2737 D.t1107 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2738 D.t1106 G.t2738 S.t1868 S.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2739 S.t1867 G.t2739 D.t1105 S.t139 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2740 D.t1102 G.t2740 S.t1866 S.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2741 S.t1865 G.t2741 D.t1101 S.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2742 S.t1864 G.t2742 D.t1100 S.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2743 S.t1863 G.t2743 D.t1097 S.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2744 D.t1096 G.t2744 S.t1862 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2745 D.t1095 G.t2745 S.t1861 S.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2746 S.t1860 G.t2746 D.t1093 S.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2747 S.t1859 G.t2747 D.t1092 S.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2748 D.t1091 G.t2748 S.t1858 S.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2749 S.t1857 G.t2749 D.t1088 S.t443 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2750 D.t1087 G.t2750 S.t1856 S.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2751 D.t1086 G.t2751 S.t1855 S.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2752 S.t1854 G.t2752 D.t1083 S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2753 D.t1082 G.t2753 S.t1853 S.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2754 S.t1852 G.t2754 D.t1081 S.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2755 D.t1080 G.t2755 S.t1851 S.t388 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2756 D.t1079 G.t2756 S.t1850 S.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2757 S.t1849 G.t2757 D.t1078 S.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2758 S.t1848 G.t2758 D.t1075 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2759 D.t1074 G.t2759 S.t1847 S.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2760 D.t1073 G.t2760 S.t1846 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2761 D.t1070 G.t2761 S.t1845 S.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2762 D.t1069 G.t2762 S.t1844 S.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2763 D.t1068 G.t2763 S.t1843 S.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2764 S.t1842 G.t2764 D.t1067 S.t79 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2765 D.t1066 G.t2765 S.t1841 S.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2766 S.t1840 G.t2766 D.t1065 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2767 D.t1062 G.t2767 S.t1839 S.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2768 D.t1061 G.t2768 S.t1838 S.t216 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2769 D.t1060 G.t2769 S.t1837 S.t176 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2770 D.t2333 G.t2770 S.t1836 S.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2771 S.t1835 G.t2771 D.t2332 S.t270 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2772 S.t1834 G.t2772 D.t2331 S.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2773 D.t2453 G.t2773 S.t1833 S.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2774 S.t1832 G.t2774 D.t2452 S.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2775 D.t2451 G.t2775 S.t1831 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2776 S.t1830 G.t2776 D.t2424 S.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2777 S.t1829 G.t2777 D.t2423 S.t79 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2778 S.t1828 G.t2778 D.t2422 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2779 D.t2220 G.t2779 S.t1827 S.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2780 D.t2219 G.t2780 S.t1826 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2781 D.t2218 G.t2781 S.t1825 S.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2782 S.t1824 G.t2782 D.t1660 S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2783 D.t1659 G.t2783 S.t1823 S.t150 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2784 S.t1822 G.t2784 D.t1658 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2785 S.t1821 G.t2785 D.t1890 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2786 D.t1889 G.t2786 S.t1820 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2787 S.t1819 G.t2787 D.t1888 S.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2788 D.t1886 G.t2788 S.t1818 S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2789 S.t1817 G.t2789 D.t1885 S.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2790 D.t1884 G.t2790 S.t1816 S.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2791 S.t1815 G.t2791 D.t1632 S.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2792 D.t1631 G.t2792 S.t1814 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2793 D.t1630 G.t2793 S.t1813 S.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2794 S.t1812 G.t2794 D.t1354 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2795 D.t1353 G.t2795 S.t1811 S.t388 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2796 D.t1352 G.t2796 S.t1810 S.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2797 D.t670 G.t2797 S.t1809 S.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2798 D.t669 G.t2798 S.t1808 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2799 D.t668 G.t2799 S.t1807 S.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2800 S.t1806 G.t2800 D.t499 S.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2801 S.t1805 G.t2801 D.t498 S.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2802 D.t497 G.t2802 S.t1804 S.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2803 D.t291 G.t2803 S.t1803 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2804 D.t290 G.t2804 S.t1802 S.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2805 S.t1801 G.t2805 D.t289 S.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2806 D.t162 G.t2806 S.t1800 S.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2807 S.t1799 G.t2807 D.t161 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2808 D.t160 G.t2808 S.t1798 S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2809 D.t183 G.t2809 S.t1797 S.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2810 S.t1796 G.t2810 D.t182 S.t231 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2811 S.t1795 G.t2811 D.t181 S.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2812 D.t285 G.t2812 S.t1794 S.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2813 D.t284 G.t2813 S.t1793 S.t231 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2814 D.t283 G.t2814 S.t1792 S.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2815 S.t1791 G.t2815 D.t3186 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2816 S.t1790 G.t2816 D.t3185 S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2817 S.t1789 G.t2817 D.t3184 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2818 D.t2618 G.t2818 S.t1788 S.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2819 S.t1787 G.t2819 D.t2617 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2820 D.t2616 G.t2820 S.t1786 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2821 S.t1785 G.t2821 D.t662 S.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2822 S.t1784 G.t2822 D.t661 S.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2823 S.t1783 G.t2823 D.t660 S.t218 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2824 S.t1782 G.t2824 D.t2439 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2825 D.t2438 G.t2825 S.t1781 S.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2826 D.t2437 G.t2826 S.t1780 S.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2827 S.t1779 G.t2827 D.t2436 S.t158 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2828 S.t1778 G.t2828 D.t2435 S.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2829 S.t1777 G.t2829 D.t2434 S.t209 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2830 S.t1776 G.t2830 D.t2433 S.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2831 S.t1775 G.t2831 D.t2432 S.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2832 D.t2431 G.t2832 S.t1774 S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2833 S.t1773 G.t2833 D.t2430 S.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2834 S.t1772 G.t2834 D.t2429 S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2835 D.t2428 G.t2835 S.t1771 S.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2836 S.t1770 G.t2836 D.t2421 S.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2837 S.t1769 G.t2837 D.t2420 S.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2838 S.t1768 G.t2838 D.t2419 S.t198 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2839 D.t2418 G.t2839 S.t1767 S.t176 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2840 D.t2417 G.t2840 S.t1766 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2841 S.t1765 G.t2841 D.t2416 S.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2842 S.t1764 G.t2842 D.t2413 S.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2843 D.t2412 G.t2843 S.t1763 S.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2844 S.t1762 G.t2844 D.t2411 S.t183 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2845 D.t2405 G.t2845 S.t1761 S.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2846 S.t1760 G.t2846 D.t2404 S.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2847 D.t2403 G.t2847 S.t1759 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2848 S.t1758 G.t2848 D.t2402 S.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2849 D.t2401 G.t2849 S.t1757 S.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2850 S.t1756 G.t2850 D.t2400 S.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2851 D.t2396 G.t2851 S.t1755 S.t183 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2852 D.t2395 G.t2852 S.t1754 S.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2853 D.t2394 G.t2853 S.t1753 S.t231 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2854 S.t1752 G.t2854 D.t2393 S.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2855 S.t1751 G.t2855 D.t2392 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2856 S.t1750 G.t2856 D.t2391 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2857 D.t2390 G.t2857 S.t1749 S.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2858 D.t2389 G.t2858 S.t1748 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2859 D.t2388 G.t2859 S.t1747 S.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2860 S.t1746 G.t2860 D.t2370 S.t332 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2861 D.t2369 G.t2861 S.t1745 S.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2862 D.t2368 G.t2862 S.t1744 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2863 S.t1743 G.t2863 D.t2363 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2864 D.t2362 G.t2864 S.t1742 S.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2865 S.t1741 G.t2865 D.t2361 S.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2866 S.t1740 G.t2866 D.t2353 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2867 S.t1739 G.t2867 D.t2352 S.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2868 D.t2351 G.t2868 S.t1738 S.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2869 D.t2350 G.t2869 S.t1737 S.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2870 D.t2349 G.t2870 S.t1736 S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2871 S.t1735 G.t2871 D.t2348 S.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2872 D.t2245 G.t2872 S.t1734 S.t150 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2873 D.t2244 G.t2873 S.t1733 S.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2874 S.t1732 G.t2874 D.t2243 S.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2875 D.t2269 G.t2875 S.t1731 S.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2876 D.t2268 G.t2876 S.t1730 S.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2877 S.t1729 G.t2877 D.t2267 S.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2878 S.t1728 G.t2878 D.t2257 S.t150 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2879 S.t1727 G.t2879 D.t2256 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2880 D.t2255 G.t2880 S.t1726 S.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2881 S.t1725 G.t2881 D.t2252 S.t139 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2882 D.t2251 G.t2882 S.t1724 S.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2883 S.t1723 G.t2883 D.t2250 S.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2884 S.t1722 G.t2884 D.t2235 S.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2885 D.t2234 G.t2885 S.t1721 S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2886 D.t2233 G.t2886 S.t1720 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2887 S.t1719 G.t2887 D.t2215 S.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2888 D.t2214 G.t2888 S.t1718 S.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2889 S.t1717 G.t2889 D.t2213 S.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2890 S.t1716 G.t2890 D.t2025 S.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2891 S.t1715 G.t2891 D.t2024 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2892 S.t1714 G.t2892 D.t2023 S.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2893 D.t1989 G.t2893 S.t1713 S.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2894 S.t1712 G.t2894 D.t1988 S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2895 D.t1987 G.t2895 S.t1711 S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2896 D.t1963 G.t2896 S.t1710 S.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2897 S.t1709 G.t2897 D.t1962 S.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2898 S.t1708 G.t2898 D.t1961 S.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2899 S.t1707 G.t2899 D.t1712 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2900 D.t1711 G.t2900 S.t1706 S.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2901 D.t1710 G.t2901 S.t1705 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2902 S.t1704 G.t2902 D.t984 S.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2903 D.t983 G.t2903 S.t1703 S.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2904 D.t982 G.t2904 S.t1702 S.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2905 D.t1213 G.t2905 S.t1701 S.t538 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2906 S.t1700 G.t2906 D.t1212 S.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2907 S.t1699 G.t2907 D.t1211 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2908 D.t2450 G.t2908 S.t1698 S.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2909 D.t2449 G.t2909 S.t1697 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2910 S.t1696 G.t2910 D.t2448 S.t79 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2911 S.t1695 G.t2911 D.t414 S.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2912 D.t413 G.t2912 S.t1694 S.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2913 D.t412 G.t2913 S.t1693 S.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2914 S.t1692 G.t2914 D.t821 S.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2915 S.t1691 G.t2915 D.t820 S.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2916 S.t1690 G.t2916 D.t819 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2917 S.t1689 G.t2917 D.t987 S.t79 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2918 D.t986 G.t2918 S.t1688 S.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2919 S.t1687 G.t2919 D.t985 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2920 S.t1686 G.t2920 D.t857 S.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2921 D.t856 G.t2921 S.t1685 S.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2922 D.t855 G.t2922 S.t1684 S.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2923 S.t1683 G.t2923 D.t839 S.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2924 S.t1682 G.t2924 D.t838 S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2925 D.t837 G.t2925 S.t1681 S.t150 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2926 S.t1680 G.t2926 D.t529 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2927 S.t1679 G.t2927 D.t528 S.t139 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2928 D.t527 G.t2928 S.t1678 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2929 D.t3227 G.t2929 S.t1677 S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2930 D.t3226 G.t2930 S.t1676 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2931 S.t1675 G.t2931 D.t3225 S.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2932 S.t1674 G.t2932 D.t3758 S.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2933 S.t1673 G.t2933 D.t3757 S.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2934 S.t1672 G.t2934 D.t3756 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2935 D.t3828 G.t2935 S.t1671 S.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2936 D.t3827 G.t2936 S.t1670 S.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2937 S.t1669 G.t2937 D.t3826 S.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2938 S.t1668 G.t2938 D.t3271 S.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2939 S.t1667 G.t2939 D.t3270 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2940 S.t1666 G.t2940 D.t3269 S.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2941 S.t1665 G.t2941 D.t3811 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2942 S.t1664 G.t2942 D.t3810 S.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2943 D.t3809 G.t2943 S.t1663 S.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2944 S.t1662 G.t2944 D.t3274 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2945 S.t1661 G.t2945 D.t3273 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2946 D.t3272 G.t2946 S.t1660 S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2947 D.t326 G.t2947 S.t1659 S.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2948 S.t1658 G.t2948 D.t325 S.t231 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2949 S.t1657 G.t2949 D.t324 S.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2950 D.t187 G.t2950 S.t1656 S.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2951 S.t1655 G.t2951 D.t186 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2952 S.t1654 G.t2952 D.t185 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2953 S.t1653 G.t2953 D.t2587 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2954 S.t1652 G.t2954 D.t2586 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2955 S.t1651 G.t2955 D.t2585 S.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2956 S.t1650 G.t2956 D.t273 S.t218 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2957 S.t1649 G.t2957 D.t272 S.t216 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2958 S.t1648 G.t2958 D.t271 S.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2959 D.t3211 G.t2959 S.t1647 S.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2960 S.t1646 G.t2960 D.t3210 S.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2961 S.t1645 G.t2961 D.t3209 S.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2962 S.t1644 G.t2962 D.t1048 S.t158 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2963 D.t1047 G.t2963 S.t1643 S.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2964 S.t1642 G.t2964 D.t1046 S.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2965 S.t1641 G.t2965 D.t2324 S.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2966 S.t1640 G.t2966 D.t2323 S.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2967 S.t1639 G.t2967 D.t2322 S.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2968 D.t2319 G.t2968 S.t1638 S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2969 S.t1637 G.t2969 D.t2318 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2970 S.t1636 G.t2970 D.t2317 S.t209 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2971 S.t1635 G.t2971 D.t2312 S.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2972 S.t1634 G.t2972 D.t2311 S.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2973 D.t2310 G.t2973 S.t1633 S.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2974 S.t1632 G.t2974 D.t386 S.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2975 D.t385 G.t2975 S.t1631 S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2976 S.t1630 G.t2976 D.t384 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2977 D.t2636 G.t2977 S.t1629 S.t406 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2978 D.t2635 G.t2978 S.t1628 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2979 S.t1627 G.t2979 D.t2607 S.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2980 S.t1626 G.t2980 D.t2606 S.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2981 S.t1625 G.t2981 D.t2605 S.t183 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2982 S.t1624 G.t2982 D.t2604 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2983 D.t627 G.t2983 S.t1623 S.t538 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2984 D.t626 G.t2984 S.t1622 S.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2985 S.t1621 G.t2985 D.t2222 S.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2986 S.t1620 G.t2986 D.t2221 S.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2987 D.t2249 G.t2987 S.t1619 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2988 D.t2248 G.t2988 S.t1618 S.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2989 S.t1617 G.t2989 D.t2093 S.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2990 S.t1616 G.t2990 D.t2092 S.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2991 S.t1615 G.t2991 D.t2446 S.t216 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2992 S.t1614 G.t2992 D.t2445 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2993 D.t2443 G.t2993 S.t1613 S.t183 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2994 S.t1612 G.t2994 D.t2442 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2995 S.t1611 G.t2995 D.t2441 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2996 S.t1610 G.t2996 D.t2440 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2997 S.t1609 G.t2997 D.t2426 S.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2998 D.t2425 G.t2998 S.t1608 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2999 D.t2415 G.t2999 S.t1607 S.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3000 S.t1606 G.t3000 D.t2414 S.t176 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3001 S.t1605 G.t3001 D.t2410 S.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3002 D.t2409 G.t3002 S.t1604 S.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3003 S.t1603 G.t3003 D.t2407 S.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3004 D.t2406 G.t3004 S.t1602 S.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3005 S.t1601 G.t3005 D.t2398 S.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3006 S.t1600 G.t3006 D.t2397 S.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3007 D.t2387 G.t3007 S.t1599 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3008 D.t2386 G.t3008 S.t1598 S.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3009 S.t1597 G.t3009 D.t2382 S.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3010 S.t1596 G.t3010 D.t2381 S.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3011 D.t2380 G.t3011 S.t1595 S.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3012 S.t1594 G.t3012 D.t2379 S.t158 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3013 D.t2377 G.t3013 S.t1593 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3014 S.t1592 G.t3014 D.t2376 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3015 D.t2375 G.t3015 S.t1591 S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3016 D.t2374 G.t3016 S.t1590 S.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3017 S.t1589 G.t3017 D.t2372 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3018 D.t2371 G.t3018 S.t1588 S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3019 S.t1587 G.t3019 D.t2367 S.t150 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3020 S.t1586 G.t3020 D.t2366 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3021 D.t2365 G.t3021 S.t1585 S.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3022 S.t1584 G.t3022 D.t2364 S.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3023 D.t2360 G.t3023 S.t1583 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3024 S.t1582 G.t3024 D.t2359 S.t357 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3025 S.t1581 G.t3025 D.t2357 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3026 S.t1580 G.t3026 D.t2356 S.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3027 D.t2355 G.t3027 S.t1579 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3028 D.t2354 G.t3028 S.t1578 S.t79 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3029 S.t1577 G.t3029 D.t2347 S.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3030 D.t2346 G.t3030 S.t1576 S.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3031 S.t1575 G.t3031 D.t2345 S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3032 S.t1574 G.t3032 D.t2344 S.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3033 S.t1573 G.t3033 D.t1335 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3034 S.t1572 G.t3034 D.t1334 S.t321 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3035 S.t1571 G.t3035 D.t1323 S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3036 D.t1322 G.t3036 S.t1570 S.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3037 S.t1569 G.t3037 D.t2288 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3038 S.t1568 G.t3038 D.t2287 S.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3039 S.t1567 G.t3039 D.t2285 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3040 D.t2284 G.t3040 S.t1566 S.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3041 D.t2281 G.t3041 S.t1565 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3042 S.t1564 G.t3042 D.t2280 S.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3043 S.t1563 G.t3043 D.t2277 S.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3044 S.t1562 G.t3044 D.t2276 S.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3045 D.t2273 G.t3045 S.t1561 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3046 S.t1560 G.t3046 D.t2272 S.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3047 D.t2264 G.t3047 S.t1559 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3048 D.t2263 G.t3048 S.t1558 S.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3049 S.t1557 G.t3049 D.t2261 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3050 D.t2260 G.t3050 S.t1556 S.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3051 S.t1555 G.t3051 D.t2247 S.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3052 S.t1554 G.t3052 D.t2246 S.t79 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3053 D.t2241 G.t3053 S.t1553 S.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3054 D.t2240 G.t3054 S.t1552 S.t139 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3055 S.t1551 G.t3055 D.t2237 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3056 D.t2236 G.t3056 S.t1550 S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3057 D.t2229 G.t3057 S.t1549 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3058 D.t2228 G.t3058 S.t1548 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3059 S.t1547 G.t3059 D.t2225 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3060 S.t1546 G.t3060 D.t2224 S.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3061 S.t1545 G.t3061 D.t2140 S.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3062 S.t1544 G.t3062 D.t2139 S.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3063 D.t2138 G.t3063 S.t1543 S.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3064 S.t1542 G.t3064 D.t2137 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3065 S.t1541 G.t3065 D.t2135 S.t79 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3066 D.t2134 G.t3066 S.t1540 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3067 S.t1539 G.t3067 D.t2132 S.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3068 S.t1538 G.t3068 D.t2131 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3069 S.t1537 G.t3069 D.t2128 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3070 D.t2127 G.t3070 S.t1536 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3071 S.t1535 G.t3071 D.t2126 S.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3072 S.t1534 G.t3072 D.t2125 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3073 S.t1533 G.t3073 D.t2124 S.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3074 S.t1532 G.t3074 D.t2123 S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3075 D.t2121 G.t3075 S.t1531 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3076 D.t2120 G.t3076 S.t1530 S.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3077 S.t1529 G.t3077 D.t2118 S.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3078 S.t1528 G.t3078 D.t2117 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3079 D.t2116 G.t3079 S.t1527 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3080 S.t1526 G.t3080 D.t2115 S.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3081 D.t2113 G.t3081 S.t1525 S.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3082 S.t1524 G.t3082 D.t2112 S.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3083 S.t1523 G.t3083 D.t2110 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3084 S.t1522 G.t3084 D.t2109 S.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3085 D.t2108 G.t3085 S.t1521 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3086 D.t2107 G.t3086 S.t1520 S.t218 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3087 S.t1519 G.t3087 D.t2105 S.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3088 S.t1518 G.t3088 D.t2104 S.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3089 S.t1517 G.t3089 D.t2102 S.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3090 D.t2101 G.t3090 S.t1516 S.t443 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3091 S.t1515 G.t3091 D.t2099 S.t209 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3092 D.t2098 G.t3092 S.t1514 S.t158 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3093 D.t2095 G.t3093 S.t1513 S.t270 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3094 D.t2094 G.t3094 S.t1512 S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3095 D.t2091 G.t3095 S.t1511 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3096 D.t2090 G.t3096 S.t1510 S.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3097 S.t1509 G.t3097 D.t2089 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3098 D.t2088 G.t3098 S.t1508 S.t209 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3099 S.t1507 G.t3099 D.t2078 S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3100 S.t1506 G.t3100 D.t2077 S.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3101 D.t2020 G.t3101 S.t1505 S.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3102 S.t1504 G.t3102 D.t2019 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3103 S.t1503 G.t3103 D.t1978 S.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3104 D.t1977 G.t3104 S.t1502 S.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3105 D.t1974 G.t3105 S.t1501 S.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3106 D.t1973 G.t3106 S.t1500 S.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3107 D.t2030 G.t3107 S.t1499 S.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3108 S.t1498 G.t3108 D.t2029 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3109 S.t1497 G.t3109 D.t2027 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3110 D.t2026 G.t3110 S.t1496 S.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3111 D.t2015 G.t3111 S.t1495 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3112 S.t1494 G.t3112 D.t2014 S.t538 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3113 D.t1968 G.t3113 S.t1493 S.t198 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3114 D.t1967 G.t3114 S.t1492 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3115 S.t1491 G.t3115 D.t1952 S.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3116 S.t1490 G.t3116 D.t1951 S.t218 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3117 D.t1881 G.t3117 S.t1489 S.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3118 D.t1880 G.t3118 S.t1488 S.t79 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3119 S.t1487 G.t3119 D.t1869 S.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3120 D.t1868 G.t3120 S.t1486 S.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3121 D.t1839 G.t3121 S.t1485 S.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3122 S.t1484 G.t3122 D.t1838 S.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3123 S.t1483 G.t3123 D.t1824 S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3124 S.t1482 G.t3124 D.t1823 S.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3125 D.t1816 G.t3125 S.t1481 S.t139 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3126 S.t1480 G.t3126 D.t1815 S.t158 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3127 S.t1479 G.t3127 D.t1799 S.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3128 S.t1478 G.t3128 D.t1798 S.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3129 S.t1477 G.t3129 D.t1586 S.t321 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3130 D.t1585 G.t3130 S.t1476 S.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3131 D.t1619 G.t3131 S.t1475 S.t79 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3132 D.t1618 G.t3132 S.t1474 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3133 S.t1473 G.t3133 D.t1513 S.t209 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3134 S.t1472 G.t3134 D.t1512 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3135 S.t1471 G.t3135 D.t1559 S.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3136 D.t1558 G.t3136 S.t1470 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3137 S.t1469 G.t3137 D.t1506 S.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3138 S.t1468 G.t3138 D.t1505 S.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3139 D.t1339 G.t3139 S.t1467 S.t406 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3140 D.t1338 G.t3140 S.t1466 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3141 D.t1315 G.t3141 S.t1465 S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3142 D.t1314 G.t3142 S.t1464 S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3143 S.t1463 G.t3143 D.t1117 S.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3144 D.t1116 G.t3144 S.t1462 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3145 D.t1114 G.t3145 S.t1461 S.t198 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3146 S.t1460 G.t3146 D.t1113 S.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3147 D.t989 G.t3147 S.t1459 S.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3148 S.t1458 G.t3148 D.t988 S.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3149 S.t1457 G.t3149 D.t1720 S.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3150 D.t1719 G.t3150 S.t1456 S.t332 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3151 S.t1455 G.t3151 D.t235 S.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3152 D.t234 G.t3152 S.t1454 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3153 S.t1453 G.t3153 D.t2574 S.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3154 D.t2573 G.t3154 S.t1452 S.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3155 D.t2578 G.t3155 S.t1451 S.t150 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3156 D.t2577 G.t3156 S.t1450 S.t198 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3157 S.t1449 G.t3157 D.t2580 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3158 S.t1448 G.t3158 D.t2579 S.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3159 D.t2582 G.t3159 S.t1447 S.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3160 S.t1446 G.t3160 D.t2581 S.t176 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3161 D.t40 G.t3161 S.t1445 S.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3162 D.t39 G.t3162 S.t1444 S.t332 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3163 S.t1443 G.t3163 D.t2455 S.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3164 D.t2454 G.t3164 S.t1442 S.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3165 D.t4 G.t3165 S.t1441 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3166 S.t1440 G.t3166 D.t3 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3167 D.t6 G.t3167 S.t1439 S.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3168 D.t5 G.t3168 S.t1438 S.t231 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3169 D.t13 G.t3169 S.t1437 S.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3170 S.t1436 G.t3170 D.t12 S.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3171 D.t1776 G.t3171 S.t1435 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3172 S.t1434 G.t3172 D.t1775 S.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3173 S.t1433 G.t3173 D.t496 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3174 D.t495 G.t3174 S.t1432 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3175 D.t938 G.t3175 S.t1431 S.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3176 S.t1430 G.t3176 D.t937 S.t158 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3177 D.t955 G.t3177 S.t1429 S.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3178 D.t954 G.t3178 S.t1428 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3179 D.t1623 G.t3179 S.t1427 S.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3180 D.t1622 G.t3180 S.t1426 S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3181 D.t1578 G.t3181 S.t1425 S.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3182 S.t1424 G.t3182 D.t1577 S.t388 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3183 S.t1423 G.t3183 D.t1533 S.t150 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3184 D.t1532 G.t3184 S.t1422 S.t218 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3185 D.t1706 G.t3185 S.t1421 S.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3186 S.t1420 G.t3186 D.t1705 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3187 D.t1163 G.t3187 S.t1419 S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3188 D.t1162 G.t3188 S.t1418 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3189 S.t1417 G.t3189 D.t958 S.t209 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3190 S.t1416 G.t3190 D.t957 S.t139 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3191 D.t879 G.t3191 S.t1415 S.t158 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3192 D.t878 G.t3192 S.t1414 S.t332 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3193 S.t1413 G.t3193 D.t655 S.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3194 D.t654 G.t3194 S.t1412 S.t209 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3195 S.t1411 G.t3195 D.t645 S.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3196 S.t1410 G.t3196 D.t644 S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3197 S.t1409 G.t3197 D.t625 S.t357 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3198 D.t624 G.t3198 S.t1408 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3199 S.t1407 G.t3199 D.t616 S.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3200 D.t615 G.t3200 S.t1406 S.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3201 D.t597 G.t3201 S.t1405 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3202 S.t1404 G.t3202 D.t596 S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3203 D.t588 G.t3203 S.t1403 S.t79 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3204 D.t587 G.t3204 S.t1402 S.t198 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3205 D.t567 G.t3205 S.t1401 S.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3206 D.t566 G.t3206 S.t1400 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3207 S.t1399 G.t3207 D.t532 S.t321 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3208 D.t531 G.t3208 S.t1398 S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3209 D.t516 G.t3209 S.t1397 S.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3210 D.t515 G.t3210 S.t1396 S.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3211 D.t503 G.t3211 S.t1395 S.t79 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3212 D.t502 G.t3212 S.t1394 S.t216 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3213 S.t1393 G.t3213 D.t487 S.t218 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3214 D.t486 G.t3214 S.t1392 S.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3215 D.t449 G.t3215 S.t1391 S.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3216 D.t448 G.t3216 S.t1390 S.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3217 S.t1389 G.t3217 D.t145 S.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3218 S.t1388 G.t3218 D.t144 S.t183 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3219 S.t1387 G.t3219 D.t2610 S.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3220 D.t2609 G.t3220 S.t1386 S.t139 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3221 D.t2341 G.t3221 S.t1385 S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3222 D.t2340 G.t3222 S.t1384 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3223 D.t2335 G.t3223 S.t1383 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3224 D.t2334 G.t3224 S.t1382 S.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3225 D.t2314 G.t3225 S.t1381 S.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3226 S.t1380 G.t3226 D.t2313 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3227 S.t1379 G.t3227 D.t2309 S.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3228 S.t1378 G.t3228 D.t2308 S.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3229 D.t345 G.t3229 S.t1377 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3230 D.t344 G.t3230 S.t1376 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3231 D.t331 G.t3231 S.t1375 S.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3232 S.t1374 G.t3232 D.t330 S.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3233 D.t2307 G.t3233 S.t1373 S.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3234 D.t2306 G.t3234 S.t1372 S.t270 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3235 D.t2316 G.t3235 S.t1371 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3236 D.t2315 G.t3236 S.t1370 S.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3237 S.t1369 G.t3237 D.t2321 S.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3238 D.t2320 G.t3238 S.t1368 S.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3239 S.t1367 G.t3239 D.t2338 S.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3240 S.t1366 G.t3240 D.t2337 S.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3241 S.t1365 G.t3241 D.t428 S.t270 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3242 S.t1364 G.t3242 D.t427 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3243 D.t3930 G.t3243 S.t1363 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3244 D.t3929 G.t3244 S.t1362 S.t332 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3245 S.t1361 G.t3245 D.t3702 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3246 D.t3701 G.t3246 S.t1360 S.t388 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3247 S.t1359 G.t3247 D.t3525 S.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3248 D.t3524 G.t3248 S.t1358 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3249 D.t3969 G.t3249 S.t1357 S.t150 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3250 S.t1356 G.t3250 D.t3968 S.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3251 D.t1361 G.t3251 S.t1355 S.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3252 S.t1354 G.t3252 D.t1360 S.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3253 D.t469 G.t3253 S.t1353 S.t198 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3254 D.t468 G.t3254 S.t1352 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3255 D.t460 G.t3255 S.t1351 S.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3256 S.t1350 G.t3256 D.t459 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3257 D.t2018 G.t3257 S.t1349 S.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3258 S.t1348 G.t3258 D.t2017 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3259 D.t1985 G.t3259 S.t1347 S.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3260 D.t1984 G.t3260 S.t1346 S.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3261 D.t1634 G.t3261 S.t1345 S.t218 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3262 D.t1633 G.t3262 S.t1344 S.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3263 S.t1343 G.t3263 D.t1581 S.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3264 S.t1342 G.t3264 D.t1580 S.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3265 D.t1557 G.t3265 S.t1341 S.t443 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3266 S.t1340 G.t3266 D.t1556 S.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3267 D.t1672 G.t3267 S.t1339 S.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3268 D.t1671 G.t3268 S.t1338 S.t158 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3269 D.t1636 G.t3269 S.t1337 S.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3270 D.t1635 G.t3270 S.t1336 S.t270 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3271 D.t1543 G.t3271 S.t1335 S.t321 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3272 D.t1542 G.t3272 S.t1334 S.t209 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3273 S.t1333 G.t3273 D.t1522 S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3274 D.t1521 G.t3274 S.t1332 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3275 S.t1331 G.t3275 D.t1520 S.t388 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3276 D.t1519 G.t3276 S.t1330 S.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3277 S.t1329 G.t3277 D.t1583 S.t216 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3278 D.t1582 G.t3278 S.t1328 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3279 D.t1161 G.t3279 S.t1327 S.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3280 S.t1326 G.t3280 D.t1160 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3281 D.t1159 G.t3281 S.t1325 S.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3282 D.t1158 G.t3282 S.t1324 S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3283 S.t1323 G.t3283 D.t518 S.t406 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3284 S.t1322 G.t3284 D.t517 S.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3285 D.t875 G.t3285 S.t1321 S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3286 D.t874 G.t3286 S.t1320 S.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3287 S.t1319 G.t3287 D.t747 S.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3288 S.t1318 G.t3288 D.t746 S.t538 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3289 D.t734 G.t3289 S.t1317 S.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3290 S.t1316 G.t3290 D.t733 S.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3291 D.t732 G.t3291 S.t1315 S.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3292 D.t731 G.t3292 S.t1314 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3293 D.t610 G.t3293 S.t1313 S.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3294 S.t1312 G.t3294 D.t609 S.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3295 D.t485 G.t3295 S.t1311 S.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3296 D.t484 G.t3296 S.t1310 S.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3297 D.t269 G.t3297 S.t1309 S.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3298 S.t1308 G.t3298 D.t268 S.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3299 S.t1307 G.t3299 D.t674 S.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3300 D.t673 G.t3300 S.t1306 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3301 D.t2652 G.t3301 S.t1305 S.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3302 D.t2651 G.t3302 S.t1304 S.t139 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3303 D.t2598 G.t3303 S.t1303 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3304 S.t1302 G.t3304 D.t2597 S.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3305 S.t1301 G.t3305 D.t2343 S.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3306 D.t2342 G.t3306 S.t1300 S.t176 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3307 S.t1299 G.t3307 D.t2305 S.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3308 D.t2304 G.t3308 S.t1298 S.t79 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3309 D.t2299 G.t3309 S.t1297 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3310 D.t2298 G.t3310 S.t1296 S.t216 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3311 D.t3499 G.t3311 S.t1295 S.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3312 S.t1294 G.t3312 D.t3498 S.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3313 D.t221 G.t3313 S.t1293 S.t406 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3314 D.t220 G.t3314 S.t1292 S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3315 D.t304 G.t3315 S.t1291 S.t198 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3316 S.t1290 G.t3316 D.t303 S.t150 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3317 D.t317 G.t3317 S.t1289 S.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3318 S.t1288 G.t3318 D.t316 S.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3319 D.t311 G.t3319 S.t1287 S.t158 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3320 S.t1286 G.t3320 D.t310 S.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3321 S.t1285 G.t3321 D.t302 S.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3322 D.t301 G.t3322 S.t1284 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3323 D.t3208 G.t3323 S.t1283 S.t332 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3324 S.t1282 G.t3324 D.t3207 S.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3325 D.t3213 G.t3325 S.t1281 S.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3326 D.t3212 G.t3326 S.t1280 S.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3327 D.t296 G.t3327 S.t1279 S.t198 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3328 D.t295 G.t3328 S.t1278 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3329 S.t1277 G.t3329 D.t1268 S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3330 D.t1267 G.t3330 S.t1276 S.t270 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3331 S.t1275 G.t3331 D.t1608 S.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3332 S.t1274 G.t3332 D.t1607 S.t176 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3333 D.t1342 G.t3333 S.t1273 S.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3334 D.t1341 G.t3334 S.t1272 S.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3335 D.t1325 G.t3335 S.t1271 S.t209 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3336 S.t1270 G.t3336 D.t1324 S.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3337 D.t1546 G.t3337 S.t1269 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3338 S.t1268 G.t3338 D.t1545 S.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3339 D.t1059 G.t3339 S.t1267 S.t357 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3340 S.t1266 G.t3340 D.t1058 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3341 D.t1237 G.t3341 S.t1265 S.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3342 S.t1264 G.t3342 D.t1236 S.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3343 D.t1166 G.t3343 S.t1263 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3344 S.t1262 G.t3344 D.t1165 S.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3345 S.t1261 G.t3345 D.t1179 S.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3346 D.t1178 G.t3346 S.t1260 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3347 D.t1245 G.t3347 S.t1259 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3348 S.t1258 G.t3348 D.t1244 S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3349 S.t1257 G.t3349 D.t1274 S.t158 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3350 D.t1273 G.t3350 S.t1256 S.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3351 D.t1252 G.t3351 S.t1255 S.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3352 S.t1254 G.t3352 D.t1251 S.t388 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3353 D.t2758 G.t3353 S.t1253 S.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3354 D.t2757 G.t3354 S.t1252 S.t218 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3355 S.t1251 G.t3355 D.t119 S.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3356 S.t1250 G.t3356 D.t118 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3357 D.t2594 G.t3357 S.t1249 S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3358 D.t2593 G.t3358 S.t1248 S.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3359 D.t861 G.t3359 S.t1247 S.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3360 D.t860 G.t3360 S.t1246 S.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3361 S.t1245 G.t3361 D.t2211 S.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3362 S.t1244 G.t3362 D.t2210 S.t139 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3363 D.t1875 G.t3363 S.t1243 S.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3364 D.t1874 G.t3364 S.t1242 S.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3365 D.t1867 G.t3365 S.t1241 S.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3366 S.t1240 G.t3366 D.t1866 S.t231 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3367 S.t1239 G.t3367 D.t1859 S.t357 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3368 S.t1238 G.t3368 D.t1858 S.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3369 D.t1851 G.t3369 S.t1237 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3370 D.t1850 G.t3370 S.t1236 S.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3371 S.t1235 G.t3371 D.t1844 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3372 D.t1843 G.t3372 S.t1234 S.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3373 S.t1233 G.t3373 D.t1837 S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3374 D.t1836 G.t3374 S.t1232 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3375 S.t1231 G.t3375 D.t1829 S.t406 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3376 D.t1828 G.t3376 S.t1230 S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3377 S.t1229 G.t3377 D.t1822 S.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3378 D.t1821 G.t3378 S.t1228 S.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3379 D.t1814 G.t3379 S.t1227 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3380 S.t1226 G.t3380 D.t1813 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3381 S.t1225 G.t3381 D.t1805 S.t332 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3382 D.t1804 G.t3382 S.t1224 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3383 S.t1223 G.t3383 D.t1680 S.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3384 D.t1679 G.t3384 S.t1222 S.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3385 D.t1077 G.t3385 S.t1221 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3386 S.t1220 G.t3386 D.t1076 S.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3387 S.t1219 G.t3387 D.t1085 S.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3388 D.t1084 G.t3388 S.t1218 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3389 D.t1090 G.t3389 S.t1217 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3390 S.t1216 G.t3390 D.t1089 S.t198 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3391 S.t1215 G.t3391 D.t1294 S.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3392 S.t1214 G.t3392 D.t1293 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3393 D.t1283 G.t3393 S.t1213 S.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3394 D.t1282 G.t3394 S.t1212 S.t321 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3395 D.t1277 G.t3395 S.t1211 S.t176 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3396 S.t1210 G.t3396 D.t1276 S.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3397 S.t1209 G.t3397 D.t1266 S.t332 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3398 D.t1265 G.t3398 S.t1208 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3399 D.t1256 G.t3399 S.t1207 S.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3400 D.t1255 G.t3400 S.t1206 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3401 S.t1205 G.t3401 D.t1200 S.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3402 S.t1204 G.t3402 D.t1199 S.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3403 S.t1203 G.t3403 D.t1194 S.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3404 S.t1202 G.t3404 D.t1193 S.t176 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3405 D.t1183 G.t3405 S.t1201 S.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3406 S.t1200 G.t3406 D.t1182 S.t443 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3407 D.t960 G.t3407 S.t1199 S.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3408 D.t959 G.t3408 S.t1198 S.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3409 D.t881 G.t3409 S.t1197 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3410 D.t880 G.t3410 S.t1196 S.t158 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3411 S.t1195 G.t3411 D.t859 S.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3412 S.t1194 G.t3412 D.t858 S.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3413 D.t841 G.t3413 S.t1193 S.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3414 S.t1192 G.t3414 D.t840 S.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3415 D.t489 G.t3415 S.t1191 S.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3416 D.t488 G.t3416 S.t1190 S.t388 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3417 D.t447 G.t3417 S.t1189 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3418 S.t1188 G.t3418 D.t446 S.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3419 S.t1187 G.t3419 D.t3771 S.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3420 D.t3770 G.t3420 S.t1186 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3421 S.t1185 G.t3421 D.t3661 S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3422 S.t1184 G.t3422 D.t3660 S.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3423 S.t1183 G.t3423 D.t3224 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3424 S.t1182 G.t3424 D.t3223 S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3425 D.t3294 G.t3425 S.t1181 S.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3426 D.t3293 G.t3426 S.t1180 S.t357 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3427 S.t1179 G.t3427 D.t3336 S.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3428 D.t3335 G.t3428 S.t1178 S.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3429 S.t1177 G.t3429 D.t3472 S.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3430 D.t3471 G.t3430 S.t1176 S.t216 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3431 D.t4106 G.t3431 S.t1175 S.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3432 S.t1174 G.t3432 D.t4105 S.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3433 S.t1173 G.t3433 D.t3474 S.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3434 S.t1172 G.t3434 D.t3473 S.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3435 D.t3920 G.t3435 S.t1171 S.t443 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3436 D.t3919 G.t3436 S.t1170 S.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3437 D.t3835 G.t3437 S.t1169 S.t321 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3438 D.t3834 G.t3438 S.t1168 S.t270 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3439 D.t3799 G.t3439 S.t1167 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3440 D.t3798 G.t3440 S.t1166 S.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3441 S.t1165 G.t3441 D.t3861 S.t216 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3442 D.t3860 G.t3442 S.t1164 S.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3443 S.t1163 G.t3443 D.t3979 S.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3444 S.t1162 G.t3444 D.t3978 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3445 D.t3623 G.t3445 S.t1161 S.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3446 D.t3622 G.t3446 S.t1160 S.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3447 S.t1159 G.t3447 D.t3637 S.t406 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3448 D.t3636 G.t3448 S.t1158 S.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3449 D.t3252 G.t3449 S.t1157 S.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3450 D.t3251 G.t3450 S.t1156 S.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3451 D.t3501 G.t3451 S.t1155 S.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3452 S.t1154 G.t3452 D.t3500 S.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3453 S.t1153 G.t3453 D.t3416 S.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3454 D.t3415 G.t3454 S.t1152 S.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3455 D.t3576 G.t3455 S.t1151 S.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3456 S.t1150 G.t3456 D.t3575 S.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3457 S.t1149 G.t3457 D.t3904 S.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3458 S.t1148 G.t3458 D.t3903 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3459 D.t3750 G.t3459 S.t1147 S.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3460 S.t1146 G.t3460 D.t3749 S.t270 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3461 D.t3942 G.t3461 S.t1145 S.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3462 D.t3941 G.t3462 S.t1144 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3463 D.t3940 G.t3463 S.t1143 S.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3464 S.t1142 G.t3464 D.t3939 S.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3465 D.t3958 G.t3465 S.t1141 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3466 S.t1140 G.t3466 D.t3957 S.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3467 S.t1139 G.t3467 D.t437 S.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3468 D.t436 G.t3468 S.t1138 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3469 S.t1137 G.t3469 D.t2576 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3470 D.t2575 G.t3470 S.t1136 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3471 D.t2584 G.t3471 S.t1135 S.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3472 D.t2583 G.t3472 S.t1134 S.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3473 S.t1133 G.t3473 D.t319 S.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3474 D.t318 G.t3474 S.t1132 S.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3475 S.t1131 G.t3475 D.t294 S.t150 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3476 S.t1130 G.t3476 D.t293 S.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3477 S.t1129 G.t3477 D.t93 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3478 S.t1128 G.t3478 D.t92 S.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3479 S.t1127 G.t3479 D.t3195 S.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3480 S.t1126 G.t3480 D.t3194 S.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3481 S.t1125 G.t3481 D.t2044 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3482 D.t2043 G.t3482 S.t1124 S.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3483 S.t1123 G.t3483 D.t115 S.t357 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3484 D.t114 G.t3484 S.t1122 S.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3485 D.t2290 G.t3485 S.t1121 S.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3486 S.t1120 G.t3486 D.t2289 S.t443 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3487 S.t1119 G.t3487 D.t2647 S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3488 S.t1118 G.t3488 D.t2646 S.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3489 S.t1117 G.t3489 D.t2631 S.t270 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3490 D.t2630 G.t3490 S.t1116 S.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3491 D.t603 G.t3491 S.t1115 S.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3492 D.t602 G.t3492 S.t1114 S.t209 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3493 S.t1113 G.t3493 D.t2639 S.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3494 S.t1112 G.t3494 D.t2638 S.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3495 D.t2217 G.t3495 S.t1111 S.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3496 D.t2216 G.t3496 S.t1110 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3497 D.t2271 G.t3497 S.t1109 S.t357 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3498 S.t1108 G.t3498 D.t2270 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3499 S.t1107 G.t3499 D.t2034 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3500 S.t1106 G.t3500 D.t2033 S.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3501 S.t1105 G.t3501 D.t2032 S.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3502 S.t1104 G.t3502 D.t2031 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3503 S.t1103 G.t3503 D.t2022 S.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3504 D.t2021 G.t3504 S.t1102 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3505 S.t1101 G.t3505 D.t2009 S.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3506 S.t1100 G.t3506 D.t2008 S.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3507 S.t1099 G.t3507 D.t2007 S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3508 S.t1098 G.t3508 D.t2006 S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3509 D.t2005 G.t3509 S.t1097 S.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3510 D.t2004 G.t3510 S.t1096 S.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3511 S.t1095 G.t3511 D.t1993 S.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3512 D.t1992 G.t3512 S.t1094 S.t216 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3513 S.t1093 G.t3513 D.t1983 S.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3514 S.t1092 G.t3514 D.t1982 S.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3515 S.t1091 G.t3515 D.t1981 S.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3516 D.t1980 G.t3516 S.t1090 S.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3517 S.t1089 G.t3517 D.t1976 S.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3518 D.t1975 G.t3518 S.t1088 S.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3519 S.t1087 G.t3519 D.t1972 S.t139 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3520 D.t1971 G.t3520 S.t1086 S.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3521 S.t1085 G.t3521 D.t1970 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3522 S.t1084 G.t3522 D.t1969 S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3523 D.t1965 G.t3523 S.t1083 S.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3524 S.t1082 G.t3524 D.t1964 S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3525 D.t1960 G.t3525 S.t1081 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3526 S.t1080 G.t3526 D.t1959 S.t198 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3527 D.t1958 G.t3527 S.t1079 S.t176 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3528 D.t1957 G.t3528 S.t1078 S.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3529 S.t1077 G.t3529 D.t1861 S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3530 D.t1860 G.t3530 S.t1076 S.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3531 S.t1075 G.t3531 D.t1853 S.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3532 D.t1852 G.t3532 S.t1074 S.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3533 S.t1073 G.t3533 D.t1846 S.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3534 S.t1072 G.t3534 D.t1845 S.t332 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3535 S.t1071 G.t3535 D.t1682 S.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3536 D.t1681 G.t3536 S.t1070 S.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3537 S.t1069 G.t3537 D.t1676 S.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3538 S.t1068 G.t3538 D.t1675 S.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3539 S.t1067 G.t3539 D.t1625 S.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3540 D.t1624 G.t3540 S.t1066 S.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3541 D.t1704 G.t3541 S.t1065 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3542 S.t1064 G.t3542 D.t1703 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3543 S.t1063 G.t3543 D.t1156 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3544 S.t1062 G.t3544 D.t1155 S.t198 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3545 D.t1154 G.t3545 S.t1061 S.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3546 S.t1060 G.t3546 D.t1153 S.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3547 S.t1059 G.t3547 D.t1151 S.t332 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3548 S.t1058 G.t3548 D.t1150 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3549 S.t1057 G.t3549 D.t1149 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3550 D.t1148 G.t3550 S.t1056 S.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3551 S.t1055 G.t3551 D.t1144 S.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3552 D.t1143 G.t3552 S.t1054 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3553 S.t1053 G.t3553 D.t1140 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3554 D.t1139 G.t3554 S.t1052 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3555 D.t1137 G.t3555 S.t1051 S.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3556 D.t1136 G.t3556 S.t1050 S.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3557 S.t1049 G.t3557 D.t1135 S.t443 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3558 D.t1134 G.t3558 S.t1048 S.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3559 S.t1047 G.t3559 D.t1133 S.t270 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3560 S.t1046 G.t3560 D.t1132 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3561 S.t1045 G.t3561 D.t1128 S.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3562 D.t1127 G.t3562 S.t1044 S.t388 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3563 D.t1125 G.t3563 S.t1043 S.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3564 D.t1124 G.t3564 S.t1042 S.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3565 S.t1041 G.t3565 D.t494 S.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3566 S.t1040 G.t3566 D.t493 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3567 S.t1039 G.t3567 D.t513 S.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3568 D.t512 G.t3568 S.t1038 S.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3569 S.t1037 G.t3569 D.t523 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3570 S.t1036 G.t3570 D.t522 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3571 D.t541 G.t3571 S.t1035 S.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3572 S.t1034 G.t3572 D.t540 S.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3573 D.t981 G.t3573 S.t1033 S.t216 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3574 S.t1032 G.t3574 D.t980 S.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3575 D.t979 G.t3575 S.t1031 S.t321 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3576 S.t1030 G.t3576 D.t978 S.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3577 S.t1029 G.t3577 D.t853 S.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3578 S.t1028 G.t3578 D.t852 S.t216 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3579 D.t834 G.t3579 S.t1027 S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3580 D.t833 G.t3580 S.t1026 S.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3581 S.t1025 G.t3581 D.t2259 S.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3582 S.t1024 G.t3582 D.t2258 S.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3583 S.t1023 G.t3583 D.t2254 S.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3584 D.t2253 G.t3584 S.t1022 S.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3585 D.t2232 G.t3585 S.t1021 S.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3586 D.t2231 G.t3586 S.t1020 S.t150 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3587 S.t1019 G.t3587 D.t2227 S.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3588 D.t2226 G.t3588 S.t1018 S.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3589 S.t1017 G.t3589 D.t2275 S.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3590 S.t1016 G.t3590 D.t2274 S.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3591 D.t683 G.t3591 S.t1015 S.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3592 D.t682 G.t3592 S.t1014 S.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3593 S.t1013 G.t3593 D.t672 S.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3594 D.t671 G.t3594 S.t1012 S.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3595 S.t1011 G.t3595 D.t652 S.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3596 D.t651 G.t3596 S.t1010 S.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3597 S.t1009 G.t3597 D.t642 S.t270 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3598 S.t1008 G.t3598 D.t641 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3599 D.t622 G.t3599 S.t1007 S.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3600 S.t1006 G.t3600 D.t621 S.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3601 S.t1005 G.t3601 D.t612 S.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3602 D.t611 G.t3602 S.t1004 S.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3603 S.t1003 G.t3603 D.t585 S.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3604 D.t584 G.t3604 S.t1002 S.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3605 S.t1001 G.t3605 D.t564 S.t231 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3606 S.t1000 G.t3606 D.t563 S.t150 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3607 S.t999 G.t3607 D.t539 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3608 D.t538 G.t3608 S.t998 S.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3609 S.t997 G.t3609 D.t521 S.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3610 S.t996 G.t3610 D.t520 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3611 S.t995 G.t3611 D.t511 S.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3612 S.t994 G.t3612 D.t510 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3613 D.t2283 G.t3613 S.t993 S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3614 S.t992 G.t3614 D.t2282 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3615 S.t991 G.t3615 D.t492 S.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3616 S.t990 G.t3616 D.t491 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3617 S.t989 G.t3617 D.t2279 S.t357 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3618 S.t988 G.t3618 D.t2278 S.t216 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3619 S.t987 G.t3619 D.t444 S.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3620 D.t443 G.t3620 S.t986 S.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3621 S.t985 G.t3621 D.t108 S.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3622 S.t984 G.t3622 D.t107 S.t270 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3623 S.t983 G.t3623 D.t339 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3624 D.t338 G.t3624 S.t982 S.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3625 S.t981 G.t3625 D.t477 S.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3626 S.t980 G.t3626 D.t476 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3627 S.t979 G.t3627 D.t1678 S.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3628 S.t978 G.t3628 D.t1677 S.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3629 D.t1639 G.t3629 S.t977 S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3630 S.t976 G.t3630 D.t1638 S.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3631 S.t975 G.t3631 D.t1949 S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3632 S.t974 G.t3632 D.t1948 S.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3633 S.t973 G.t3633 D.t1945 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3634 D.t1944 G.t3634 S.t972 S.t538 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3635 S.t971 G.t3635 D.t1943 S.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3636 D.t1942 G.t3636 S.t970 S.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3637 D.t1936 G.t3637 S.t969 S.t443 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3638 S.t968 G.t3638 D.t1935 S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3639 D.t1912 G.t3639 S.t967 S.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3640 S.t966 G.t3640 D.t1911 S.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3641 S.t965 G.t3641 D.t1657 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3642 D.t1656 G.t3642 S.t964 S.t183 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3643 D.t1515 G.t3643 S.t963 S.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3644 S.t962 G.t3644 D.t1514 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3645 D.t1064 G.t3645 S.t961 S.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3646 D.t1063 G.t3646 S.t960 S.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3647 D.t1072 G.t3647 S.t959 S.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3648 D.t1071 G.t3648 S.t958 S.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3649 S.t957 G.t3649 D.t1104 S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3650 D.t1103 G.t3650 S.t956 S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3651 S.t955 G.t3651 D.t1239 S.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3652 D.t1238 G.t3652 S.t954 S.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3653 D.t1109 G.t3653 S.t953 S.t150 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3654 S.t952 G.t3654 D.t1108 S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3655 D.t1292 G.t3655 S.t951 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3656 D.t1291 G.t3656 S.t950 S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3657 S.t949 G.t3657 D.t1281 S.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3658 D.t1280 G.t3658 S.t948 S.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3659 S.t947 G.t3659 D.t1264 S.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3660 S.t946 G.t3660 D.t1263 S.t332 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3661 S.t945 G.t3661 D.t1254 S.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3662 D.t1253 G.t3662 S.t944 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3663 S.t943 G.t3663 D.t1192 S.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3664 D.t1191 G.t3664 S.t942 S.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3665 S.t941 G.t3665 D.t1181 S.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3666 S.t940 G.t3666 D.t1180 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3667 S.t939 G.t3667 D.t1169 S.t198 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3668 D.t1168 G.t3668 S.t938 S.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3669 D.t1099 G.t3669 S.t937 S.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3670 D.t1098 G.t3670 S.t936 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3671 D.t836 G.t3671 S.t935 S.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3672 S.t934 G.t3672 D.t835 S.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3673 S.t933 G.t3673 D.t877 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3674 S.t932 G.t3674 D.t876 S.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3675 S.t931 G.t3675 D.t1231 S.t231 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3676 D.t1230 G.t3676 S.t930 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3677 D.t1202 G.t3677 S.t929 S.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3678 S.t928 G.t3678 D.t1201 S.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3679 D.t1196 G.t3679 S.t927 S.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3680 D.t1195 G.t3680 S.t926 S.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3681 S.t925 G.t3681 D.t1172 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3682 S.t924 G.t3682 D.t1171 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3683 S.t923 G.t3683 D.t1209 S.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3684 D.t1208 G.t3684 S.t922 S.t406 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3685 D.t1215 G.t3685 S.t921 S.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3686 S.t920 G.t3686 D.t1214 S.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3687 D.t1285 G.t3687 S.t919 S.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3688 D.t1284 G.t3688 S.t918 S.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3689 S.t917 G.t3689 D.t467 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3690 D.t466 G.t3690 S.t916 S.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3691 S.t915 G.t3691 D.t439 S.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3692 D.t438 G.t3692 S.t914 S.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3693 S.t913 G.t3693 D.t397 S.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3694 S.t912 G.t3694 D.t396 S.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3695 S.t911 G.t3695 D.t4060 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3696 S.t910 G.t3696 D.t4059 S.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3697 S.t909 G.t3697 D.t3795 S.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3698 S.t908 G.t3698 D.t3794 S.t158 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3699 S.t907 G.t3699 D.t3633 S.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3700 D.t3632 G.t3700 S.t906 S.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3701 S.t905 G.t3701 D.t3574 S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3702 S.t904 G.t3702 D.t3573 S.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3703 S.t903 G.t3703 D.t244 S.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3704 D.t243 G.t3704 S.t902 S.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3705 D.t167 G.t3705 S.t901 S.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3706 D.t166 G.t3706 S.t900 S.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3707 D.t180 G.t3707 S.t899 S.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3708 S.t898 G.t3708 D.t179 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3709 D.t248 G.t3709 S.t897 S.t183 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3710 D.t247 G.t3710 S.t896 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3711 D.t192 G.t3711 S.t895 S.t150 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3712 D.t191 G.t3712 S.t894 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3713 D.t38 G.t3713 S.t893 S.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3714 D.t37 G.t3714 S.t892 S.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3715 S.t891 G.t3715 D.t128 S.t321 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3716 D.t127 G.t3716 S.t890 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3717 S.t889 G.t3717 D.t139 S.t79 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3718 S.t888 G.t3718 D.t138 S.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3719 S.t887 G.t3719 D.t111 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3720 D.t110 G.t3720 S.t886 S.t538 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3721 S.t885 G.t3721 D.t121 S.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3722 D.t120 G.t3722 S.t884 S.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3723 S.t883 G.t3723 D.t102 S.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3724 S.t882 G.t3724 D.t101 S.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3725 D.t106 G.t3725 S.t881 S.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3726 D.t105 G.t3726 S.t880 S.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3727 S.t879 G.t3727 D.t99 S.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3728 S.t878 G.t3728 D.t98 S.t231 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3729 D.t82 G.t3729 S.t877 S.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3730 S.t876 G.t3730 D.t81 S.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3731 D.t88 G.t3731 S.t875 S.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3732 D.t87 G.t3732 S.t874 S.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3733 D.t75 G.t3733 S.t873 S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3734 D.t74 G.t3734 S.t872 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3735 S.t871 G.t3735 D.t78 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3736 S.t870 G.t3736 D.t77 S.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3737 S.t869 G.t3737 D.t69 S.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3738 S.t868 G.t3738 D.t68 S.t357 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3739 S.t867 G.t3739 D.t71 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3740 S.t866 G.t3740 D.t70 S.t216 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3741 D.t66 G.t3741 S.t865 S.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3742 D.t65 G.t3742 S.t864 S.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3743 S.t863 G.t3743 D.t8 S.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3744 S.t862 G.t3744 D.t7 S.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3745 D.t11 G.t3745 S.t861 S.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3746 S.t860 G.t3746 D.t10 S.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3747 D.t15 G.t3747 S.t859 S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3748 S.t858 G.t3748 D.t14 S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3749 D.t17 G.t3749 S.t857 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3750 S.t856 G.t3750 D.t16 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3751 S.t855 G.t3751 D.t20 S.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3752 S.t854 G.t3752 D.t19 S.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3753 D.t1796 G.t3753 S.t853 S.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3754 S.t852 G.t3754 D.t1795 S.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3755 D.t1793 G.t3755 S.t851 S.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3756 S.t850 G.t3756 D.t1792 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3757 D.t1790 G.t3757 S.t849 S.t538 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3758 S.t848 G.t3758 D.t1789 S.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3759 D.t1787 G.t3759 S.t847 S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3760 D.t1786 G.t3760 S.t846 S.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3761 D.t1784 G.t3761 S.t845 S.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3762 D.t1783 G.t3762 S.t844 S.t443 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3763 D.t1781 G.t3763 S.t843 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3764 S.t842 G.t3764 D.t1780 S.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3765 S.t841 G.t3765 D.t1778 S.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3766 S.t840 G.t3766 D.t1777 S.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3767 S.t839 G.t3767 D.t3215 S.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3768 D.t3214 G.t3768 S.t838 S.t183 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3769 S.t837 G.t3769 D.t1740 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3770 S.t836 G.t3770 D.t1739 S.t158 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3771 D.t2146 G.t3771 S.t835 S.t139 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3772 S.t834 G.t3772 D.t2145 S.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3773 D.t1744 G.t3773 S.t833 S.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3774 S.t832 G.t3774 D.t1743 S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3775 S.t831 G.t3775 D.t1747 S.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3776 D.t1746 G.t3776 S.t830 S.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3777 S.t829 G.t3777 D.t1750 S.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3778 D.t1749 G.t3778 S.t828 S.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3779 D.t1753 G.t3779 S.t827 S.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3780 D.t1752 G.t3780 S.t826 S.t231 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3781 D.t1756 G.t3781 S.t825 S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3782 D.t1755 G.t3782 S.t824 S.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3783 S.t823 G.t3783 D.t1759 S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3784 D.t1758 G.t3784 S.t822 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3785 D.t1762 G.t3785 S.t821 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3786 D.t1761 G.t3786 S.t820 S.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3787 S.t819 G.t3787 D.t1765 S.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3788 D.t1764 G.t3788 S.t818 S.t357 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3789 D.t1768 G.t3789 S.t817 S.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3790 D.t1767 G.t3790 S.t816 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3791 D.t1770 G.t3791 S.t815 S.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3792 D.t1769 G.t3792 S.t814 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3793 S.t813 G.t3793 D.t1003 S.t209 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3794 S.t812 G.t3794 D.t1002 S.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3795 S.t811 G.t3795 D.t1005 S.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3796 D.t1004 G.t3796 S.t810 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3797 D.t1007 G.t3797 S.t809 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3798 D.t1006 G.t3798 S.t808 S.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3799 D.t1009 G.t3799 S.t807 S.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3800 D.t1008 G.t3800 S.t806 S.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3801 D.t1011 G.t3801 S.t805 S.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3802 S.t804 G.t3802 D.t1010 S.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3803 D.t1013 G.t3803 S.t803 S.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3804 D.t1012 G.t3804 S.t802 S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3805 S.t801 G.t3805 D.t1015 S.t218 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3806 S.t800 G.t3806 D.t1014 S.t388 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3807 D.t1017 G.t3807 S.t799 S.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3808 S.t798 G.t3808 D.t1016 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3809 D.t1019 G.t3809 S.t797 S.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3810 S.t796 G.t3810 D.t1018 S.t183 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3811 S.t795 G.t3811 D.t1021 S.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3812 D.t1020 G.t3812 S.t794 S.t406 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3813 S.t793 G.t3813 D.t1023 S.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3814 D.t1022 G.t3814 S.t792 S.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3815 S.t791 G.t3815 D.t1025 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3816 D.t1024 G.t3816 S.t790 S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3817 D.t1027 G.t3817 S.t789 S.t183 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3818 S.t788 G.t3818 D.t1026 S.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3819 S.t787 G.t3819 D.t1029 S.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3820 D.t1028 G.t3820 S.t786 S.t79 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3821 S.t785 G.t3821 D.t1031 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3822 S.t784 G.t3822 D.t1030 S.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3823 S.t783 G.t3823 D.t1033 S.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3824 S.t782 G.t3824 D.t1032 S.t218 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3825 D.t1035 G.t3825 S.t781 S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3826 D.t1034 G.t3826 S.t780 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3827 S.t779 G.t3827 D.t1037 S.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3828 S.t778 G.t3828 D.t1036 S.t321 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3829 D.t2615 G.t3829 S.t777 S.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3830 S.t776 G.t3830 D.t1340 S.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3831 S.t775 G.t3831 D.t1316 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3832 D.t2300 G.t3832 S.t774 S.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3833 D.t2302 G.t3833 S.t773 S.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3834 S.t772 G.t3834 D.t475 S.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3835 D.t328 G.t3835 S.t771 S.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3836 D.t327 G.t3836 S.t770 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3837 S.t769 G.t3837 D.t112 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3838 D.t150 G.t3838 S.t768 S.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3839 D.t2696 G.t3839 S.t767 S.t406 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3840 D.t2752 G.t3840 S.t766 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3841 D.t2672 G.t3841 S.t765 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3842 S.t764 G.t3842 D.t2634 S.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3843 S.t763 G.t3843 D.t2645 S.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3844 D.t2608 G.t3844 S.t762 S.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3845 S.t761 G.t3845 D.t2038 S.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3846 S.t760 G.t3846 D.t2012 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3847 D.t2010 G.t3847 S.t759 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3848 D.t1986 G.t3848 S.t758 S.t357 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3849 S.t757 G.t3849 D.t1947 S.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3850 D.t1946 G.t3850 S.t756 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3851 D.t1938 G.t3851 S.t755 S.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3852 D.t1937 G.t3852 S.t754 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3853 S.t753 G.t3853 D.t1934 S.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3854 S.t752 G.t3854 D.t1933 S.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3855 S.t751 G.t3855 D.t1932 S.t388 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3856 D.t1910 G.t3856 S.t750 S.t538 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3857 S.t749 G.t3857 D.t1891 S.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3858 S.t748 G.t3858 D.t1609 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3859 S.t747 G.t3859 D.t1621 S.t321 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3860 S.t746 G.t3860 D.t1606 S.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3861 S.t745 G.t3861 D.t1576 S.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3862 S.t744 G.t3862 D.t1561 S.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3863 D.t1534 G.t3863 S.t743 S.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3864 S.t742 G.t3864 D.t1530 S.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3865 D.t1707 G.t3865 S.t741 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3866 S.t740 G.t3866 D.t1718 S.t231 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3867 D.t1504 G.t3867 S.t739 S.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3868 D.t1569 G.t3868 S.t738 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3869 D.t1555 G.t3869 S.t737 S.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3870 S.t736 G.t3870 D.t1517 S.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3871 D.t1516 G.t3871 S.t735 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3872 D.t2238 G.t3872 S.t734 S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3873 S.t733 G.t3873 D.t1173 S.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3874 S.t732 G.t3874 D.t1167 S.t538 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3875 D.t1617 G.t3875 S.t731 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3876 D.t1186 G.t3876 S.t730 S.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3877 S.t729 G.t3877 D.t1210 S.t218 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3878 D.t1222 G.t3878 S.t728 S.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3879 S.t727 G.t3879 D.t1232 S.t216 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3880 S.t726 G.t3880 D.t1226 S.t357 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3881 D.t1319 G.t3881 S.t725 S.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3882 D.t1246 G.t3882 S.t724 S.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3883 D.t1950 G.t3883 S.t723 S.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3884 D.t1257 G.t3884 S.t722 S.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3885 S.t721 G.t3885 D.t1669 S.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3886 S.t720 G.t3886 D.t1575 S.t176 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3887 D.t1507 G.t3887 S.t719 S.t158 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3888 S.t718 G.t3888 D.t1509 S.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3889 D.t1197 G.t3889 S.t717 S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3890 S.t716 G.t3890 D.t1510 S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3891 S.t715 G.t3891 D.t1511 S.t357 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3892 D.t1279 G.t3892 S.t714 S.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3893 D.t1286 G.t3893 S.t713 S.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3894 S.t712 G.t3894 D.t1146 S.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3895 D.t1142 G.t3895 S.t711 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3896 S.t710 G.t3896 D.t1131 S.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3897 D.t595 G.t3897 S.t709 S.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3898 S.t708 G.t3898 D.t613 S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3899 D.t643 G.t3899 S.t707 S.t198 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3900 D.t900 G.t3900 S.t706 S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3901 D.t1348 G.t3901 S.t705 S.t538 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3902 S.t704 G.t3902 D.t976 S.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3903 D.t681 G.t3903 S.t703 S.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3904 S.t702 G.t3904 D.t573 S.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3905 D.t519 G.t3905 S.t701 S.t443 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3906 S.t700 G.t3906 D.t1321 S.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3907 D.t500 G.t3907 S.t699 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3908 D.t1296 G.t3908 S.t698 S.t388 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3909 S.t697 G.t3909 D.t1278 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3910 D.t995 G.t3910 S.t696 S.t139 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3911 D.t482 G.t3911 S.t695 S.t270 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3912 S.t694 G.t3912 D.t483 S.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3913 D.t371 G.t3913 S.t693 S.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3914 S.t692 G.t3914 D.t253 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3915 S.t691 G.t3915 D.t261 S.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3916 D.t3723 G.t3916 S.t690 S.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3917 D.t3287 G.t3917 S.t689 S.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3918 D.t4132 G.t3918 S.t688 S.t332 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3919 D.t4133 G.t3919 S.t687 S.t231 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3920 D.t3917 G.t3920 S.t686 S.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3921 D.t4136 G.t3921 S.t685 S.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3922 D.t3295 G.t3922 S.t684 S.t406 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3923 D.t3538 G.t3923 S.t683 S.t231 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3924 S.t682 G.t3924 D.t4109 S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3925 S.t681 G.t3925 D.t3662 S.t321 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3926 S.t680 G.t3926 D.t259 S.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3927 D.t4079 G.t3927 S.t679 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3928 S.t678 G.t3928 D.t3520 S.t183 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3929 S.t677 G.t3929 D.t3868 S.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3930 D.t3699 G.t3930 S.t676 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3931 S.t675 G.t3931 D.t3911 S.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3932 D.t3261 G.t3932 S.t674 S.t357 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3933 D.t3625 G.t3933 S.t673 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3934 D.t4082 G.t3934 S.t672 S.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3935 S.t671 G.t3935 D.t3442 S.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3936 S.t670 G.t3936 D.t3793 S.t388 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3937 S.t669 G.t3937 D.t3631 S.t406 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3938 S.t668 G.t3938 D.t3262 S.t209 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3939 D.t3620 G.t3939 S.t667 S.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3940 S.t666 G.t3940 D.t4063 S.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3941 D.t4156 G.t3941 S.t665 S.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3942 D.t4126 G.t3942 S.t664 S.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3943 S.t663 G.t3943 D.t4073 S.t231 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3944 D.t3621 G.t3944 S.t662 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3945 S.t661 G.t3945 D.t3639 S.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3946 D.t3878 G.t3946 S.t660 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3947 S.t659 G.t3947 D.t3487 S.t538 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3948 D.t3971 G.t3948 S.t658 S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3949 S.t657 G.t3949 D.t3522 S.t218 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3950 S.t656 G.t3950 D.t3726 S.t443 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3951 D.t3691 G.t3951 S.t655 S.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3952 S.t654 G.t3952 D.t3263 S.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3953 D.t3517 G.t3953 S.t653 S.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3954 S.t652 G.t3954 D.t411 S.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3955 D.t163 G.t3955 S.t651 S.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3956 S.t650 G.t3956 D.t254 S.t388 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3957 D.t142 G.t3957 S.t649 S.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3958 D.t1050 G.t3958 S.t648 S.t406 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3959 S.t647 G.t3959 D.t1054 S.t183 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3960 S.t646 G.t3960 D.t1055 S.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3961 D.t196 G.t3961 S.t645 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3962 S.t644 G.t3962 D.t1053 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3963 S.t643 G.t3963 D.t1051 S.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3964 S.t642 G.t3964 D.t1052 S.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3965 S.t641 G.t3965 D.t210 S.t332 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3966 S.t640 G.t3966 D.t266 S.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3967 D.t33 G.t3967 S.t639 S.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3968 S.t638 G.t3968 D.t2456 S.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3969 S.t637 G.t3969 D.t3203 S.t357 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3970 S.t636 G.t3970 D.t3200 S.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3971 S.t635 G.t3971 D.t3196 S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3972 D.t3177 G.t3972 S.t634 S.t198 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3973 S.t633 G.t3973 D.t3188 S.t176 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3974 S.t632 G.t3974 D.t3198 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3975 S.t631 G.t3975 D.t1794 S.t538 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3976 D.t1791 G.t3976 S.t630 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3977 D.t1788 G.t3977 S.t629 S.t321 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3978 S.t628 G.t3978 D.t1785 S.t321 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3979 S.t627 G.t3979 D.t1782 S.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3980 S.t626 G.t3980 D.t1779 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3981 S.t625 G.t3981 D.t3197 S.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3982 D.t2209 G.t3982 S.t624 S.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3983 S.t623 G.t3983 D.t399 S.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3984 S.t622 G.t3984 D.t95 S.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3985 S.t621 G.t3985 D.t2722 S.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3986 S.t620 G.t3986 D.t2703 S.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3987 D.t2687 G.t3987 S.t619 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3988 S.t618 G.t3988 D.t450 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3989 S.t617 G.t3989 D.t1797 S.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3990 S.t616 G.t3990 D.t1646 S.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3991 S.t615 G.t3991 D.t586 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3992 D.t465 G.t3992 S.t614 S.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3993 S.t613 G.t3993 D.t1297 S.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3994 S.t612 G.t3994 D.t346 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3995 D.t329 G.t3995 S.t611 S.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3996 S.t610 G.t3996 D.t135 S.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3997 D.t2755 G.t3997 S.t609 S.t332 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3998 S.t608 G.t3998 D.t2764 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3999 D.t2689 G.t3999 S.t607 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4000 S.t606 G.t4000 D.t2763 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4001 S.t605 G.t4001 D.t2663 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4002 D.t2658 G.t4002 S.t604 S.t538 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4003 S.t603 G.t4003 D.t977 S.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4004 D.t1356 G.t4004 S.t602 S.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4005 D.t2301 G.t4005 S.t601 S.t538 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4006 S.t600 G.t4006 D.t2086 S.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4007 S.t599 G.t4007 D.t2085 S.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4008 S.t598 G.t4008 D.t2084 S.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4009 D.t2083 G.t4009 S.t597 S.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4010 S.t596 G.t4010 D.t1953 S.t321 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4011 S.t595 G.t4011 D.t2039 S.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4012 D.t2028 G.t4012 S.t594 S.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4013 D.t2016 G.t4013 S.t593 S.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4014 D.t1990 G.t4014 S.t592 S.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4015 S.t591 G.t4015 D.t1955 S.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4016 S.t590 G.t4016 D.t1118 S.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4017 D.t975 G.t4017 S.t589 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4018 S.t588 G.t4018 D.t1318 S.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4019 S.t587 G.t4019 D.t1336 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4020 D.t1306 G.t4020 S.t586 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4021 D.t1299 G.t4021 S.t585 S.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4022 S.t584 G.t4022 D.t1311 S.t406 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4023 S.t583 G.t4023 D.t2702 S.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4024 D.t369 G.t4024 S.t582 S.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4025 S.t581 G.t4025 D.t267 S.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4026 D.t188 G.t4026 S.t580 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4027 S.t579 G.t4027 D.t246 S.t538 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4028 D.t236 G.t4028 S.t578 S.t139 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4029 D.t255 G.t4029 S.t577 S.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4030 S.t576 G.t4030 D.t2566 S.t443 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4031 D.t270 G.t4031 S.t575 S.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4032 D.t190 G.t4032 S.t574 S.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4033 D.t129 G.t4033 S.t573 S.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4034 S.t572 G.t4034 D.t178 S.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4035 D.t189 G.t4035 S.t571 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4036 D.t195 G.t4036 S.t570 S.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4037 D.t313 G.t4037 S.t569 S.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4038 D.t308 G.t4038 S.t568 S.t443 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4039 D.t321 G.t4039 S.t567 S.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4040 S.t566 G.t4040 D.t320 S.t139 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4041 D.t322 G.t4041 S.t565 S.t158 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4042 D.t315 G.t4042 S.t564 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4043 D.t314 G.t4043 S.t563 S.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4044 S.t562 G.t4044 D.t307 S.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4045 D.t306 G.t4045 S.t561 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4046 S.t560 G.t4046 D.t31 S.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4047 S.t559 G.t4047 D.t337 S.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4048 D.t299 G.t4048 S.t558 S.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4049 S.t557 G.t4049 D.t286 S.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4050 D.t298 G.t4050 S.t556 S.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4051 D.t292 G.t4051 S.t555 S.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4052 S.t554 G.t4052 D.t32 S.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4053 S.t553 G.t4053 D.t2291 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4054 D.t25 G.t4054 S.t552 S.t198 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4055 S.t551 G.t4055 D.t300 S.t176 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4056 S.t550 G.t4056 D.t27 S.t406 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4057 S.t549 G.t4057 D.t1742 S.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4058 D.t1745 G.t4058 S.t548 S.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4059 D.t1748 G.t4059 S.t547 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4060 D.t1751 G.t4060 S.t546 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4061 S.t545 G.t4061 D.t1754 S.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4062 D.t1757 G.t4062 S.t544 S.t183 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4063 D.t1760 G.t4063 S.t543 S.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4064 S.t542 G.t4064 D.t1763 S.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4065 D.t1766 G.t4065 S.t541 S.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4066 D.t1057 G.t4066 S.t540 S.t388 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4067 S.t539 G.t4067 D.t1056 S.t538 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4068 D.t1000 G.t4068 S.t537 S.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4069 D.t153 G.t4069 S.t536 S.t270 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4070 D.t2096 G.t4070 S.t535 S.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4071 D.t2671 G.t4071 S.t534 S.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4072 D.t2738 G.t4072 S.t533 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4073 D.t2685 G.t4073 S.t532 S.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4074 D.t2668 G.t4074 S.t531 S.t209 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4075 D.t2648 G.t4075 S.t530 S.t332 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4076 S.t529 G.t4076 D.t2665 S.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4077 S.t528 G.t4077 D.t2644 S.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4078 D.t2653 G.t4078 S.t527 S.t231 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4079 S.t526 G.t4079 D.t2656 S.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4080 D.t2650 G.t4080 S.t525 S.t231 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4081 S.t524 G.t4081 D.t2642 S.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4082 D.t2641 G.t4082 S.t523 S.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4083 D.t2640 G.t4083 S.t522 S.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4084 S.t521 G.t4084 D.t2666 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4085 S.t520 G.t4085 D.t2621 S.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4086 S.t519 G.t4086 D.t2627 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4087 S.t518 G.t4087 D.t2614 S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4088 S.t517 G.t4088 D.t2612 S.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4089 S.t516 G.t4089 D.t2601 S.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4090 D.t2600 G.t4090 S.t515 S.t218 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4091 D.t2595 G.t4091 S.t514 S.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4092 D.t2133 G.t4092 S.t513 S.t388 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4093 D.t2262 G.t4093 S.t512 S.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4094 S.t511 G.t4094 D.t2286 S.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4095 S.t510 G.t4095 D.t2106 S.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4096 S.t509 G.t4096 D.t2111 S.t406 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4097 D.t2119 G.t4097 S.t508 S.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4098 S.t507 G.t4098 D.t2103 S.t209 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4099 D.t2129 G.t4099 S.t506 S.t139 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4100 S.t505 G.t4100 D.t2136 S.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4101 S.t504 G.t4101 D.t2076 S.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4102 D.t2075 G.t4102 S.t503 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4103 D.t2074 G.t4103 S.t502 S.t357 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4104 S.t501 G.t4104 D.t2073 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4105 S.t500 G.t4105 D.t2072 S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4106 S.t499 G.t4106 D.t2071 S.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4107 S.t498 G.t4107 D.t1563 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4108 S.t497 G.t4108 D.t1502 S.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4109 S.t496 G.t4109 D.t1485 S.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4110 D.t1469 G.t4110 S.t495 S.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4111 D.t1453 G.t4111 S.t494 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4112 S.t493 G.t4112 D.t1437 S.t198 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4113 D.t1421 G.t4113 S.t492 S.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4114 S.t491 G.t4114 D.t1405 S.t443 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4115 S.t490 G.t4115 D.t1355 S.t183 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4116 D.t1931 G.t4116 S.t489 S.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4117 S.t488 G.t4117 D.t1882 S.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4118 D.t1275 G.t4118 S.t487 S.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4119 D.t1223 G.t4119 S.t486 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4120 S.t485 G.t4120 D.t1198 S.t183 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4121 S.t484 G.t4121 D.t1170 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4122 D.t1224 G.t4122 S.t483 S.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4123 S.t482 G.t4123 D.t956 S.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4124 S.t481 G.t4124 D.t474 S.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4125 D.t445 G.t4125 S.t480 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4126 S.t479 G.t4126 D.t375 S.t139 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4127 S.t478 G.t4127 D.t2122 S.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4128 D.t2620 G.t4128 S.t477 S.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4129 S.t476 G.t4129 D.t2649 S.t332 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4130 D.t2736 G.t4130 S.t475 S.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4131 S.t474 G.t4131 D.t365 S.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4132 D.t347 G.t4132 S.t473 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4133 D.t3088 G.t4133 S.t472 S.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4134 S.t471 G.t4134 D.t2985 S.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4135 S.t470 G.t4135 D.t176 S.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4136 S.t469 G.t4136 D.t194 S.t176 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4137 D.t174 G.t4137 S.t468 S.t321 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4138 D.t3217 G.t4138 S.t467 S.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4139 S.t466 G.t4139 D.t3218 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4140 D.t113 G.t4140 S.t465 S.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4141 D.t2726 G.t4141 S.t464 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4142 S.t463 G.t4142 D.t131 S.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4143 D.t158 G.t4143 S.t462 S.t183 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4144 S.t461 G.t4144 D.t94 S.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4145 D.t2725 G.t4145 S.t460 S.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4146 D.t2759 G.t4146 S.t459 S.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4147 D.t2940 G.t4147 S.t458 S.t209 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4148 S.t457 G.t4148 D.t2820 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4149 S.t456 G.t4149 D.t2699 S.t139 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4150 D.t2704 G.t4150 S.t455 S.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4151 S.t454 G.t4151 D.t2730 S.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4152 S.t453 G.t4152 D.t2720 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4153 D.t2710 G.t4153 S.t452 S.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4154 S.t451 G.t4154 D.t2748 S.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4155 D.t2701 G.t4155 S.t450 S.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4156 S.t449 G.t4156 D.t2700 S.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4157 S.t448 G.t4157 D.t2694 S.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4158 D.t2688 G.t4158 S.t447 S.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4159 D.t2690 G.t4159 S.t446 S.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4160 D.t2708 G.t4160 S.t445 S.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4161 S.t444 G.t4161 D.t2669 S.t443 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4162 D.t2721 G.t4162 S.t442 S.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4163 D.t2633 G.t4163 S.t441 S.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4164 D.t2622 G.t4164 S.t440 S.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4165 D.t2011 G.t4165 S.t439 S.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4166 D.t1994 G.t4166 S.t438 S.t218 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4167 S.t437 G.t4167 D.t1991 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4168 S.t436 G.t4168 D.t1887 S.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4169 D.t1610 G.t4169 S.t435 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4170 D.t1600 G.t4170 S.t434 S.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4171 D.t1579 G.t4171 S.t433 S.t388 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4172 S.t432 G.t4172 D.t1535 S.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4173 S.t431 G.t4173 D.t1503 S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4174 S.t430 G.t4174 D.t1518 S.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4175 D.t1529 G.t4175 S.t429 S.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4176 D.t1709 G.t4176 S.t428 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4177 D.t1523 G.t4177 S.t427 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4178 D.t565 G.t4178 S.t426 S.t139 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4179 S.t425 G.t4179 D.t1590 S.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4180 D.t1531 G.t4180 S.t424 S.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4181 D.t1152 G.t4181 S.t423 S.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4182 D.t1147 G.t4182 S.t422 S.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4183 D.t1145 G.t4183 S.t421 S.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4184 D.t1141 G.t4184 S.t420 S.t216 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4185 D.t1138 G.t4185 S.t419 S.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4186 D.t1129 G.t4186 S.t418 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4187 D.t1119 G.t4187 S.t417 S.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4188 S.t416 G.t4188 D.t653 S.t270 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4189 D.t697 G.t4189 S.t415 S.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4190 D.t922 G.t4190 S.t414 S.t321 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4191 D.t847 G.t4191 S.t413 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4192 D.t827 G.t4192 S.t412 S.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4193 D.t601 G.t4193 S.t411 S.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4194 D.t594 G.t4194 S.t410 S.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4195 D.t530 G.t4195 S.t409 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4196 D.t2080 G.t4196 S.t408 S.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4197 S.t407 G.t4197 D.t124 S.t406 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4198 S.t405 G.t4198 D.t2750 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4199 D.t2753 G.t4199 S.t404 S.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4200 S.t403 G.t4200 D.t3741 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4201 D.t3745 G.t4201 S.t402 S.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4202 D.t4094 G.t4202 S.t401 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4203 S.t400 G.t4203 D.t3288 S.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4204 D.t3906 G.t4204 S.t399 S.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4205 S.t398 G.t4205 D.t3724 S.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4206 S.t397 G.t4206 D.t3506 S.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4207 D.t3539 G.t4207 S.t396 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4208 S.t395 G.t4208 D.t3334 S.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4209 S.t394 G.t4209 D.t4108 S.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4210 S.t393 G.t4210 D.t264 S.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4211 D.t3663 G.t4211 S.t392 S.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4212 D.t3475 G.t4212 S.t391 S.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4213 D.t3228 G.t4213 S.t390 S.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4214 D.t3337 G.t4214 S.t389 S.t388 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4215 D.t3931 G.t4215 S.t387 S.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4216 D.t3918 G.t4216 S.t386 S.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4217 D.t3497 G.t4217 S.t385 S.t270 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4218 D.t3439 G.t4218 S.t384 S.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4219 S.t383 G.t4219 D.t3562 S.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4220 D.t3747 G.t4220 S.t382 S.t209 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4221 D.t3839 G.t4221 S.t381 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4222 S.t380 G.t4222 D.t3837 S.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4223 D.t3268 G.t4223 S.t379 S.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4224 S.t378 G.t4224 D.t3829 S.t150 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4225 S.t377 G.t4225 D.t3414 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4226 D.t3693 G.t4226 S.t376 S.t231 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4227 D.t3961 G.t4227 S.t375 S.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4228 S.t374 G.t4228 D.t3753 S.t150 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4229 S.t373 G.t4229 D.t3836 S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4230 S.t372 G.t4230 D.t3959 S.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4231 D.t370 G.t4231 S.t371 S.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4232 D.t245 G.t4232 S.t370 S.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4233 S.t369 G.t4233 D.t148 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4234 D.t237 G.t4234 S.t368 S.t218 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4235 D.t233 G.t4235 S.t367 S.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4236 S.t365 G.t4236 D.t126 S.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4237 D.t116 G.t4237 S.t364 S.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4238 S.t363 G.t4238 D.t134 S.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4239 D.t146 G.t4239 S.t362 S.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4240 D.t147 G.t4240 S.t361 S.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4241 D.t149 G.t4241 S.t360 S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4242 D.t151 G.t4242 S.t359 S.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4243 D.t152 G.t4243 S.t358 S.t357 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4244 S.t356 G.t4244 D.t169 S.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4245 S.t355 G.t4245 D.t172 S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4246 S.t354 G.t4246 D.t170 S.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4247 S.t353 G.t4247 D.t171 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4248 D.t173 G.t4248 S.t352 S.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4249 S.t351 G.t4249 D.t1049 S.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4250 S.t350 G.t4250 D.t177 S.t198 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4251 D.t2588 G.t4251 S.t349 S.t176 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4252 D.t193 G.t4252 S.t348 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4253 D.t256 G.t4253 S.t347 S.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4254 D.t257 G.t4254 S.t346 S.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4255 S.t345 G.t4255 D.t258 S.t183 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4256 S.t344 G.t4256 D.t263 S.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4257 S.t343 G.t4257 D.t265 S.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4258 D.t287 G.t4258 S.t342 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4259 D.t288 G.t4259 S.t341 S.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4260 D.t41 G.t4260 S.t340 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4261 D.t42 G.t4261 S.t339 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4262 S.t338 G.t4262 D.t43 S.t270 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4263 S.t337 G.t4263 D.t44 S.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4264 S.t336 G.t4264 D.t45 S.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4265 D.t28 G.t4265 S.t335 S.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4266 S.t334 G.t4266 D.t73 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4267 S.t333 G.t4267 D.t3205 S.t332 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4268 D.t3178 G.t4268 S.t331 S.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4269 D.t9 G.t4269 S.t329 S.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4270 D.t18 G.t4270 S.t328 S.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4271 D.t2564 G.t4271 S.t327 S.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4272 D.t2565 G.t4272 S.t326 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4273 S.t325 G.t4273 D.t2 S.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4274 S.t324 G.t4274 D.t24 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4275 S.t323 G.t4275 D.t26 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4276 D.t3202 G.t4276 S.t322 S.t321 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4277 S.t320 G.t4277 D.t297 S.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4278 D.t305 G.t4278 S.t319 S.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4279 S.t318 G.t4279 D.t309 S.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4280 S.t317 G.t4280 D.t312 S.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4281 D.t2045 G.t4281 S.t316 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4282 D.t323 G.t4282 S.t315 S.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4283 D.t1362 G.t4283 S.t314 S.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4284 S.t313 G.t4284 D.t2144 S.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4285 S.t312 G.t4285 D.t1741 S.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4286 D.t1001 G.t4286 S.t311 S.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4287 D.t136 G.t4287 S.t310 S.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4288 S.t309 G.t4288 D.t156 S.t150 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4289 S.t308 G.t4289 D.t2625 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4290 S.t307 G.t4290 D.t2686 S.t139 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4291 D.t2673 G.t4291 S.t306 S.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4292 D.t2674 G.t4292 S.t305 S.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4293 S.t304 G.t4293 D.t2659 S.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4294 S.t303 G.t4294 D.t2623 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4295 S.t302 G.t4295 D.t2662 S.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4296 D.t1651 G.t4296 S.t301 S.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4297 S.t300 G.t4297 D.t1734 S.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4298 S.t299 G.t4298 D.t1956 S.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4299 D.t1941 G.t4299 S.t298 S.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4300 S.t297 G.t4300 D.t1940 S.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4301 D.t1899 G.t4301 S.t296 S.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4302 D.t1883 G.t4302 S.t295 S.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4303 D.t1588 G.t4303 S.t294 S.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4304 S.t293 G.t4304 D.t1544 S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4305 D.t1536 G.t4305 S.t292 S.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4306 S.t291 G.t4306 D.t2041 S.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4307 S.t290 G.t4307 D.t2079 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4308 S.t289 G.t4308 D.t748 S.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4309 D.t1298 G.t4309 S.t287 S.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4310 D.t1673 G.t4310 S.t286 S.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4311 D.t155 G.t4311 S.t285 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4312 D.t2664 G.t4312 S.t284 S.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4313 S.t283 G.t4313 D.t2670 S.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4314 D.t4384 G.t4314 S.t282 S.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4315 D.t398 G.t4315 S.t281 S.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4316 D.t366 G.t4316 S.t280 S.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4317 D.t125 G.t4317 S.t279 S.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4318 S.t278 G.t4318 D.t154 S.t79 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4319 S.t277 G.t4319 D.t3216 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4320 D.t0 G.t4320 S.t276 S.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4321 S.t275 G.t4321 D.t67 S.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4322 D.t89 G.t4322 S.t274 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4323 D.t123 G.t4323 S.t273 S.t176 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4324 D.t86 G.t4324 S.t272 S.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4325 S.t271 G.t4325 D.t96 S.t270 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4326 D.t2749 G.t4326 S.t269 S.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4327 S.t268 G.t4327 D.t90 S.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4328 D.t2744 G.t4328 S.t267 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4329 S.t266 G.t4329 D.t2679 S.t79 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4330 S.t265 G.t4330 D.t2740 S.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4331 D.t3175 G.t4331 S.t264 S.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4332 D.t2743 G.t4332 S.t263 S.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4333 S.t261 G.t4333 D.t2735 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4334 D.t2734 G.t4334 S.t260 S.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4335 D.t2719 G.t4335 S.t259 S.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4336 D.t2715 G.t4336 S.t258 S.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4337 D.t2723 G.t4337 S.t257 S.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4338 S.t256 G.t4338 D.t91 S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4339 D.t2697 G.t4339 S.t255 S.t150 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4340 S.t254 G.t4340 D.t2677 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4341 S.t253 G.t4341 D.t2681 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4342 D.t2849 G.t4342 S.t252 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4343 S.t251 G.t4343 D.t2602 S.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4344 D.t991 G.t4344 S.t250 S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4345 S.t249 G.t4345 D.t1954 S.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4346 S.t248 G.t4346 D.t1620 S.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4347 S.t247 G.t4347 D.t1605 S.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4348 S.t246 G.t4348 D.t1560 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4349 D.t1304 G.t4349 S.t245 S.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4350 S.t244 G.t4350 D.t2081 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4351 D.t604 G.t4351 S.t243 S.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4352 D.t575 G.t4352 S.t242 S.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4353 D.t1320 G.t4353 S.t241 S.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4354 S.t240 G.t4354 D.t1317 S.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4355 S.t239 G.t4355 D.t1312 S.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4356 D.t1295 G.t4356 S.t238 S.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4357 D.t1300 G.t4357 S.t237 S.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4358 S.t236 G.t4358 D.t1357 S.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4359 S.t235 G.t4359 D.t685 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4360 S.t234 G.t4360 D.t514 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4361 D.t542 G.t4361 S.t233 S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4362 S.t232 G.t4362 D.t614 S.t231 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4363 D.t2737 G.t4363 S.t230 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4364 S.t229 G.t4364 D.t3171 S.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4365 D.t2741 G.t4365 S.t228 S.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4366 D.t2746 G.t4366 S.t227 S.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4367 S.t226 G.t4367 D.t85 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4368 S.t225 G.t4368 D.t109 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4369 S.t224 G.t4369 D.t83 S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4370 S.t223 G.t4370 D.t3253 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4371 S.t222 G.t4371 D.t3577 S.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4372 S.t220 G.t4372 D.t4062 S.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4373 S.t219 G.t4373 D.t3034 S.t218 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4374 S.t217 G.t4374 D.t2705 S.t216 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4375 D.t368 G.t4375 S.t215 S.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4376 S.t213 G.t4376 D.t226 S.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4377 S.t212 G.t4377 D.t130 S.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4378 S.t211 G.t4378 D.t222 S.t158 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4379 S.t210 G.t4379 D.t132 S.t209 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4380 S.t208 G.t4380 D.t159 S.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4381 D.t133 G.t4381 S.t207 S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4382 S.t206 G.t4382 D.t219 S.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4383 D.t175 G.t4383 S.t205 S.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4384 S.t204 G.t4384 D.t164 S.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4385 D.t137 G.t4385 S.t203 S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4386 S.t202 G.t4386 D.t143 S.t79 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4387 D.t165 G.t4387 S.t201 S.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4388 S.t199 G.t4388 D.t168 S.t198 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4389 D.t184 G.t4389 S.t197 S.t176 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4390 S.t196 G.t4390 D.t215 S.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4391 S.t195 G.t4391 D.t260 S.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4392 D.t262 G.t4392 S.t194 S.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4393 S.t192 G.t4393 D.t36 S.t183 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4394 D.t35 G.t4394 S.t191 S.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4395 S.t190 G.t4395 D.t34 S.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4396 S.t189 G.t4396 D.t30 S.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4397 D.t29 G.t4397 S.t188 S.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4398 S.t186 G.t4398 D.t2297 S.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4399 D.t2292 G.t4399 S.t185 S.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4400 D.t2082 G.t4400 S.t184 S.t183 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4401 S.t182 G.t4401 D.t3193 S.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4402 S.t180 G.t4402 D.t3199 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4403 D.t3201 G.t4403 S.t179 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4404 D.t3204 G.t4404 S.t178 S.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4405 S.t177 G.t4405 D.t3206 S.t176 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4406 D.t2563 G.t4406 S.t175 S.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4407 D.t80 G.t4407 S.t173 S.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4408 S.t171 G.t4408 D.t97 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4409 S.t170 G.t4409 D.t104 S.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4410 S.t168 G.t4410 D.t359 S.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4411 D.t332 G.t4411 S.t166 S.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4412 D.t122 G.t4412 S.t164 S.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4413 D.t2747 G.t4413 S.t162 S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4414 S.t161 G.t4414 D.t2693 S.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4415 S.t159 G.t4415 D.t2691 S.t158 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4416 S.t157 G.t4416 D.t2724 S.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4417 D.t2739 G.t4417 S.t156 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4418 S.t155 G.t4418 D.t2729 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4419 D.t2596 G.t4419 S.t154 S.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4420 D.t2742 G.t4420 S.t153 S.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4421 S.t151 G.t4421 D.t2626 S.t150 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4422 D.t2667 G.t4422 S.t149 S.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4423 S.t147 G.t4423 D.t2682 S.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4424 D.t2678 G.t4424 S.t146 S.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4425 S.t145 G.t4425 D.t2683 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4426 D.t2628 G.t4426 S.t144 S.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4427 D.t1305 G.t4427 S.t142 S.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4428 S.t140 G.t4428 D.t1939 S.t139 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4429 S.t138 G.t4429 D.t1999 S.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4430 S.t136 G.t4430 D.t1541 S.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4431 S.t135 G.t4431 D.t1190 S.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4432 D.t1584 G.t4432 S.t133 S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4433 D.t1587 G.t4433 S.t132 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4434 S.t131 G.t4434 D.t1670 S.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4435 D.t1702 G.t4435 S.t129 S.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4436 S.t127 G.t4436 D.t623 S.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4437 D.t1126 G.t4437 S.t125 S.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4438 S.t124 G.t4438 D.t1130 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4439 S.t123 G.t4439 D.t1508 S.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4440 S.t121 G.t4440 D.t1216 S.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4441 S.t120 G.t4441 D.t968 S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4442 D.t814 G.t4442 S.t119 S.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4443 D.t862 G.t4443 S.t117 S.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4444 S.t115 G.t4444 D.t882 S.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4445 S.t113 G.t4445 D.t907 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4446 S.t112 G.t4446 D.t2042 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4447 D.t2717 G.t4447 S.t111 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4448 S.t110 G.t4448 D.t376 S.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4449 S.t108 G.t4449 D.t628 S.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4450 D.t745 G.t4450 S.t107 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4451 D.t749 G.t4451 S.t106 S.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4452 D.t2745 G.t4452 S.t104 S.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4453 S.t103 G.t4453 D.t100 S.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4454 D.t2718 G.t4454 S.t101 S.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4455 S.t99 G.t4455 D.t367 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4456 D.t2765 G.t4456 S.t98 S.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4457 D.t2923 G.t4457 S.t96 S.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4458 S.t94 G.t4458 D.t2814 S.t79 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4459 D.t2784 G.t4459 S.t93 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4460 S.t92 G.t4460 D.t2967 S.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4461 S.t90 G.t4461 D.t2903 S.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4462 D.t2751 G.t4462 S.t89 S.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4463 S.t87 G.t4463 D.t1549 S.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4464 S.t86 G.t4464 D.t2762 S.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4465 S.t85 G.t4465 D.t3074 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4466 S.t84 G.t4466 D.t2760 S.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4467 S.t82 G.t4467 D.t2707 S.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4468 S.t80 G.t4468 D.t1225 S.t79 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4469 D.t1337 G.t4469 S.t78 S.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4470 S.t76 G.t4470 D.t901 S.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4471 S.t74 G.t4471 D.t501 S.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4472 D.t1592 G.t4472 S.t72 S.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4473 D.t2040 G.t4473 S.t71 S.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4474 S.t69 G.t4474 D.t1548 S.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4475 S.t68 G.t4475 D.t1562 S.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4476 S.t66 G.t4476 D.t2100 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4477 S.t65 G.t4477 D.t1655 S.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4478 D.t1261 G.t4478 S.t63 S.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4479 S.t61 G.t4479 D.t1966 S.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4480 S.t59 G.t4480 D.t1979 S.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4481 D.t2013 G.t4481 S.t57 S.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4482 D.t1591 G.t4482 S.t55 S.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4483 S.t53 G.t4483 D.t1716 S.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4484 S.t52 G.t4484 D.t1708 S.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4485 S.t50 G.t4485 D.t1184 S.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4486 D.t1550 G.t4486 S.t48 S.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4487 S.t46 G.t4487 D.t1637 S.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4488 S.t44 G.t4488 D.t1589 S.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4489 D.t1547 G.t4489 S.t42 S.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4490 S.t40 G.t4490 D.t2130 S.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4491 S.t38 G.t4491 D.t2266 S.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4492 S.t36 G.t4492 D.t2097 S.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4493 S.t34 G.t4493 D.t2114 S.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4494 S.t32 G.t4494 D.t2239 S.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4495 D.t1262 G.t4495 S.t30 S.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4496 S.t28 G.t4496 D.t1157 S.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4497 S.t26 G.t4497 D.t1164 S.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4498 D.t1115 G.t4498 S.t24 S.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4499 S.t22 G.t4499 D.t854 S.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4500 D.t969 G.t4500 S.t20 S.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4501 S.t18 G.t4501 D.t1359 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4502 S.t17 G.t4502 D.t2713 S.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4503 S.t15 G.t4503 D.t684 S.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4504 D.t970 G.t4504 S.t13 S.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4505 S.t12 G.t4505 D.t895 S.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4506 S.t10 G.t4506 D.t828 S.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4507 D.t663 G.t4507 S.t8 S.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4508 S.t6 G.t4508 D.t2706 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4509 S.t5 G.t4509 D.t2695 S.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4510 S.t3 G.t4510 D.t490 S.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4511 S.t1 G.t4511 D.t574 S.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
R0 G.n2306 G.t2035 132.223
R1 G.n3565 G.t1815 132.223
R2 G.n3569 G.t496 132.223
R3 G.n2309 G.t672 132.223
R4 G.n2313 G.t3349 132.223
R5 G.n3576 G.t680 132.223
R6 G.n3586 G.t3746 132.223
R7 G.n2320 G.t1920 132.223
R8 G.n2327 G.t1784 132.223
R9 G.n3599 G.t3648 132.223
R10 G.n3615 G.t2197 132.223
R11 G.n2337 G.t369 132.223
R12 G.n2347 G.t230 132.223
R13 G.n3634 G.t2098 132.223
R14 G.n3656 G.t661 132.223
R15 G.n2360 G.t3319 132.223
R16 G.n2375 G.t3176 132.223
R17 G.n3681 G.t557 132.223
R18 G.n3706 G.t3628 132.223
R19 G.n2391 G.t1755 132.223
R20 G.n2410 G.t1616 132.223
R21 G.n3734 G.t3523 132.223
R22 G.n3765 G.t2262 132.223
R23 G.n2429 G.t456 132.223
R24 G.n2451 G.t55 132.223
R25 G.n3799 G.t1964 132.223
R26 G.n3836 G.t729 132.223
R27 G.n2473 G.t3410 132.223
R28 G.n2498 G.t3012 132.223
R29 G.n3876 G.t415 132.223
R30 G.n3919 G.t3691 132.223
R31 G.n2525 G.t1851 132.223
R32 G.n2553 G.t1457 132.223
R33 G.n3965 G.t3370 132.223
R34 G.n4011 G.t2146 132.223
R35 G.n2583 G.t292 132.223
R36 G.n2614 G.t4415 132.223
R37 G.n4060 G.t1807 132.223
R38 G.n4112 G.t3232 132.223
R39 G.n2648 G.t1877 132.223
R40 G.n2682 G.t1480 132.223
R41 G.n4167 G.t2864 132.223
R42 G.n4225 G.t1667 132.223
R43 G.n2719 G.t319 132.223
R44 G.n2756 G.t180 132.223
R45 G.n4286 G.t1536 132.223
R46 G.n4350 G.t111 132.223
R47 G.n2796 G.t3268 132.223
R48 G.n2838 G.t3126 132.223
R49 G.n4417 G.t4489 132.223
R50 G.n4487 G.t3060 132.223
R51 G.n2881 G.t1701 132.223
R52 G.n2927 G.t1568 132.223
R53 G.n4557 G.t2935 132.223
R54 G.n4630 G.t1507 132.223
R55 G.n2973 G.t147 132.223
R56 G.n3022 G.t8 132.223
R57 G.n4706 G.t1385 132.223
R58 G.n4784 G.t4461 132.223
R59 G.n3070 G.t3092 132.223
R60 G.n3115 G.t2962 132.223
R61 G.n4856 G.t4352 132.223
R62 G.n4925 G.t3153 132.223
R63 G.n3158 G.t1796 132.223
R64 G.n3198 G.t1414 132.223
R65 G.n4988 G.t2796 132.223
R66 G.n5048 G.t1592 132.223
R67 G.n3235 G.t243 132.223
R68 G.n3270 G.t4378 132.223
R69 G.n5102 G.t1251 132.223
R70 G.n5153 G.t33 132.223
R71 G.n3302 G.t3191 132.223
R72 G.n3332 G.t2827 132.223
R73 G.n5200 G.t4211 132.223
R74 G.n5242 G.t896 132.223
R75 G.n3359 G.t4041 132.223
R76 G.n3383 G.t3698 132.223
R77 G.n5280 G.t588 132.223
R78 G.n5313 G.t3853 132.223
R79 G.n3404 G.t2474 132.223
R80 G.n3422 G.t2153 132.223
R81 G.n5343 G.t3555 132.223
R82 G.n5367 G.t2294 132.223
R83 G.n3437 G.t927 132.223
R84 G.n3449 G.t808 132.223
R85 G.n5388 G.t2193 132.223
R86 G.n5415 G.t655 132.223
R87 G.n5403 G.t757 132.223
R88 G.n3458 G.t3887 132.223
R89 G.n3465 G.t3770 132.223
R90 G.n5424 G.t3620 132.223
R91 G.n5421 G.t3718 132.223
R92 G.n3469 G.t2323 132.223
R93 G.n3470 G.t2216 132.223
R94 G.n2300 G.t2135 132.208
R95 G.n2291 G.t4429 132.208
R96 G.n2277 G.t44 132.208
R97 G.n2257 G.t2367 132.208
R98 G.n2233 G.t2491 132.208
R99 G.n2203 G.t350 132.208
R100 G.n2168 G.t478 132.208
R101 G.n2127 G.t3886 132.208
R102 G.n2082 G.t2873 132.208
R103 G.n2031 G.t331 132.208
R104 G.n1974 G.t3789 132.208
R105 G.n1912 G.t2741 132.208
R106 G.n1844 G.t1744 132.208
R107 G.n1772 G.t695 132.208
R108 G.n1694 G.t4180 132.208
R109 G.n1611 G.t3123 132.208
R110 G.n1524 G.t2129 132.208
R111 G.n1436 G.t1065 132.208
R112 G.n1348 G.t1184 132.208
R113 G.n1260 G.t3549 132.208
R114 G.n1172 G.t3646 132.208
R115 G.n1084 G.t1427 132.208
R116 G.n999 G.t1552 132.208
R117 G.n917 G.t3880 132.208
R118 G.n841 G.t4002 132.208
R119 G.n768 G.t1855 132.208
R120 G.n698 G.t1979 132.208
R121 G.n631 G.t1006 132.208
R122 G.n567 G.t4495 132.208
R123 G.n506 G.t3498 132.208
R124 G.n448 G.t2426 132.208
R125 G.n393 G.t1379 132.208
R126 G.n344 G.t417 132.208
R127 G.n298 G.t3824 132.208
R128 G.n255 G.t2820 132.208
R129 G.n215 G.t1792 132.208
R130 G.n178 G.t759 132.208
R131 G.n144 G.t4224 132.208
R132 G.n113 G.t4332 132.208
R133 G.n88 G.t2167 132.208
R134 G.n66 G.t2257 132.208
R135 G.n47 G.t80 132.208
R136 G.n31 G.t224 132.208
R137 G.n18 G.t2526 132.208
R138 G.n8 G.t1139 132.208
R139 G.n1 G.t610 132.208
R140 G.n3567 G.t3753 132.208
R141 G.n5 G.t4300 132.208
R142 G.n15 G.t1200 132.208
R143 G.n28 G.t3418 132.208
R144 G.n44 G.t3282 132.208
R145 G.n63 G.t925 132.208
R146 G.n85 G.t809 132.208
R147 G.n110 G.t2985 132.208
R148 G.n141 G.t2872 132.208
R149 G.n175 G.t3924 132.208
R150 G.n212 G.t475 132.208
R151 G.n252 G.t1467 132.208
R152 G.n295 G.t2490 132.208
R153 G.n341 G.t3577 132.208
R154 G.n390 G.t43 132.208
R155 G.n445 G.t1110 132.208
R156 G.n503 G.t2134 132.208
R157 G.n564 G.t3173 132.208
R158 G.n628 G.t4186 132.208
R159 G.n695 G.t625 132.208
R160 G.n765 G.t525 132.208
R161 G.n838 G.t2668 132.208
R162 G.n914 G.t2542 132.208
R163 G.n996 G.t239 132.208
R164 G.n1081 G.t98 132.208
R165 G.n1169 G.t2270 132.208
R166 G.n1257 G.t2176 132.208
R167 G.n1345 G.t4345 132.208
R168 G.n1433 G.t4235 132.208
R169 G.n1521 G.t769 132.208
R170 G.n1608 G.t1812 132.208
R171 G.n1691 G.t2830 132.208
R172 G.n1769 G.t3840 132.208
R173 G.n1841 G.t431 132.208
R174 G.n1909 G.t1392 132.208
R175 G.n1971 G.t2444 132.208
R176 G.n2028 G.t3510 132.208
R177 G.n2079 G.t1533 132.208
R178 G.n2124 G.t2548 132.208
R179 G.n2165 G.t3627 132.208
R180 G.n2200 G.t3525 132.208
R181 G.n2230 G.t1164 132.208
R182 G.n2254 G.t1039 132.208
R183 G.n2274 G.t3241 132.208
R184 G.n2288 G.t3096 132.208
R185 G.n2297 G.t776 132.208
R186 G.n2311 G.t524 132.208
R187 G.n2285 G.t344 132.208
R188 G.n2271 G.t2023 132.208
R189 G.n2251 G.t1849 132.208
R190 G.n2227 G.t3536 132.208
R191 G.n2197 G.t3356 132.208
R192 G.n2162 G.t531 132.208
R193 G.n2121 G.t3332 132.208
R194 G.n2076 G.t2030 132.208
R195 G.n2025 G.t802 132.208
R196 G.n1968 G.t4012 132.208
R197 G.n1906 G.t2299 132.208
R198 G.n1838 G.t1003 132.208
R199 G.n1766 G.t3808 132.208
R200 G.n1688 G.t2510 132.208
R201 G.n1605 G.t811 132.208
R202 G.n1518 G.t4021 132.208
R203 G.n1430 G.t2302 132.208
R204 G.n1342 G.t3992 132.208
R205 G.n1254 G.t3815 132.208
R206 G.n1166 G.t984 132.208
R207 G.n1078 G.t820 132.208
R208 G.n993 G.t2493 132.208
R209 G.n911 G.t2315 132.208
R210 G.n835 G.t4005 132.208
R211 G.n762 G.t3823 132.208
R212 G.n692 G.t993 132.208
R213 G.n625 G.t159 132.208
R214 G.n561 G.t3398 132.208
R215 G.n500 G.t1663 132.208
R216 G.n442 G.t395 132.208
R217 G.n387 G.t3172 132.208
R218 G.n338 G.t1899 132.208
R219 G.n292 G.t166 132.208
R220 G.n249 G.t3409 132.208
R221 G.n209 G.t1672 132.208
R222 G.n172 G.t402 132.208
R223 G.n138 G.t3183 132.208
R224 G.n107 G.t382 132.208
R225 G.n82 G.t183 132.208
R226 G.n60 G.t1882 132.208
R227 G.n41 G.t1683 132.208
R228 G.n25 G.t3393 132.208
R229 G.n12 G.t3193 132.208
R230 G.n3572 G.t2040 132.208
R231 G.n3574 G.t349 132.208
R232 G.n3584 G.t3436 132.208
R233 G.n3582 G.t602 132.208
R234 G.n3580 G.t1770 132.208
R235 G.n22 G.t1961 132.208
R236 G.n38 G.t270 132.208
R237 G.n57 G.t461 132.208
R238 G.n79 G.t3272 132.208
R239 G.n104 G.t3464 132.208
R240 G.n135 G.t1759 132.208
R241 G.n169 G.t3487 132.208
R242 G.n206 G.t261 132.208
R243 G.n246 G.t1978 132.208
R244 G.n289 G.t3261 132.208
R245 G.n335 G.t477 132.208
R246 G.n384 G.t1752 132.208
R247 G.n439 G.t3480 132.208
R248 G.n497 G.t253 132.208
R249 G.n558 G.t1968 132.208
R250 G.n622 G.t3254 132.208
R251 G.n689 G.t4088 132.208
R252 G.n759 G.t2387 132.208
R253 G.n832 G.t2576 132.208
R254 G.n908 G.t893 132.208
R255 G.n990 G.t1078 132.208
R256 G.n1075 G.t3900 132.208
R257 G.n1163 G.t4079 132.208
R258 G.n1251 G.t2379 132.208
R259 G.n1339 G.t2566 132.208
R260 G.n1427 G.t884 132.208
R261 G.n1515 G.t2588 132.208
R262 G.n1602 G.t3889 132.208
R263 G.n1685 G.t1091 132.208
R264 G.n1763 G.t2374 132.208
R265 G.n1835 G.t4096 132.208
R266 G.n1903 G.t875 132.208
R267 G.n1965 G.t2584 132.208
R268 G.n2022 G.t3883 132.208
R269 G.n2073 G.t597 132.208
R270 G.n2118 G.t1907 132.208
R271 G.n2159 G.t3600 132.208
R272 G.n2194 G.t1930 132.208
R273 G.n2224 G.t2090 132.208
R274 G.n2248 G.t428 132.208
R275 G.n2268 G.t591 132.208
R276 G.n2316 G.t3431 132.208
R277 G.n2318 G.t3593 132.208
R278 G.n2325 G.t3484 132.208
R279 G.n2323 G.t3294 132.208
R280 G.n2265 G.t480 132.208
R281 G.n2245 G.t293 132.208
R282 G.n2221 G.t1983 132.208
R283 G.n2191 G.t1793 132.208
R284 G.n2156 G.t3491 132.208
R285 G.n2115 G.t1763 132.208
R286 G.n2070 G.t488 132.208
R287 G.n2019 G.t3764 132.208
R288 G.n1962 G.t2450 132.208
R289 G.n1900 G.t762 132.208
R290 G.n1832 G.t3958 132.208
R291 G.n1760 G.t2253 132.208
R292 G.n1682 G.t961 132.208
R293 G.n1599 G.t3774 132.208
R294 G.n1512 G.t2458 132.208
R295 G.n1424 G.t767 132.208
R296 G.n1336 G.t2431 132.208
R297 G.n1248 G.t2261 132.208
R298 G.n1160 G.t3942 132.208
R299 G.n1072 G.t3783 132.208
R300 G.n987 G.t944 132.208
R301 G.n905 G.t777 132.208
R302 G.n829 G.t2446 132.208
R303 G.n756 G.t2271 132.208
R304 G.n686 G.t3953 132.208
R305 G.n619 G.t3109 132.208
R306 G.n555 G.t1838 132.208
R307 G.n494 G.t106 132.208
R308 G.n436 G.t3350 132.208
R309 G.n381 G.t1612 132.208
R310 G.n332 G.t345 132.208
R311 G.n286 G.t3116 132.208
R312 G.n243 G.t1850 132.208
R313 G.n203 G.t120 132.208
R314 G.n166 G.t3357 132.208
R315 G.n132 G.t1622 132.208
R316 G.n101 G.t3333 132.208
R317 G.n76 G.t3133 132.208
R318 G.n54 G.t328 132.208
R319 G.n35 G.t129 132.208
R320 G.n3591 G.t1833 132.208
R321 G.n3593 G.t1627 132.208
R322 G.n3595 G.t498 132.208
R323 G.n3597 G.t3299 132.208
R324 G.n3613 G.t1878 132.208
R325 G.n3611 G.t3567 132.208
R326 G.n3609 G.t215 132.208
R327 G.n3607 G.t413 132.208
R328 G.n3605 G.t3221 132.208
R329 G.n51 G.t3419 132.208
R330 G.n73 G.t1707 132.208
R331 G.n98 G.t1908 132.208
R332 G.n129 G.t207 132.208
R333 G.n163 G.t1931 132.208
R334 G.n200 G.t3211 132.208
R335 G.n240 G.t429 132.208
R336 G.n283 G.t1697 132.208
R337 G.n329 G.t3432 132.208
R338 G.n378 G.t199 132.208
R339 G.n433 G.t1921 132.208
R340 G.n491 G.t3201 132.208
R341 G.n552 G.t418 132.208
R342 G.n616 G.t1689 132.208
R343 G.n683 G.t2523 132.208
R344 G.n753 G.t844 132.208
R345 G.n826 G.t1024 132.208
R346 G.n902 G.t3848 132.208
R347 G.n984 G.t4030 132.208
R348 G.n1069 G.t2336 132.208
R349 G.n1157 G.t2514 132.208
R350 G.n1245 G.t835 132.208
R351 G.n1333 G.t1011 132.208
R352 G.n1421 G.t3838 132.208
R353 G.n1509 G.t1040 132.208
R354 G.n1596 G.t2326 132.208
R355 G.n1679 G.t4047 132.208
R356 G.n1757 G.t829 132.208
R357 G.n1829 G.t2532 132.208
R358 G.n1897 G.t3832 132.208
R359 G.n1959 G.t1033 132.208
R360 G.n2016 G.t2320 132.208
R361 G.n2067 G.t3565 132.208
R362 G.n2112 G.t357 132.208
R363 G.n2153 G.t2052 132.208
R364 G.n2188 G.t378 132.208
R365 G.n2218 G.t549 132.208
R366 G.n2242 G.t3379 132.208
R367 G.n2331 G.t3559 132.208
R368 G.n2333 G.t1871 132.208
R369 G.n2335 G.t2046 132.208
R370 G.n2345 G.t1927 132.208
R371 G.n2343 G.t1727 132.208
R372 G.n2341 G.t3438 132.208
R373 G.n2239 G.t3242 132.208
R374 G.n2215 G.t434 132.208
R375 G.n2185 G.t240 132.208
R376 G.n2150 G.t1936 132.208
R377 G.n2109 G.t208 132.208
R378 G.n2064 G.t3442 132.208
R379 G.n2013 G.t2211 132.208
R380 G.n1956 G.t903 132.208
R381 G.n1894 G.t3723 132.208
R382 G.n1826 G.t2396 132.208
R383 G.n1754 G.t716 132.208
R384 G.n1676 G.t3916 132.208
R385 G.n1593 G.t2218 132.208
R386 G.n1506 G.t911 132.208
R387 G.n1418 G.t3730 132.208
R388 G.n1330 G.t887 132.208
R389 G.n1242 G.t726 132.208
R390 G.n1154 G.t2382 132.208
R391 G.n1066 G.t2227 132.208
R392 G.n981 G.t3905 132.208
R393 G.n899 G.t3738 132.208
R394 G.n823 G.t900 132.208
R395 G.n750 G.t733 132.208
R396 G.n680 G.t2392 132.208
R397 G.n613 G.t1556 132.208
R398 G.n549 G.t282 132.208
R399 G.n488 G.t3055 132.208
R400 G.n430 G.t1785 132.208
R401 G.n375 G.t54 132.208
R402 G.n326 G.t3295 132.208
R403 G.n280 G.t1561 132.208
R404 G.n237 G.t294 132.208
R405 G.n197 G.t3065 132.208
R406 G.n160 G.t1794 132.208
R407 G.n126 G.t62 132.208
R408 G.n95 G.t1765 132.208
R409 G.n70 G.t1574 132.208
R410 G.n3622 G.t3279 132.208
R411 G.n3624 G.t3074 132.208
R412 G.n3626 G.t278 132.208
R413 G.n3628 G.t67 132.208
R414 G.n3630 G.t3451 132.208
R415 G.n3632 G.t1732 132.208
R416 G.n3654 G.t321 132.208
R417 G.n3652 G.t2014 132.208
R418 G.n3650 G.t3164 132.208
R419 G.n3648 G.t3368 132.208
R420 G.n3646 G.t1656 132.208
R421 G.n3644 G.t1860 132.208
R422 G.n3642 G.t151 132.208
R423 G.n92 G.t358 132.208
R424 G.n123 G.t3155 132.208
R425 G.n157 G.t379 132.208
R426 G.n194 G.t1643 132.208
R427 G.n234 G.t3380 132.208
R428 G.n277 G.t141 132.208
R429 G.n323 G.t1872 132.208
R430 G.n372 G.t3147 132.208
R431 G.n427 G.t370 132.208
R432 G.n485 G.t1633 132.208
R433 G.n546 G.t3371 132.208
R434 G.n610 G.t134 132.208
R435 G.n677 G.t970 132.208
R436 G.n747 G.t3800 132.208
R437 G.n820 G.t3975 132.208
R438 G.n896 G.t2288 132.208
R439 G.n978 G.t2466 132.208
R440 G.n1063 G.t798 132.208
R441 G.n1151 G.t963 132.208
R442 G.n1239 G.t3796 132.208
R443 G.n1327 G.t3964 132.208
R444 G.n1415 G.t2283 132.208
R445 G.n1503 G.t3990 132.208
R446 G.n1590 G.t787 132.208
R447 G.n1673 G.t2479 132.208
R448 G.n1751 G.t3790 132.208
R449 G.n1823 G.t977 132.208
R450 G.n1891 G.t2276 132.208
R451 G.n1953 G.t3984 132.208
R452 G.n2010 G.t782 132.208
R453 G.n2061 G.t2012 132.208
R454 G.n2106 G.t3306 132.208
R455 G.n2147 G.t511 132.208
R456 G.n2182 G.t3328 132.208
R457 G.n2212 G.t3514 132.208
R458 G.n2352 G.t1819 132.208
R459 G.n2354 G.t2005 132.208
R460 G.n2356 G.t313 132.208
R461 G.n2358 G.t504 132.208
R462 G.n2373 G.t374 132.208
R463 G.n2371 G.t171 132.208
R464 G.n2369 G.t1879 132.208
R465 G.n2367 G.t1677 132.208
R466 G.n2209 G.t3384 132.208
R467 G.n2179 G.t3186 132.208
R468 G.n2144 G.t384 132.208
R469 G.n2103 G.t3160 132.208
R470 G.n2058 G.t1886 132.208
R471 G.n2007 G.t674 132.208
R472 G.n1950 G.t3863 132.208
R473 G.n1888 G.t2180 132.208
R474 G.n1820 G.t859 132.208
R475 G.n1748 G.t3681 132.208
R476 G.n1670 G.t2360 132.208
R477 G.n1587 G.t678 132.208
R478 G.n1500 G.t3867 132.208
R479 G.n1412 G.t2183 132.208
R480 G.n1324 G.t3844 132.208
R481 G.n1236 G.t3689 132.208
R482 G.n1148 G.t839 132.208
R483 G.n1060 G.t691 132.208
R484 G.n975 G.t2343 132.208
R485 G.n893 G.t2190 132.208
R486 G.n817 G.t3856 132.208
R487 G.n744 G.t3696 132.208
R488 G.n674 G.t849 132.208
R489 G.n607 G.t4511 132.208
R490 G.n543 G.t3230 132.208
R491 G.n482 G.t1502 132.208
R492 G.n424 G.t231 132.208
R493 G.n369 G.t3009 132.208
R494 G.n320 G.t1728 132.208
R495 G.n274 G.t2 132.208
R496 G.n231 G.t3243 132.208
R497 G.n191 G.t1514 132.208
R498 G.n154 G.t241 132.208
R499 G.n120 G.t3019 132.208
R500 G.n3665 G.t210 132.208
R501 G.n3667 G.t17 132.208
R502 G.n3669 G.t1713 132.208
R503 G.n3671 G.t1520 132.208
R504 G.n3673 G.t3225 132.208
R505 G.n3675 G.t3022 132.208
R506 G.n3677 G.t1890 132.208
R507 G.n3679 G.t177 132.208
R508 G.n3704 G.t3269 132.208
R509 G.n3702 G.t469 132.208
R510 G.n3700 G.t1605 132.208
R511 G.n3698 G.t1803 132.208
R512 G.n3696 G.t100 132.208
R513 G.n3694 G.t303 132.208
R514 G.n3692 G.t3098 132.208
R515 G.n3690 G.t3307 132.208
R516 G.n117 G.t1594 132.208
R517 G.n151 G.t3329 132.208
R518 G.n188 G.t86 132.208
R519 G.n228 G.t1820 132.208
R520 G.n271 G.t3086 132.208
R521 G.n317 G.t314 132.208
R522 G.n366 G.t1587 132.208
R523 G.n421 G.t3320 132.208
R524 G.n479 G.t73 132.208
R525 G.n540 G.t1809 132.208
R526 G.n604 G.t3079 132.208
R527 G.n671 G.t3931 132.208
R528 G.n741 G.t2246 132.208
R529 G.n814 G.t2413 132.208
R530 G.n890 G.t754 132.208
R531 G.n972 G.t921 132.208
R532 G.n1057 G.t3759 132.208
R533 G.n1145 G.t3926 132.208
R534 G.n1233 G.t2242 132.208
R535 G.n1321 G.t2406 132.208
R536 G.n1409 G.t747 132.208
R537 G.n1497 G.t2429 132.208
R538 G.n1584 G.t3747 132.208
R539 G.n1667 G.t933 132.208
R540 G.n1745 G.t2234 132.208
R541 G.n1817 G.t3937 132.208
R542 G.n1885 G.t738 132.208
R543 G.n1947 G.t2423 132.208
R544 G.n2004 G.t3741 132.208
R545 G.n2055 G.t464 132.208
R546 G.n2100 G.t1738 132.208
R547 G.n2141 G.t3467 132.208
R548 G.n2176 G.t1760 132.208
R549 G.n2381 G.t1952 132.208
R550 G.n2383 G.t262 132.208
R551 G.n2385 G.t455 132.208
R552 G.n2387 G.t3262 132.208
R553 G.n2389 G.t3457 132.208
R554 G.n2408 G.t3325 132.208
R555 G.n2406 G.t3119 132.208
R556 G.n2404 G.t322 132.208
R557 G.n2402 G.t123 132.208
R558 G.n2400 G.t1824 132.208
R559 G.n2398 G.t1623 132.208
R560 G.n2138 G.t3334 132.208
R561 G.n2097 G.t1597 132.208
R562 G.n2052 G.t332 132.208
R563 G.n2001 G.t3640 132.208
R564 G.n1944 G.t2301 132.208
R565 G.n1882 G.t638 132.208
R566 G.n1814 G.t3812 132.208
R567 G.n1742 G.t2139 132.208
R568 G.n1664 G.t817 132.208
R569 G.n1581 G.t3649 132.208
R570 G.n1494 G.t2307 132.208
R571 G.n1406 G.t646 132.208
R572 G.n1318 G.t2286 132.208
R573 G.n1230 G.t2145 132.208
R574 G.n1142 G.t3798 132.208
R575 G.n1054 G.t3654 132.208
R576 G.n969 G.t801 132.208
R577 G.n887 G.t652 132.208
R578 G.n811 G.t2293 132.208
R579 G.n738 G.t2151 132.208
R580 G.n668 G.t3803 132.208
R581 G.n601 G.t2952 132.208
R582 G.n537 G.t1665 132.208
R583 G.n476 G.t4455 132.208
R584 G.n418 G.t3177 132.208
R585 G.n363 G.t1451 132.208
R586 G.n314 G.t172 132.208
R587 G.n268 G.t2956 132.208
R588 G.n225 G.t1678 132.208
R589 G.n185 G.t4468 132.208
R590 G.n148 G.t3187 132.208
R591 G.n3716 G.t1461 132.208
R592 G.n3718 G.t3161 132.208
R593 G.n3720 G.t2970 132.208
R594 G.n3722 G.t158 132.208
R595 G.n3724 G.t4477 132.208
R596 G.n3726 G.t1661 132.208
R597 G.n3728 G.t1469 132.208
R598 G.n3730 G.t338 132.208
R599 G.n3732 G.t3127 132.208
R600 G.n3763 G.t1959 132.208
R601 G.n3761 G.t3632 132.208
R602 G.n3759 G.t308 132.208
R603 G.n3757 G.t500 132.208
R604 G.n3755 G.t3314 132.208
R605 G.n3753 G.t3500 132.208
R606 G.n3751 G.t1804 132.208
R607 G.n3749 G.t1991 132.208
R608 G.n3747 G.t304 132.208
R609 G.n3745 G.t2013 132.208
R610 G.n182 G.t3308 132.208
R611 G.n222 G.t512 132.208
R612 G.n265 G.t1790 132.208
R613 G.n311 G.t3515 132.208
R614 G.n360 G.t290 132.208
R615 G.n415 G.t2006 132.208
R616 G.n473 G.t3292 132.208
R617 G.n534 G.t505 132.208
R618 G.n598 G.t1780 132.208
R619 G.n665 G.t2610 132.208
R620 G.n735 G.t926 132.208
R621 G.n808 G.t1112 132.208
R622 G.n884 G.t3932 132.208
R623 G.n966 G.t4114 132.208
R624 G.n1051 G.t2414 132.208
R625 G.n1139 G.t2600 132.208
R626 G.n1227 G.t918 132.208
R627 G.n1315 G.t1101 132.208
R628 G.n1403 G.t3921 132.208
R629 G.n1491 G.t1123 132.208
R630 G.n1578 G.t2402 132.208
R631 G.n1661 G.t4131 132.208
R632 G.n1739 G.t908 132.208
R633 G.n1811 G.t2620 132.208
R634 G.n1879 G.t3917 132.208
R635 G.n1941 G.t1119 132.208
R636 G.n1998 G.t2397 132.208
R637 G.n2049 G.t3630 132.208
R638 G.n2094 G.t442 132.208
R639 G.n2135 G.t2120 132.208
R640 G.n2417 G.t465 132.208
R641 G.n2419 G.t617 132.208
R642 G.n2421 G.t3468 132.208
R643 G.n2423 G.t3622 132.208
R644 G.n2425 G.t1953 132.208
R645 G.n2427 G.t2113 132.208
R646 G.n2449 G.t1757 132.208
R647 G.n2447 G.t1562 132.208
R648 G.n2445 G.t3270 132.208
R649 G.n2443 G.t3069 132.208
R650 G.n2441 G.t266 132.208
R651 G.n2439 G.t64 132.208
R652 G.n2437 G.t1766 132.208
R653 G.n2091 G.t39 132.208
R654 G.n2046 G.t3281 132.208
R655 G.n1995 G.t2092 132.208
R656 G.n1938 G.t763 132.208
R657 G.n1876 G.t3601 132.208
R658 G.n1808 G.t2255 132.208
R659 G.n1736 G.t598 132.208
R660 G.n1658 G.t3776 132.208
R661 G.n1575 G.t2099 132.208
R662 G.n1488 G.t770 132.208
R663 G.n1400 G.t3609 132.208
R664 G.n1312 G.t749 132.208
R665 G.n1224 G.t604 132.208
R666 G.n1136 G.t2244 132.208
R667 G.n1048 G.t2106 132.208
R668 G.n963 G.t3762 132.208
R669 G.n881 G.t3617 132.208
R670 G.n805 G.t756 132.208
R671 G.n732 G.t611 132.208
R672 G.n662 G.t2248 132.208
R673 G.n595 G.t1402 132.208
R674 G.n531 G.t109 132.208
R675 G.n470 G.t2907 132.208
R676 G.n412 G.t1617 132.208
R677 G.n357 G.t4410 132.208
R678 G.n308 G.t3120 132.208
R679 G.n262 G.t1407 132.208
R680 G.n219 G.t124 132.208
R681 G.n3777 G.t2917 132.208
R682 G.n3779 G.t1624 132.208
R683 G.n3781 G.t4421 132.208
R684 G.n3783 G.t1598 132.208
R685 G.n3785 G.t1418 132.208
R686 G.n3787 G.t3105 132.208
R687 G.n3789 G.t2924 132.208
R688 G.n3791 G.t105 132.208
R689 G.n3793 G.t4430 132.208
R690 G.n3795 G.t3289 132.208
R691 G.n3797 G.t1570 132.208
R692 G.n3834 G.t410 132.208
R693 G.n3832 G.t2084 132.208
R694 G.n3830 G.t3257 132.208
R695 G.n3828 G.t3453 132.208
R696 G.n3826 G.t1746 132.208
R697 G.n3824 G.t1943 132.208
R698 G.n3822 G.t247 132.208
R699 G.n3820 G.t443 132.208
R700 G.n3818 G.t3249 132.208
R701 G.n3816 G.t466 132.208
R702 G.n3814 G.t1739 132.208
R703 G.n3812 G.t3469 132.208
R704 G.n259 G.t238 132.208
R705 G.n305 G.t1954 132.208
R706 G.n354 G.t3238 132.208
R707 G.n409 G.t457 132.208
R708 G.n467 G.t1724 132.208
R709 G.n528 G.t3458 132.208
R710 G.n592 G.t228 132.208
R711 G.n659 G.t1061 132.208
R712 G.n729 G.t3884 132.208
R713 G.n802 G.t4067 132.208
R714 G.n878 G.t2370 132.208
R715 G.n960 G.t2550 132.208
R716 G.n1045 G.t868 132.208
R717 G.n1133 G.t1050 132.208
R718 G.n1221 G.t3875 132.208
R719 G.n1309 G.t4057 132.208
R720 G.n1397 G.t2365 132.208
R721 G.n1485 G.t4081 132.208
R722 G.n1572 G.t864 132.208
R723 G.n1655 G.t2570 132.208
R724 G.n1733 G.t3868 132.208
R725 G.n1805 G.t1070 132.208
R726 G.n1873 G.t2354 132.208
R727 G.n1935 G.t4076 132.208
R728 G.n1992 G.t857 132.208
R729 G.n2043 G.t2082 132.208
R730 G.n2088 G.t3395 132.208
R731 G.n2459 G.t579 132.208
R732 G.n2461 G.t3420 132.208
R733 G.n2463 G.t3581 132.208
R734 G.n2465 G.t1909 132.208
R735 G.n2467 G.t2072 132.208
R736 G.n2469 G.t403 132.208
R737 G.n2471 G.t571 132.208
R738 G.n2496 G.t204 132.208
R739 G.n2494 G.t6 132.208
R740 G.n2492 G.t1702 132.208
R741 G.n2490 G.t1515 132.208
R742 G.n2488 G.t3214 132.208
R743 G.n2486 G.t3020 132.208
R744 G.n2484 G.t212 132.208
R745 G.n2482 G.t3000 132.208
R746 G.n2040 G.t1716 132.208
R747 G.n1989 G.t550 132.208
R748 G.n1932 G.t3726 132.208
R749 G.n1870 G.t2053 132.208
R750 G.n1802 G.t719 132.208
R751 G.n1730 G.t3566 132.208
R752 G.n1652 G.t2220 132.208
R753 G.n1569 G.t558 132.208
R754 G.n1482 G.t3731 132.208
R755 G.n1394 G.t2062 132.208
R756 G.n1306 G.t3713 132.208
R757 G.n1218 G.t3569 132.208
R758 G.n1130 G.t710 132.208
R759 G.n1042 G.t564 132.208
R760 G.n957 G.t2208 132.208
R761 G.n875 G.t2068 132.208
R762 G.n799 G.t3720 132.208
R763 G.n726 G.t3576 132.208
R764 G.n656 G.t712 132.208
R765 G.n589 G.t4367 132.208
R766 G.n525 G.t3058 132.208
R767 G.n464 G.t1352 132.208
R768 G.n406 G.t56 132.208
R769 G.n351 G.t2867 132.208
R770 G.n302 G.t1563 132.208
R771 G.n3850 G.t4373 132.208
R772 G.n3852 G.t3070 132.208
R773 G.n3854 G.t1366 132.208
R774 G.n3856 G.t65 132.208
R775 G.n3858 G.t2878 132.208
R776 G.n3860 G.t40 132.208
R777 G.n3862 G.t4379 132.208
R778 G.n3864 G.t1550 132.208
R779 G.n3866 G.t1373 132.208
R780 G.n3868 G.t3050 132.208
R781 G.n3870 G.t2883 132.208
R782 G.n3872 G.t1721 132.208
R783 G.n3874 G.t10 132.208
R784 G.n3917 G.t3363 132.208
R785 G.n3915 G.t546 132.208
R786 G.n3913 G.t1692 132.208
R787 G.n3911 G.t1895 132.208
R788 G.n3909 G.t194 132.208
R789 G.n3907 G.t392 132.208
R790 G.n3905 G.t3194 132.208
R791 G.n3903 G.t3396 132.208
R792 G.n3901 G.t1684 132.208
R793 G.n3899 G.t3421 132.208
R794 G.n3897 G.t184 132.208
R795 G.n3895 G.t1910 132.208
R796 G.n3893 G.t3184 132.208
R797 G.n3891 G.t404 132.208
R798 G.n348 G.t1674 132.208
R799 G.n403 G.t3411 132.208
R800 G.n461 G.t167 132.208
R801 G.n522 G.t1900 132.208
R802 G.n586 G.t3174 132.208
R803 G.n653 G.t4015 132.208
R804 G.n723 G.t2321 132.208
R805 G.n796 G.t2500 132.208
R806 G.n872 G.t826 132.208
R807 G.n954 G.t995 132.208
R808 G.n1039 G.t3825 132.208
R809 G.n1127 G.t4011 132.208
R810 G.n1215 G.t2316 132.208
R811 G.n1303 G.t2497 132.208
R812 G.n1391 G.t821 132.208
R813 G.n1479 G.t2516 132.208
R814 G.n1566 G.t3816 132.208
R815 G.n1649 G.t1014 132.208
R816 G.n1727 G.t2303 132.208
R817 G.n1799 G.t4022 132.208
R818 G.n1867 G.t812 132.208
R819 G.n1929 G.t2511 132.208
R820 G.n1986 G.t3809 132.208
R821 G.n2037 G.t541 132.208
R822 G.n2509 G.t1834 132.208
R823 G.n2511 G.t3546 132.208
R824 G.n2513 G.t1861 132.208
R825 G.n2515 G.t2031 132.208
R826 G.n2517 G.t359 132.208
R827 G.n2519 G.t532 132.208
R828 G.n2521 G.t3358 132.208
R829 G.n2523 G.t3537 132.208
R830 G.n2551 G.t3154 132.208
R831 G.n2549 G.t2960 132.208
R832 G.n2547 G.t148 132.208
R833 G.n2545 G.t4470 132.208
R834 G.n2543 G.t1651 132.208
R835 G.n2541 G.t1464 132.208
R836 G.n2539 G.t3159 132.208
R837 G.n2537 G.t1445 132.208
R838 G.n2535 G.t157 132.208
R839 G.n1983 G.t3513 132.208
R840 G.n1926 G.t2179 132.208
R841 G.n1864 G.t510 132.208
R842 G.n1796 G.t3684 132.208
R843 G.n1724 G.t2011 132.208
R844 G.n1646 G.t679 132.208
R845 G.n1563 G.t3522 132.208
R846 G.n1476 G.t2185 132.208
R847 G.n1388 G.t519 132.208
R848 G.n1300 G.t2166 132.208
R849 G.n1212 G.t2018 132.208
R850 G.n1124 G.t3677 132.208
R851 G.n1036 G.t3529 132.208
R852 G.n951 G.t670 132.208
R853 G.n869 G.t526 132.208
R854 G.n793 G.t2172 132.208
R855 G.n720 G.t2025 132.208
R856 G.n650 G.t3679 132.208
R857 G.n583 G.t2817 132.208
R858 G.n519 G.t1505 132.208
R859 G.n458 G.t4319 132.208
R860 G.n400 G.t3011 132.208
R861 G.n3935 G.t1320 132.208
R862 G.n3937 G.t5 132.208
R863 G.n3939 G.t2823 132.208
R864 G.n3941 G.t1516 132.208
R865 G.n3943 G.t4329 132.208
R866 G.n3945 G.t3018 132.208
R867 G.n3947 G.t1327 132.208
R868 G.n3949 G.t2999 132.208
R869 G.n3951 G.t2829 132.208
R870 G.n3953 G.t4504 132.208
R871 G.n3955 G.t4338 132.208
R872 G.n3957 G.t1498 132.208
R873 G.n3959 G.t1331 132.208
R874 G.n3961 G.t162 132.208
R875 G.n3963 G.t2964 132.208
R876 G.n4009 G.t1798 132.208
R877 G.n4007 G.t3506 132.208
R878 G.n4005 G.t137 132.208
R879 G.n4003 G.t341 132.208
R880 G.n4001 G.t3142 132.208
R881 G.n3999 G.t3344 132.208
R882 G.n3997 G.t1626 132.208
R883 G.n3995 G.t1832 132.208
R884 G.n3993 G.t128 132.208
R885 G.n3991 G.t1859 132.208
R886 G.n3989 G.t3131 132.208
R887 G.n3987 G.t356 132.208
R888 G.n3985 G.t1620 132.208
R889 G.n3983 G.t3355 132.208
R890 G.n3981 G.t116 132.208
R891 G.n397 G.t1848 132.208
R892 G.n455 G.t3114 132.208
R893 G.n516 G.t347 132.208
R894 G.n580 G.t1610 132.208
R895 G.n647 G.t2451 132.208
R896 G.n717 G.t785 132.208
R897 G.n790 G.t950 132.208
R898 G.n866 G.t3788 132.208
R899 G.n948 G.t3950 132.208
R900 G.n1033 G.t2269 132.208
R901 G.n1121 G.t2443 132.208
R902 G.n1209 G.t775 132.208
R903 G.n1297 G.t942 132.208
R904 G.n1385 G.t3782 132.208
R905 G.n1473 G.t965 132.208
R906 G.n1560 G.t2260 132.208
R907 G.n1643 G.t3966 132.208
R908 G.n1721 G.t766 132.208
R909 G.n1793 G.t2456 132.208
R910 G.n1861 G.t3773 132.208
R911 G.n1923 G.t959 132.208
R912 G.n1980 G.t2252 132.208
R913 G.n2565 G.t3503 132.208
R914 G.n2567 G.t276 132.208
R915 G.n2569 G.t1992 132.208
R916 G.n2571 G.t302 132.208
R917 G.n2573 G.t487 132.208
R918 G.n2575 G.t3309 132.208
R919 G.n2577 G.t3489 132.208
R920 G.n2579 G.t1791 132.208
R921 G.n2581 G.t1982 132.208
R922 G.n2612 G.t1591 132.208
R923 G.n2610 G.t1409 132.208
R924 G.n2608 G.t3093 132.208
R925 G.n2606 G.t2919 132.208
R926 G.n2604 G.t94 132.208
R927 G.n2602 G.t4425 132.208
R928 G.n2600 G.t1601 132.208
R929 G.n2598 G.t4405 132.208
R930 G.n2596 G.t3106 132.208
R931 G.n2594 G.t1951 132.208
R932 G.n1920 G.t641 132.208
R933 G.n1858 G.t3466 132.208
R934 G.n1790 G.t2138 132.208
R935 G.n1718 G.t463 132.208
R936 G.n1640 G.t3647 132.208
R937 G.n1557 G.t1962 132.208
R938 G.n1470 G.t645 132.208
R939 G.n1382 G.t3476 132.208
R940 G.n1294 G.t626 132.208
R941 G.n1206 G.t472 132.208
R942 G.n1118 G.t2128 132.208
R943 G.n1030 G.t1973 132.208
R944 G.n945 G.t3637 132.208
R945 G.n863 G.t3483 132.208
R946 G.n787 G.t632 132.208
R947 G.n714 G.t483 132.208
R948 G.n644 G.t2133 132.208
R949 G.n577 G.t1270 132.208
R950 G.n513 G.t4459 132.208
R951 G.n452 G.t2766 132.208
R952 G.n4028 G.t1456 132.208
R953 G.n4030 G.t4280 132.208
R954 G.n4032 G.t2959 132.208
R955 G.n4034 G.t1275 132.208
R956 G.n4036 G.t4469 132.208
R957 G.n4038 G.t2777 132.208
R958 G.n4040 G.t1463 132.208
R959 G.n4042 G.t4288 132.208
R960 G.n4044 G.t1444 132.208
R961 G.n4046 G.t1280 132.208
R962 G.n4048 G.t2947 132.208
R963 G.n4050 G.t2782 132.208
R964 G.n4052 G.t4451 132.208
R965 G.n4054 G.t4293 132.208
R966 G.n4056 G.t3110 132.208
R967 G.n4058 G.t1411 132.208
R968 G.n4110 G.t300 132.208
R969 G.n4108 G.t1639 132.208
R970 G.n4106 G.t2264 132.208
R971 G.n4104 G.t784 132.208
R972 G.n4102 G.t1786 132.208
R973 G.n4100 G.t301 132.208
R974 G.n4098 G.t1257 132.208
R975 G.n4096 G.t4273 132.208
R976 G.n4094 G.t746 132.208
R977 G.n4092 G.t3273 132.208
R978 G.n4090 G.t252 132.208
R979 G.n4088 G.t2737 132.208
R980 G.n4086 G.t4234 132.208
R981 G.n4084 G.t2229 132.208
R982 G.n4082 G.t3725 132.208
R983 G.n4080 G.t1726 132.208
R984 G.n4078 G.t3223 132.208
R985 G.n510 G.t1212 132.208
R986 G.n574 G.t2698 132.208
R987 G.n641 G.t1577 132.208
R988 G.n711 G.t2557 132.208
R989 G.n784 G.t1076 132.208
R990 G.n860 G.t2077 132.208
R991 G.n942 G.t590 132.208
R992 G.n1027 G.t1529 132.208
R993 G.n1115 G.t34 132.208
R994 G.n1203 G.t1026 132.208
R995 G.n1291 G.t4046 132.208
R996 G.n1379 G.t552 132.208
R997 G.n1467 G.t3010 132.208
R998 G.n1554 G.t4500 132.208
R999 G.n1637 G.t2507 132.208
R1000 G.n1715 G.t3999 132.208
R1001 G.n1787 G.t2038 132.208
R1002 G.n1855 G.t3532 132.208
R1003 G.n2626 G.t1474 132.208
R1004 G.n2628 G.t2963 132.208
R1005 G.n2630 G.t2898 132.208
R1006 G.n2632 G.t4389 132.208
R1007 G.n2634 G.t2378 132.208
R1008 G.n2636 G.t3417 132.208
R1009 G.n2638 G.t1919 132.208
R1010 G.n2640 G.t2862 132.208
R1011 G.n2642 G.t1361 132.208
R1012 G.n2644 G.t2341 132.208
R1013 G.n2646 G.t855 132.208
R1014 G.n2680 G.t551 132.208
R1015 G.n2678 G.t2042 132.208
R1016 G.n2676 G.t1025 132.208
R1017 G.n2674 G.t2512 132.208
R1018 G.n2672 G.t1528 132.208
R1019 G.n2670 G.t3017 132.208
R1020 G.n2668 G.t2076 132.208
R1021 G.n2666 G.t4055 132.208
R1022 G.n2664 G.t2559 132.208
R1023 G.n2662 G.t2635 132.208
R1024 G.n2660 G.t1149 132.208
R1025 G.n1852 G.t3146 132.208
R1026 G.n1784 G.t1655 132.208
R1027 G.n1712 G.t3673 132.208
R1028 G.n1634 G.t2175 132.208
R1029 G.n1551 G.t4173 132.208
R1030 G.n1464 G.t2675 132.208
R1031 G.n1376 G.t175 132.208
R1032 G.n1288 G.t3707 132.208
R1033 G.n1200 G.t694 132.208
R1034 G.n1112 G.t4213 132.208
R1035 G.n1024 G.t1194 132.208
R1036 G.n939 G.t227 132.208
R1037 G.n857 G.t1711 132.208
R1038 G.n781 G.t723 132.208
R1039 G.n708 G.t2213 132.208
R1040 G.n638 G.t1234 132.208
R1041 G.n571 G.t2335 132.208
R1042 G.n4131 G.t854 132.208
R1043 G.n4133 G.t2856 132.208
R1044 G.n4135 G.t1358 132.208
R1045 G.n4137 G.t3412 132.208
R1046 G.n4139 G.t1918 132.208
R1047 G.n4141 G.t3877 132.208
R1048 G.n4143 G.t2377 132.208
R1049 G.n4145 G.t4386 132.208
R1050 G.n4147 G.t2895 132.208
R1051 G.n4149 G.t439 132.208
R1052 G.n4151 G.t3920 132.208
R1053 G.n4153 G.t902 132.208
R1054 G.n4155 G.t4424 132.208
R1055 G.n4157 G.t1403 132.208
R1056 G.n4159 G.t482 132.208
R1057 G.n4161 G.t1967 132.208
R1058 G.n4163 G.t1289 132.208
R1059 G.n4165 G.t4423 132.208
R1060 G.n4223 G.t3251 132.208
R1061 G.n4221 G.t79 132.208
R1062 G.n4219 G.t728 132.208
R1063 G.n4217 G.t3744 132.208
R1064 G.n4215 G.t234 132.208
R1065 G.n4213 G.t3252 132.208
R1066 G.n4211 G.t4220 132.208
R1067 G.n4209 G.t2719 132.208
R1068 G.n4207 G.t3711 132.208
R1069 G.n4205 G.t1706 132.208
R1070 G.n4203 G.t3203 132.208
R1071 G.n4201 G.t1193 132.208
R1072 G.n4199 G.t2680 132.208
R1073 G.n4197 G.t693 132.208
R1074 G.n4195 G.t2178 132.208
R1075 G.n4193 G.t174 132.208
R1076 G.n4191 G.t1658 132.208
R1077 G.n4189 G.t4167 132.208
R1078 G.n4187 G.t1154 132.208
R1079 G.n635 G.t15 132.208
R1080 G.n705 G.t1002 132.208
R1081 G.n778 G.t4027 132.208
R1082 G.n854 G.t536 132.208
R1083 G.n936 G.t3557 132.208
R1084 G.n1021 G.t4482 132.208
R1085 G.n1109 G.t2989 132.208
R1086 G.n1197 G.t3976 132.208
R1087 G.n1285 G.t2483 132.208
R1088 G.n1373 G.t3516 132.208
R1089 G.n1461 G.t1455 132.208
R1090 G.n1548 G.t2946 132.208
R1091 G.n1631 G.t954 132.208
R1092 G.n1709 G.t2435 132.208
R1093 G.n1781 G.t494 132.208
R1094 G.n2695 G.t1976 132.208
R1095 G.n2697 G.t4434 132.208
R1096 G.n2699 G.t1410 132.208
R1097 G.n2701 G.t1344 132.208
R1098 G.n2703 G.t2839 132.208
R1099 G.n2705 G.t834 132.208
R1100 G.n2707 G.t1858 132.208
R1101 G.n2709 G.t368 132.208
R1102 G.n2711 G.t1312 132.208
R1103 G.n2713 G.t4325 132.208
R1104 G.n2715 G.t799 132.208
R1105 G.n2717 G.t3811 132.208
R1106 G.n2754 G.t3706 132.208
R1107 G.n2752 G.t697 132.208
R1108 G.n2750 G.t4217 132.208
R1109 G.n2748 G.t1198 132.208
R1110 G.n2746 G.t229 132.208
R1111 G.n2744 G.t1710 132.208
R1112 G.n2742 G.t725 132.208
R1113 G.n2740 G.t2722 132.208
R1114 G.n2738 G.t1233 132.208
R1115 G.n2736 G.t1303 132.208
R1116 G.n2734 G.t4316 132.208
R1117 G.n2732 G.t1847 132.208
R1118 G.n1778 G.t364 132.208
R1119 G.n1706 G.t2313 132.208
R1120 G.n1628 G.t830 132.208
R1121 G.n1545 G.t2834 132.208
R1122 G.n1458 G.t1339 132.208
R1123 G.n1370 G.t3387 132.208
R1124 G.n1282 G.t2358 132.208
R1125 G.n1194 G.t3858 132.208
R1126 G.n1106 G.t2876 132.208
R1127 G.n1018 G.t4369 132.208
R1128 G.n933 G.t3435 132.208
R1129 G.n851 G.t414 132.208
R1130 G.n775 G.t3901 132.208
R1131 G.n702 G.t879 132.208
R1132 G.n4246 G.t4404 132.208
R1133 G.n4248 G.t1018 132.208
R1134 G.n4250 G.t4045 132.208
R1135 G.n4252 G.t1527 132.208
R1136 G.n4254 G.t32 132.208
R1137 G.n4256 G.t2074 132.208
R1138 G.n4258 G.t589 132.208
R1139 G.n4260 G.t2552 132.208
R1140 G.n4262 G.t1075 132.208
R1141 G.n4264 G.t3052 132.208
R1142 G.n4266 G.t1576 132.208
R1143 G.n4268 G.t3606 132.208
R1144 G.n4270 G.t2598 132.208
R1145 G.n4272 G.t4098 132.208
R1146 G.n4274 G.t3104 132.208
R1147 G.n4276 G.t84 132.208
R1148 G.n4278 G.t3645 132.208
R1149 G.n4280 G.t627 132.208
R1150 G.n4282 G.t4462 132.208
R1151 G.n4284 G.t3103 132.208
R1152 G.n4348 G.t1686 132.208
R1153 G.n4346 G.t3032 132.208
R1154 G.n4344 G.t3692 132.208
R1155 G.n4342 G.t2195 132.208
R1156 G.n4340 G.t3180 132.208
R1157 G.n4338 G.t1687 132.208
R1158 G.n4336 G.t2665 132.208
R1159 G.n4334 G.t1175 132.208
R1160 G.n4332 G.t2164 132.208
R1161 G.n4330 G.t150 132.208
R1162 G.n4328 G.t1635 132.208
R1163 G.n4326 G.t4148 132.208
R1164 G.n4324 G.t1133 132.208
R1165 G.n4322 G.t3657 132.208
R1166 G.n4320 G.t637 132.208
R1167 G.n4318 G.t3122 132.208
R1168 G.n4316 G.t102 132.208
R1169 G.n4314 G.t2617 132.208
R1170 G.n4312 G.t4111 132.208
R1171 G.n4310 G.t2972 132.208
R1172 G.n4308 G.t3957 132.208
R1173 G.n772 G.t2463 132.208
R1174 G.n848 G.t3497 132.208
R1175 G.n930 G.t2003 132.208
R1176 G.n1015 G.t2929 132.208
R1177 G.n1103 G.t1436 132.208
R1178 G.n1191 G.t2417 132.208
R1179 G.n1279 G.t937 132.208
R1180 G.n1367 G.t1955 132.208
R1181 G.n1455 G.t4414 132.208
R1182 G.n1542 G.t1397 132.208
R1183 G.n1625 G.t3912 132.208
R1184 G.n1703 G.t892 132.208
R1185 G.n2770 G.t3447 132.208
R1186 G.n2772 G.t426 132.208
R1187 G.n2774 G.t2887 132.208
R1188 G.n2776 G.t4375 132.208
R1189 G.n2778 G.t4308 132.208
R1190 G.n2780 G.t1288 132.208
R1191 G.n2782 G.t3794 132.208
R1192 G.n2784 G.t299 132.208
R1193 G.n2786 G.t3318 132.208
R1194 G.n2788 G.t4272 132.208
R1195 G.n2790 G.t2771 132.208
R1196 G.n2792 G.t3761 132.208
R1197 G.n2794 G.t2254 132.208
R1198 G.n2836 G.t2159 132.208
R1199 G.n2834 G.t3659 132.208
R1200 G.n2832 G.t2660 132.208
R1201 G.n2830 G.t4152 132.208
R1202 G.n2828 G.t3175 132.208
R1203 G.n2826 G.t154 132.208
R1204 G.n2824 G.t3688 132.208
R1205 G.n2822 G.t1177 132.208
R1206 G.n2820 G.t4194 132.208
R1207 G.n2818 G.t4263 132.208
R1208 G.n2816 G.t2765 132.208
R1209 G.n2814 G.t289 132.208
R1210 G.n2812 G.t3313 132.208
R1211 G.n1700 G.t773 132.208
R1212 G.n1622 G.t3791 132.208
R1213 G.n1539 G.t1282 132.208
R1214 G.n1452 G.t4301 132.208
R1215 G.n1364 G.t1825 132.208
R1216 G.n1276 G.t815 132.208
R1217 G.n1188 G.t2296 132.208
R1218 G.n1100 G.t1326 132.208
R1219 G.n1012 G.t2816 132.208
R1220 G.n927 G.t1875 132.208
R1221 G.n845 G.t3367 132.208
R1222 G.n4373 G.t2339 132.208
R1223 G.n4375 G.t3834 132.208
R1224 G.n4377 G.t2859 132.208
R1225 G.n4379 G.t3974 132.208
R1226 G.n4381 G.t2478 132.208
R1227 G.n4383 G.t4479 132.208
R1228 G.n4385 G.t2988 132.208
R1229 G.n4387 G.t533 132.208
R1230 G.n4389 G.t3556 132.208
R1231 G.n4391 G.t996 132.208
R1232 G.n4393 G.t4026 132.208
R1233 G.n4395 G.t1501 132.208
R1234 G.n4397 G.t14 132.208
R1235 G.n4399 G.t2061 132.208
R1236 G.n4401 G.t1048 132.208
R1237 G.n4403 G.t2534 132.208
R1238 G.n4405 G.t1551 132.208
R1239 G.n4407 G.t3035 132.208
R1240 G.n4409 G.t2097 132.208
R1241 G.n4411 G.t3590 132.208
R1242 G.n4413 G.t2912 132.208
R1243 G.n4415 G.t1549 132.208
R1244 G.n4485 G.t132 132.208
R1245 G.n4483 G.t1479 132.208
R1246 G.n4481 G.t2147 132.208
R1247 G.n4479 G.t658 132.208
R1248 G.n4477 G.t1618 132.208
R1249 G.n4475 G.t133 132.208
R1250 G.n4473 G.t1118 132.208
R1251 G.n4471 G.t4135 132.208
R1252 G.n4469 G.t622 132.208
R1253 G.n4467 G.t3099 132.208
R1254 G.n4465 G.t74 132.208
R1255 G.n4463 G.t2591 132.208
R1256 G.n4461 G.t4090 132.208
R1257 G.n4459 G.t2105 132.208
R1258 G.n4457 G.t3599 132.208
R1259 G.n4455 G.t1565 132.208
R1260 G.n4453 G.t3047 132.208
R1261 G.n4451 G.t1067 132.208
R1262 G.n4449 G.t2546 132.208
R1263 G.n4447 G.t1420 132.208
R1264 G.n4445 G.t2395 132.208
R1265 G.n4443 G.t917 132.208
R1266 G.n4441 G.t1939 132.208
R1267 G.n924 G.t452 132.208
R1268 G.n1009 G.t1378 132.208
R1269 G.n1097 G.t4398 132.208
R1270 G.n1185 G.t870 132.208
R1271 G.n1273 G.t3896 132.208
R1272 G.n1361 G.t405 132.208
R1273 G.n1449 G.t2871 132.208
R1274 G.n1536 G.t4361 132.208
R1275 G.n1619 G.t2353 132.208
R1276 G.n2853 G.t3847 132.208
R1277 G.n2855 G.t1888 132.208
R1278 G.n2857 G.t3378 132.208
R1279 G.n2859 G.t1334 132.208
R1280 G.n2861 G.t2826 132.208
R1281 G.n2863 G.t2757 132.208
R1282 G.n2865 G.t4251 132.208
R1283 G.n2867 G.t2240 132.208
R1284 G.n2869 G.t3248 132.208
R1285 G.n2871 G.t1751 132.208
R1286 G.n2873 G.t2718 132.208
R1287 G.n2875 G.t1226 132.208
R1288 G.n2877 G.t2207 132.208
R1289 G.n2879 G.t718 132.208
R1290 G.n2925 G.t620 132.208
R1291 G.n2923 G.t2108 132.208
R1292 G.n2921 G.t1113 132.208
R1293 G.n2919 G.t2595 132.208
R1294 G.n2917 G.t1614 132.208
R1295 G.n2915 G.t3102 132.208
R1296 G.n2913 G.t2144 132.208
R1297 G.n2911 G.t4136 132.208
R1298 G.n2909 G.t2642 132.208
R1299 G.n2907 G.t2709 132.208
R1300 G.n2905 G.t1220 132.208
R1301 G.n2903 G.t3237 132.208
R1302 G.n2901 G.t1745 132.208
R1303 G.n2899 G.t3735 132.208
R1304 G.n2897 G.t2235 132.208
R1305 G.n1533 G.t4245 132.208
R1306 G.n1446 G.t2750 132.208
R1307 G.n1358 G.t269 132.208
R1308 G.n1270 G.t3779 132.208
R1309 G.n1182 G.t758 132.208
R1310 G.n1094 G.t4286 132.208
R1311 G.n1006 G.t1269 132.208
R1312 G.n921 G.t316 132.208
R1313 G.n4511 G.t1806 132.208
R1314 G.n4513 G.t796 132.208
R1315 G.n4515 G.t2279 132.208
R1316 G.n4517 G.t1307 132.208
R1317 G.n4519 G.t2412 132.208
R1318 G.n4521 G.t932 132.208
R1319 G.n4523 G.t2926 132.208
R1320 G.n4525 G.t1435 132.208
R1321 G.n4527 G.t3493 132.208
R1322 G.n4529 G.t2002 132.208
R1323 G.n4531 G.t3949 132.208
R1324 G.n4533 G.t2462 132.208
R1325 G.n4535 G.t4458 132.208
R1326 G.n4537 G.t2968 132.208
R1327 G.n4539 G.t518 132.208
R1328 G.n4541 G.t4004 132.208
R1329 G.n4543 G.t979 132.208
R1330 G.n4545 G.t4507 132.208
R1331 G.n4547 G.t1483 132.208
R1332 G.n4549 G.t554 132.208
R1333 G.n4551 G.t2043 132.208
R1334 G.n4553 G.t1357 132.208
R1335 G.n4555 G.t4506 132.208
R1336 G.n4628 G.t3076 132.208
R1337 G.n4626 G.t4440 132.208
R1338 G.n4624 G.t605 132.208
R1339 G.n4622 G.t3621 132.208
R1340 G.n4620 G.t58 132.208
R1341 G.n4618 G.t3077 132.208
R1342 G.n4616 G.t4074 132.208
R1343 G.n4614 G.t2573 132.208
R1344 G.n4612 G.t3586 132.208
R1345 G.n4610 G.t1545 132.208
R1346 G.n4608 G.t3028 132.208
R1347 G.n4606 G.t1045 132.208
R1348 G.n4604 G.t2525 132.208
R1349 G.n4602 G.t563 132.208
R1350 G.n4600 G.t2055 132.208
R1351 G.n4598 G.t4 132.208
R1352 G.n4596 G.t1494 132.208
R1353 G.n4594 G.t4019 132.208
R1354 G.n4592 G.t988 132.208
R1355 G.n4590 G.t4382 132.208
R1356 G.n4588 G.t853 132.208
R1357 G.n4586 G.t3874 132.208
R1358 G.n4584 G.t388 132.208
R1359 G.n4582 G.t3406 132.208
R1360 G.n1003 G.t4344 132.208
R1361 G.n1091 G.t2850 132.208
R1362 G.n1179 G.t3826 132.208
R1363 G.n1267 G.t2330 132.208
R1364 G.n1355 G.t3359 132.208
R1365 G.n1443 G.t1323 132.208
R1366 G.n1530 G.t2808 132.208
R1367 G.n2943 G.t810 132.208
R1368 G.n2945 G.t2287 132.208
R1369 G.n2947 G.t333 132.208
R1370 G.n2949 G.t1818 132.208
R1371 G.n2951 G.t4295 132.208
R1372 G.n2953 G.t1278 132.208
R1373 G.n2955 G.t1214 132.208
R1374 G.n2957 G.t2697 132.208
R1375 G.n2959 G.t706 132.208
R1376 G.n2961 G.t1682 132.208
R1377 G.n2963 G.t200 132.208
R1378 G.n2965 G.t1172 132.208
R1379 G.n2967 G.t4188 132.208
R1380 G.n2969 G.t669 132.208
R1381 G.n2971 G.t3683 132.208
R1382 G.n3020 G.t3584 132.208
R1383 G.n3018 G.t565 132.208
R1384 G.n3016 G.t4069 132.208
R1385 G.n3014 G.t1047 132.208
R1386 G.n3012 G.t52 132.208
R1387 G.n3010 G.t1548 132.208
R1388 G.n3008 G.t603 132.208
R1389 G.n3006 G.t2575 132.208
R1390 G.n3004 G.t1093 132.208
R1391 G.n3002 G.t1163 132.208
R1392 G.n3000 G.t4182 132.208
R1393 G.n2998 G.t1671 132.208
R1394 G.n2996 G.t192 132.208
R1395 G.n2994 G.t2189 132.208
R1396 G.n2992 G.t703 132.208
R1397 G.n2990 G.t2692 132.208
R1398 G.n1440 G.t1207 132.208
R1399 G.n1352 G.t3217 132.208
R1400 G.n1264 G.t2224 132.208
R1401 G.n1176 G.t3719 132.208
R1402 G.n1088 G.t2732 132.208
R1403 G.n4656 G.t4229 132.208
R1404 G.n4658 G.t3265 132.208
R1405 G.n4660 G.t248 132.208
R1406 G.n4662 G.t3757 132.208
R1407 G.n4664 G.t740 132.208
R1408 G.n4666 G.t4271 132.208
R1409 G.n4668 G.t867 132.208
R1410 G.n4670 G.t3895 132.208
R1411 G.n4672 G.t1375 132.208
R1412 G.n4674 G.t4397 132.208
R1413 G.n4676 G.t1935 132.208
R1414 G.n4678 G.t451 132.208
R1415 G.n4680 G.t2393 132.208
R1416 G.n4682 G.t915 132.208
R1417 G.n4684 G.t2910 132.208
R1418 G.n4686 G.t1417 132.208
R1419 G.n4688 G.t3475 132.208
R1420 G.n4690 G.t2440 132.208
R1421 G.n4692 G.t3938 132.208
R1422 G.n4694 G.t2950 132.208
R1423 G.n4696 G.t4441 132.208
R1424 G.n4698 G.t3518 132.208
R1425 G.n4700 G.t503 132.208
R1426 G.n4702 G.t4324 132.208
R1427 G.n4704 G.t2949 132.208
R1428 G.n4782 G.t1522 132.208
R1429 G.n4780 G.t2892 132.208
R1430 G.n4778 G.t3571 132.208
R1431 G.n4776 G.t2073 132.208
R1432 G.n4774 G.t3015 132.208
R1433 G.n4772 G.t1523 132.208
R1434 G.n4770 G.t2508 132.208
R1435 G.n4768 G.t1017 132.208
R1436 G.n4766 G.t2037 132.208
R1437 G.n4764 G.t4499 132.208
R1438 G.n4762 G.t1473 132.208
R1439 G.n4760 G.t3998 132.208
R1440 G.n4758 G.t972 132.208
R1441 G.n4756 G.t3531 132.208
R1442 G.n4754 G.t514 132.208
R1443 G.n4752 G.t2958 132.208
R1444 G.n4750 G.t4450 132.208
R1445 G.n4748 G.t2454 132.208
R1446 G.n4746 G.t3944 132.208
R1447 G.n4744 G.t2833 132.208
R1448 G.n4742 G.t3807 132.208
R1449 G.n4740 G.t2312 132.208
R1450 G.n4738 G.t3339 132.208
R1451 G.n4736 G.t1846 132.208
R1452 G.n4734 G.t2788 132.208
R1453 G.n4732 G.t1299 132.208
R1454 G.n6138 G.t2273 132.208
R1455 G.n6192 G.t790 132.208
R1456 G.n6246 G.t1797 132.208
R1457 G.n6300 G.t4284 132.208
R1458 G.n3038 G.t1262 132.208
R1459 G.n3040 G.t3772 132.208
R1460 G.n3042 G.t750 132.208
R1461 G.n3044 G.t3283 132.208
R1462 G.n3046 G.t259 132.208
R1463 G.n3048 G.t2742 132.208
R1464 G.n3050 G.t4239 132.208
R1465 G.n3052 G.t4172 132.208
R1466 G.n3054 G.t1153 132.208
R1467 G.n3056 G.t3672 132.208
R1468 G.n3058 G.t127 132.208
R1469 G.n3060 G.t3148 132.208
R1470 G.n3062 G.t4132 132.208
R1471 G.n3064 G.t2638 132.208
R1472 G.n3066 G.t3636 132.208
R1473 G.n3068 G.t2137 132.208
R1474 G.n3113 G.t2034 132.208
R1475 G.n3111 G.t3533 132.208
R1476 G.n3109 G.t2502 132.208
R1477 G.n3107 G.t4000 132.208
R1478 G.n3105 G.t3008 132.208
R1479 G.n3103 G.t4503 132.208
R1480 G.n3101 G.t3568 132.208
R1481 G.n3099 G.t1022 132.208
R1482 G.n3097 G.t4048 132.208
R1483 G.n3095 G.t4123 132.208
R1484 G.n3093 G.t2628 132.208
R1485 G.n3091 G.t122 132.208
R1486 G.n3089 G.t3139 132.208
R1487 G.n3087 G.t651 132.208
R1488 G.n3085 G.t3669 132.208
R1489 G.n6356 G.t1146 132.208
R1490 G.n6303 G.t4163 132.208
R1491 G.n6249 G.t1650 132.208
R1492 G.n6195 G.t683 132.208
R1493 G.n6141 G.t2171 132.208
R1494 G.n6087 G.t1187 132.208
R1495 G.n6035 G.t2674 132.208
R1496 G.n4808 G.t1699 132.208
R1497 G.n4810 G.t3197 132.208
R1498 G.n4812 G.t2206 132.208
R1499 G.n4814 G.t3703 132.208
R1500 G.n4816 G.t2717 132.208
R1501 G.n4818 G.t3821 132.208
R1502 G.n4820 G.t2329 132.208
R1503 G.n4822 G.t4340 132.208
R1504 G.n4824 G.t2849 132.208
R1505 G.n4826 G.t385 132.208
R1506 G.n4828 G.t3405 132.208
R1507 G.n4830 G.t851 132.208
R1508 G.n4832 G.t3871 132.208
R1509 G.n4834 G.t1355 132.208
R1510 G.n4836 G.t4381 132.208
R1511 G.n4838 G.t1915 132.208
R1512 G.n4840 G.t895 132.208
R1513 G.n4842 G.t2375 132.208
R1514 G.n4844 G.t1400 132.208
R1515 G.n4846 G.t2894 132.208
R1516 G.n4848 G.t1957 132.208
R1517 G.n4850 G.t3456 132.208
R1518 G.n4852 G.t2770 132.208
R1519 G.n4854 G.t1399 132.208
R1520 G.n4923 G.t222 132.208
R1521 G.n4921 G.t1564 132.208
R1522 G.n4919 G.t2210 132.208
R1523 G.n4917 G.t722 132.208
R1524 G.n4915 G.t1705 132.208
R1525 G.n4913 G.t223 132.208
R1526 G.n4911 G.t1192 132.208
R1527 G.n4909 G.t4209 132.208
R1528 G.n4907 G.t689 132.208
R1529 G.n4905 G.t3196 132.208
R1530 G.n4903 G.t169 132.208
R1531 G.n4901 G.t2672 132.208
R1532 G.n4899 G.t4166 132.208
R1533 G.n4897 G.t2170 132.208
R1534 G.n4895 G.t3668 132.208
R1535 G.n4893 G.t1649 132.208
R1536 G.n4891 G.t3144 132.208
R1537 G.n4889 G.t1145 132.208
R1538 G.n4887 G.t2633 132.208
R1539 G.n4885 G.t1499 132.208
R1540 G.n4883 G.t2481 132.208
R1541 G.n4881 G.t992 132.208
R1542 G.n4879 G.t2017 132.208
R1543 G.n5985 G.t529 132.208
R1544 G.n6034 G.t1454 132.208
R1545 G.n6085 G.t4475 132.208
R1546 G.n6137 G.t949 132.208
R1547 G.n6191 G.t3970 132.208
R1548 G.n6245 G.t492 132.208
R1549 G.n6299 G.t2940 132.208
R1550 G.n6353 G.t4432 132.208
R1551 G.n6406 G.t2428 132.208
R1552 G.n3130 G.t3930 132.208
R1553 G.n3132 G.t1970 132.208
R1554 G.n3134 G.t3461 132.208
R1555 G.n3136 G.t1406 132.208
R1556 G.n3138 G.t2903 132.208
R1557 G.n3140 G.t2836 132.208
R1558 G.n3142 G.t4323 132.208
R1559 G.n3144 G.t2311 132.208
R1560 G.n3146 G.t3343 132.208
R1561 G.n3148 G.t1845 132.208
R1562 G.n3150 G.t2792 132.208
R1563 G.n3152 G.t1302 132.208
R1564 G.n3154 G.t2272 132.208
R1565 G.n3156 G.t794 132.208
R1566 G.n3196 G.t491 132.208
R1567 G.n3194 G.t1977 132.208
R1568 G.n3192 G.t948 132.208
R1569 G.n3190 G.t2438 132.208
R1570 G.n3188 G.t1453 132.208
R1571 G.n3186 G.t2945 132.208
R1572 G.n3184 G.t2016 132.208
R1573 G.n3182 G.t3973 132.208
R1574 G.n3180 G.t2480 132.208
R1575 G.n3178 G.t2565 132.208
R1576 G.n3176 G.t1080 132.208
R1577 G.n3174 G.t3067 132.208
R1578 G.n3172 G.t1583 132.208
R1579 G.n6460 G.t3614 132.208
R1580 G.n6412 G.t2119 132.208
R1581 G.n6361 G.t4105 132.208
R1582 G.n6308 G.t2608 132.208
R1583 G.n6254 G.t93 132.208
R1584 G.n6200 G.t3652 132.208
R1585 G.n6146 G.t633 132.208
R1586 G.n6092 G.t4145 132.208
R1587 G.n6040 G.t1128 132.208
R1588 G.n5989 G.t146 132.208
R1589 G.n5940 G.t1630 132.208
R1590 G.n5894 G.t668 132.208
R1591 G.n4946 G.t2156 132.208
R1592 G.n4948 G.t1170 132.208
R1593 G.n4950 G.t2266 132.208
R1594 G.n4952 G.t789 132.208
R1595 G.n4954 G.t2785 132.208
R1596 G.n4956 G.t1298 132.208
R1597 G.n4958 G.t3336 132.208
R1598 G.n4960 G.t1843 132.208
R1599 G.n4962 G.t3805 132.208
R1600 G.n4964 G.t2310 132.208
R1601 G.n4966 G.t4318 132.208
R1602 G.n4968 G.t2832 132.208
R1603 G.n4970 G.t363 132.208
R1604 G.n4972 G.t3851 132.208
R1605 G.n4974 G.t833 132.208
R1606 G.n4976 G.t4365 132.208
R1607 G.n4978 G.t1341 132.208
R1608 G.n4980 G.t408 132.208
R1609 G.n4982 G.t1897 132.208
R1610 G.n4984 G.t1225 132.208
R1611 G.n4986 G.t4364 132.208
R1612 G.n5046 G.t3169 132.208
R1613 G.n5044 G.t7 132.208
R1614 G.n5042 G.t671 132.208
R1615 G.n5040 G.t3686 132.208
R1616 G.n5038 G.t149 132.208
R1617 G.n5036 G.t3170 132.208
R1618 G.n5034 G.t4147 132.208
R1619 G.n5032 G.t2656 132.208
R1620 G.n5030 G.t3653 132.208
R1621 G.n5028 G.t1629 132.208
R1622 G.n5026 G.t3118 132.208
R1623 G.n5024 G.t1125 132.208
R1624 G.n5022 G.t2612 132.208
R1625 G.n5020 G.t631 132.208
R1626 G.n5018 G.t2122 132.208
R1627 G.n5016 G.t92 132.208
R1628 G.n5014 G.t1582 132.208
R1629 G.n5012 G.t4104 132.208
R1630 G.n5010 G.t1085 132.208
R1631 G.n5008 G.t4453 132.208
R1632 G.n5850 G.t935 132.208
R1633 G.n5893 G.t3947 132.208
R1634 G.n5938 G.t471 132.208
R1635 G.n5984 G.t3486 132.208
R1636 G.n6033 G.t4413 132.208
R1637 G.n6084 G.t2923 132.208
R1638 G.n6136 G.t3907 132.208
R1639 G.n6190 G.t2408 132.208
R1640 G.n6244 G.t3446 132.208
R1641 G.n6298 G.t1391 132.208
R1642 G.n6352 G.t2885 132.208
R1643 G.n6405 G.t886 132.208
R1644 G.n6456 G.t2369 132.208
R1645 G.n6504 G.t419 132.208
R1646 G.n3211 G.t1906 132.208
R1647 G.n3213 G.t4372 132.208
R1648 G.n3215 G.t1348 132.208
R1649 G.n3217 G.t1283 132.208
R1650 G.n3219 G.t2769 132.208
R1651 G.n3221 G.t774 132.208
R1652 G.n3223 G.t1775 132.208
R1653 G.n3225 G.t288 132.208
R1654 G.n3227 G.t1246 132.208
R1655 G.n3229 G.t4262 132.208
R1656 G.n3231 G.t737 132.208
R1657 G.n3233 G.t3752 132.208
R1658 G.n3268 G.t3445 132.208
R1659 G.n3266 G.t427 132.208
R1660 G.n3264 G.t3911 132.208
R1661 G.n3262 G.t891 132.208
R1662 G.n3260 G.t4412 132.208
R1663 G.n3258 G.t1396 132.208
R1664 G.n3256 G.t470 132.208
R1665 G.n3254 G.t2416 132.208
R1666 G.n3252 G.t934 132.208
R1667 G.n3250 G.t1010 132.208
R1668 G.n3248 G.t4032 132.208
R1669 G.n6550 G.t1512 132.208
R1670 G.n6509 G.t23 132.208
R1671 G.n6465 G.t2067 132.208
R1672 G.n6417 G.t578 132.208
R1673 G.n6366 G.t2541 132.208
R1674 G.n6313 G.t1059 132.208
R1675 G.n6259 G.t3044 132.208
R1676 G.n6205 G.t2101 132.208
R1677 G.n6151 G.t3598 132.208
R1678 G.n6097 G.t2586 132.208
R1679 G.n6045 G.t4087 132.208
R1680 G.n5994 G.t3090 132.208
R1681 G.n5945 G.t70 132.208
R1682 G.n5899 G.t3634 132.208
R1683 G.n5854 G.t615 132.208
R1684 G.n5811 G.t4128 132.208
R1685 G.n5771 G.t732 132.208
R1686 G.n5066 G.t3749 132.208
R1687 G.n5068 G.t1240 132.208
R1688 G.n5070 G.t4259 132.208
R1689 G.n5072 G.t1769 132.208
R1690 G.n5074 G.t287 132.208
R1691 G.n5076 G.t2250 132.208
R1692 G.n5078 G.t772 132.208
R1693 G.n5080 G.t2764 132.208
R1694 G.n5082 G.t1281 132.208
R1695 G.n5084 G.t3316 132.208
R1696 G.n5086 G.t2290 132.208
R1697 G.n5088 G.t3793 132.208
R1698 G.n5090 G.t2812 132.208
R1699 G.n5092 G.t4304 132.208
R1700 G.n5094 G.t3365 132.208
R1701 G.n5096 G.t342 132.208
R1702 G.n5098 G.t4187 132.208
R1703 G.n5100 G.t2811 132.208
R1704 G.n5151 G.t1608 132.208
R1705 G.n5149 G.t2961 132.208
R1706 G.n5147 G.t3639 132.208
R1707 G.n5145 G.t2143 132.208
R1708 G.n5143 G.t3094 132.208
R1709 G.n5141 G.t1609 132.208
R1710 G.n5139 G.t2590 132.208
R1711 G.n5137 G.t1108 132.208
R1712 G.n5135 G.t2103 132.208
R1713 G.n5133 G.t69 132.208
R1714 G.n5131 G.t1560 132.208
R1715 G.n5129 G.t4086 132.208
R1716 G.n5127 G.t1063 132.208
R1717 G.n5125 G.t3595 132.208
R1718 G.n5123 G.t580 132.208
R1719 G.n5121 G.t3042 132.208
R1720 G.n5119 G.t27 132.208
R1721 G.n5733 G.t2540 132.208
R1722 G.n5770 G.t4035 132.208
R1723 G.n5809 G.t2906 132.208
R1724 G.n5849 G.t3893 132.208
R1725 G.n5892 G.t2388 132.208
R1726 G.n5937 G.t3426 132.208
R1727 G.n5983 G.t1933 132.208
R1728 G.n6032 G.t2870 132.208
R1729 G.n6083 G.t1370 132.208
R1730 G.n6135 G.t2352 132.208
R1731 G.n6189 G.t865 132.208
R1732 G.n6243 G.t1885 132.208
R1733 G.n6297 G.t4358 132.208
R1734 G.n6351 G.t1333 132.208
R1735 G.n6404 G.t3842 132.208
R1736 G.n6455 G.t825 132.208
R1737 G.n6503 G.t3375 132.208
R1738 G.n6547 G.t355 132.208
R1739 G.n6588 G.t2821 132.208
R1740 G.n3282 G.t4312 132.208
R1741 G.n3284 G.t4244 132.208
R1742 G.n3286 G.t1223 132.208
R1743 G.n3288 G.t3737 132.208
R1744 G.n3290 G.t218 132.208
R1745 G.n3292 G.t3240 132.208
R1746 G.n3294 G.t4207 132.208
R1747 G.n3296 G.t2708 132.208
R1748 G.n3298 G.t3700 132.208
R1749 G.n3300 G.t2201 132.208
R1750 G.n3330 G.t1887 132.208
R1751 G.n3328 G.t3377 132.208
R1752 G.n3326 G.t2351 132.208
R1753 G.n3324 G.t3846 132.208
R1754 G.n3322 G.t2869 132.208
R1755 G.n3320 G.t4360 132.208
R1756 G.n3318 G.t3425 132.208
R1757 G.n3316 G.t869 132.208
R1758 G.n3314 G.t3892 132.208
R1759 G.n3312 G.t3963 132.208
R1760 G.n6592 G.t2469 132.208
R1761 G.n6555 G.t4466 132.208
R1762 G.n6514 G.t2977 132.208
R1763 G.n6470 G.t522 132.208
R1764 G.n6422 G.t3545 132.208
R1765 G.n6371 G.t983 132.208
R1766 G.n6318 G.t4013 132.208
R1767 G.n6264 G.t1493 132.208
R1768 G.n6210 G.t559 132.208
R1769 G.n6156 G.t2050 132.208
R1770 G.n6102 G.t1036 132.208
R1771 G.n6050 G.t2519 132.208
R1772 G.n5999 G.t1540 132.208
R1773 G.n5950 G.t3024 132.208
R1774 G.n5904 G.t2086 132.208
R1775 G.n5859 G.t3583 132.208
R1776 G.n5816 G.t2567 132.208
R1777 G.n5776 G.t3695 132.208
R1778 G.n5737 G.t2198 132.208
R1779 G.n5700 G.t4200 132.208
R1780 G.n5168 G.t2707 132.208
R1781 G.n5170 G.t213 132.208
R1782 G.n5172 G.t3236 132.208
R1783 G.n5174 G.t713 132.208
R1784 G.n5176 G.t3734 132.208
R1785 G.n5178 G.t1222 132.208
R1786 G.n5180 G.t4241 132.208
R1787 G.n5182 G.t1749 132.208
R1788 G.n5184 G.t753 132.208
R1789 G.n5186 G.t2237 132.208
R1790 G.n5188 G.t1267 132.208
R1791 G.n5190 G.t2752 132.208
R1792 G.n5192 G.t1801 132.208
R1793 G.n5194 G.t3290 132.208
R1794 G.n5196 G.t2634 132.208
R1795 G.n5198 G.t1266 132.208
R1796 G.n5240 G.t2460 132.208
R1797 G.n5238 G.t3822 132.208
R1798 G.n5236 G.t4454 132.208
R1799 G.n5234 G.t2966 132.208
R1800 G.n5232 G.t3948 132.208
R1801 G.n5230 G.t2461 132.208
R1802 G.n5228 G.t3492 132.208
R1803 G.n5226 G.t2000 132.208
R1804 G.n5224 G.t2925 132.208
R1805 G.n5222 G.t931 132.208
R1806 G.n5220 G.t2411 132.208
R1807 G.n5218 G.t468 132.208
R1808 G.n5216 G.t1947 132.208
R1809 G.n5214 G.t4409 132.208
R1810 G.n5636 G.t1390 132.208
R1811 G.n5667 G.t3906 132.208
R1812 G.n5698 G.t885 132.208
R1813 G.n5732 G.t3444 132.208
R1814 G.n5769 G.t421 132.208
R1815 G.n5808 G.t3775 132.208
R1816 G.n5848 G.t268 132.208
R1817 G.n5891 G.t3288 132.208
R1818 G.n5936 G.t4243 132.208
R1819 G.n5982 G.t2749 132.208
R1820 G.n6031 G.t3733 132.208
R1821 G.n6082 G.t2233 132.208
R1822 G.n6134 G.t3235 132.208
R1823 G.n6188 G.t1743 132.208
R1824 G.n6242 G.t2706 132.208
R1825 G.n6296 G.t711 132.208
R1826 G.n6350 G.t2200 132.208
R1827 G.n6403 G.t211 132.208
R1828 G.n6454 G.t1693 132.208
R1829 G.n6502 G.t4197 132.208
R1830 G.n6546 G.t1180 132.208
R1831 G.n6587 G.t3693 132.208
R1832 G.n6624 G.t676 132.208
R1833 G.n3341 G.t618 132.208
R1834 G.n3343 G.t2104 132.208
R1835 G.n3345 G.t68 132.208
R1836 G.n3347 G.t1069 132.208
R1837 G.n3349 G.t4085 132.208
R1838 G.n3351 G.t582 132.208
R1839 G.n3353 G.t3597 132.208
R1840 G.n3355 G.t28 132.208
R1841 G.n3357 G.t3043 132.208
R1842 G.n3381 G.t2705 132.208
R1843 G.n3379 G.t4205 132.208
R1844 G.n3377 G.t3234 132.208
R1845 G.n3375 G.t217 132.208
R1846 G.n3373 G.t3732 132.208
R1847 G.n3371 G.t717 132.208
R1848 G.n3369 G.t4242 132.208
R1849 G.n3367 G.t1748 132.208
R1850 G.n6660 G.t267 132.208
R1851 G.n6630 G.t351 132.208
R1852 G.n6597 G.t3372 132.208
R1853 G.n6560 G.t824 132.208
R1854 G.n6519 G.t3839 132.208
R1855 G.n6475 G.t1332 132.208
R1856 G.n6427 G.t4357 132.208
R1857 G.n6376 G.t1884 132.208
R1858 G.n6323 G.t399 132.208
R1859 G.n6269 G.t2348 132.208
R1860 G.n6215 G.t1369 132.208
R1861 G.n6161 G.t2866 132.208
R1862 G.n6107 G.t1929 132.208
R1863 G.n6055 G.t3424 132.208
R1864 G.n6004 G.t2386 132.208
R1865 G.n5955 G.t3891 132.208
R1866 G.n5909 G.t2905 132.208
R1867 G.n5864 G.t4396 132.208
R1868 G.n5821 G.t3472 132.208
R1869 G.n5781 G.t22 132.208
R1870 G.n5742 G.t3041 132.208
R1871 G.n5705 G.t577 132.208
R1872 G.n5671 G.t3594 132.208
R1873 G.n5640 G.t1062 132.208
R1874 G.n5609 G.t4082 132.208
R1875 G.n5254 G.t1559 132.208
R1876 G.n5256 G.t66 132.208
R1877 G.n5258 G.t2102 132.208
R1878 G.n5260 G.t614 132.208
R1879 G.n5262 G.t2589 132.208
R1880 G.n5264 G.t1607 132.208
R1881 G.n5266 G.t3091 132.208
R1882 G.n5268 G.t2142 132.208
R1883 G.n5270 G.t3638 132.208
R1884 G.n5272 G.t2637 132.208
R1885 G.n5274 G.t4134 132.208
R1886 G.n5276 G.t3530 132.208
R1887 G.n5278 G.t2141 132.208
R1888 G.n5311 G.t912 132.208
R1889 G.n5309 G.t2268 132.208
R1890 G.n5307 G.t2908 132.208
R1891 G.n5305 G.t1413 132.208
R1892 G.n5303 G.t2389 132.208
R1893 G.n5301 G.t913 132.208
R1894 G.n5299 G.t1934 132.208
R1895 G.n5297 G.t450 132.208
R1896 G.n5295 G.t1374 132.208
R1897 G.n5293 G.t3890 132.208
R1898 G.n5291 G.t866 132.208
R1899 G.n5557 G.t3423 132.208
R1900 G.n5582 G.t401 132.208
R1901 G.n5607 G.t2865 132.208
R1902 G.n5635 G.t4356 132.208
R1903 G.n5666 G.t2347 132.208
R1904 G.n5697 G.t3841 132.208
R1905 G.n5731 G.t1883 132.208
R1906 G.n5768 G.t3374 132.208
R1907 G.n5807 G.t2222 132.208
R1908 G.n5847 G.t3216 132.208
R1909 G.n5890 G.t1719 132.208
R1910 G.n5935 G.t2691 132.208
R1911 G.n5981 G.t1206 132.208
R1912 G.n6030 G.t2188 132.208
R1913 G.n6081 G.t701 132.208
R1914 G.n6133 G.t1670 132.208
R1915 G.n6187 G.t190 132.208
R1916 G.n6241 G.t1162 132.208
R1917 G.n6295 G.t3678 132.208
R1918 G.n6349 G.t662 132.208
R1919 G.n6402 G.t3158 132.208
R1920 G.n6453 G.t139 132.208
R1921 G.n6501 G.t2646 132.208
R1922 G.n6545 G.t4140 132.208
R1923 G.n6586 G.t2149 132.208
R1924 G.n6623 G.t3643 132.208
R1925 G.n6656 G.t3582 132.208
R1926 G.n6686 G.t562 132.208
R1927 G.n3390 G.t3026 132.208
R1928 G.n3392 G.t4020 132.208
R1929 G.n3394 G.t2518 132.208
R1930 G.n3396 G.t3552 132.208
R1931 G.n3398 G.t2049 132.208
R1932 G.n3400 G.t2984 132.208
R1933 G.n3402 G.t1492 132.208
R1934 G.n3420 G.t1161 132.208
R1935 G.n3418 G.t2652 132.208
R1936 G.n3416 G.t1669 132.208
R1937 G.n3414 G.t3166 132.208
R1938 G.n3412 G.t2187 132.208
R1939 G.n3410 G.t3682 132.208
R1940 G.n6716 G.t2690 132.208
R1941 G.n6692 G.t196 132.208
R1942 G.n6665 G.t3215 132.208
R1943 G.n6635 G.t3304 132.208
R1944 G.n6602 G.t1810 132.208
R1945 G.n6565 G.t3787 132.208
R1946 G.n6524 G.t2285 132.208
R1947 G.n6480 G.t4294 132.208
R1948 G.n6432 G.t2804 132.208
R1949 G.n6381 G.t330 132.208
R1950 G.n6328 G.t3351 132.208
R1951 G.n6274 G.t805 132.208
R1952 G.n6220 G.t4335 132.208
R1953 G.n6166 G.t1319 132.208
R1954 G.n6112 G.t377 132.208
R1955 G.n6060 G.t1867 132.208
R1956 G.n6009 G.t847 132.208
R1957 G.n5960 G.t2328 132.208
R1958 G.n5914 G.t1351 132.208
R1959 G.n5869 G.t2848 132.208
R1960 G.n5826 G.t1912 132.208
R1961 G.n5786 G.t2976 132.208
R1962 G.n5747 G.t1489 132.208
R1963 G.n5710 G.t3548 132.208
R1964 G.n5676 G.t2047 132.208
R1965 G.n5645 G.t4016 132.208
R1966 G.n5614 G.t2517 132.208
R1967 G.n5586 G.t1 132.208
R1968 G.n5561 G.t3023 132.208
R1969 G.n5536 G.t560 132.208
R1970 G.n5323 G.t3579 132.208
R1971 G.n5325 G.t1038 132.208
R1972 G.n5327 G.t49 132.208
R1973 G.n5329 G.t1542 132.208
R1974 G.n5331 G.t601 132.208
R1975 G.n5333 G.t2088 132.208
R1976 G.n5335 G.t1088 132.208
R1977 G.n5337 G.t2572 132.208
R1978 G.n5339 G.t1974 132.208
R1979 G.n5341 G.t600 132.208
R1980 G.n5365 G.t3869 132.208
R1981 G.n5363 G.t734 132.208
R1982 G.n5361 G.t1353 132.208
R1983 G.n5359 G.t4377 132.208
R1984 G.n5357 G.t850 132.208
R1985 G.n5355 G.t3870 132.208
R1986 G.n5353 G.t383 132.208
R1987 G.n5351 G.t3403 132.208
R1988 G.n5497 G.t4339 132.208
R1989 G.n5515 G.t2327 132.208
R1990 G.n5534 G.t3820 132.208
R1991 G.n5556 G.t1864 132.208
R1992 G.n5581 G.t3354 132.208
R1993 G.n5606 G.t1315 132.208
R1994 G.n5634 G.t2806 132.208
R1995 G.n5665 G.t804 132.208
R1996 G.n5696 G.t2284 132.208
R1997 G.n5730 G.t329 132.208
R1998 G.n5767 G.t1814 132.208
R1999 G.n5806 G.t682 132.208
R2000 G.n5846 G.t1648 132.208
R2001 G.n5889 G.t164 132.208
R2002 G.n5934 G.t1144 132.208
R2003 G.n5980 G.t4161 132.208
R2004 G.n6029 G.t650 132.208
R2005 G.n6080 G.t3665 132.208
R2006 G.n6132 G.t113 132.208
R2007 G.n6186 G.t3137 132.208
R2008 G.n6240 G.t4122 132.208
R2009 G.n6294 G.t2131 132.208
R2010 G.n6348 G.t3629 132.208
R2011 G.n6401 G.t1599 132.208
R2012 G.n6452 G.t3085 132.208
R2013 G.n6500 G.t1097 132.208
R2014 G.n6544 G.t2583 132.208
R2015 G.n6585 G.t606 132.208
R2016 G.n6622 G.t2095 132.208
R2017 G.n6655 G.t2032 132.208
R2018 G.n6685 G.t3527 132.208
R2019 G.n6712 G.t1470 132.208
R2020 G.n6736 G.t2455 132.208
R2021 G.n3427 G.t968 132.208
R2022 G.n3429 G.t1997 132.208
R2023 G.n3431 G.t508 132.208
R2024 G.n3433 G.t1434 132.208
R2025 G.n3435 G.t4448 132.208
R2026 G.n3447 G.t4337 132.208
R2027 G.n3445 G.t1318 132.208
R2028 G.n3443 G.t381 132.208
R2029 G.n3441 G.t1866 132.208
R2030 G.n6760 G.t846 132.208
R2031 G.n6742 G.t2333 132.208
R2032 G.n6721 G.t1350 132.208
R2033 G.n6697 G.t3404 132.208
R2034 G.n6670 G.t1914 132.208
R2035 G.n6640 G.t1988 132.208
R2036 G.n6607 G.t506 132.208
R2037 G.n6570 G.t2449 132.208
R2038 G.n6529 G.t964 132.208
R2039 G.n6485 G.t2954 132.208
R2040 G.n6437 G.t1465 132.208
R2041 G.n6386 G.t3524 132.208
R2042 G.n6333 G.t2028 132.208
R2043 G.n6279 G.t3986 132.208
R2044 G.n6225 G.t3004 132.208
R2045 G.n6171 G.t4494 132.208
R2046 G.n6117 G.t3564 132.208
R2047 G.n6065 G.t544 132.208
R2048 G.n6014 G.t4038 132.208
R2049 G.n5965 G.t1015 132.208
R2050 G.n5919 G.t26 132.208
R2051 G.n5874 G.t1518 132.208
R2052 G.n5831 G.t581 132.208
R2053 G.n5791 G.t1668 132.208
R2054 G.n5752 G.t189 132.208
R2055 G.n5715 G.t2186 132.208
R2056 G.n5681 G.t700 132.208
R2057 G.n5650 G.t2688 132.208
R2058 G.n5619 G.t1205 132.208
R2059 G.n5591 G.t3213 132.208
R2060 G.n5566 G.t1718 132.208
R2061 G.n5541 G.t3717 132.208
R2062 G.n5519 G.t2219 132.208
R2063 G.n5500 G.t4228 132.208
R2064 G.n5482 G.t3260 132.208
R2065 G.n5374 G.t244 132.208
R2066 G.n5376 G.t3755 132.208
R2067 G.n5378 G.t735 132.208
R2068 G.n5380 G.t4265 132.208
R2069 G.n5382 G.t1248 132.208
R2070 G.n5384 G.t630 132.208
R2071 G.n5386 G.t3754 132.208
R2072 G.n5400 G.t2304 132.208
R2073 G.n5397 G.t3697 132.208
R2074 G.n5394 G.t4317 132.208
R2075 G.n5391 G.t2828 132.208
R2076 G.n5389 G.t3804 132.208
R2077 G.n5455 G.t2305 132.208
R2078 G.n5467 G.t3335 132.208
R2079 G.n5480 G.t1839 132.208
R2080 G.n5496 G.t2783 132.208
R2081 G.n5514 G.t788 132.208
R2082 G.n5533 G.t2265 132.208
R2083 G.n5555 G.t309 132.208
R2084 G.n5580 G.t1789 132.208
R2085 G.n5605 G.t4277 132.208
R2086 G.n5633 G.t1260 132.208
R2087 G.n5664 G.t3767 132.208
R2088 G.n5695 G.t748 132.208
R2089 G.n5729 G.t3280 132.208
R2090 G.n5766 G.t256 132.208
R2091 G.n5805 G.t3651 132.208
R2092 G.n5845 G.t90 132.208
R2093 G.n5888 G.t3112 132.208
R2094 G.n5933 G.t4103 132.208
R2095 G.n5979 G.t2607 132.208
R2096 G.n6028 G.t3613 132.208
R2097 G.n6079 G.t2116 132.208
R2098 G.n6131 G.t3066 132.208
R2099 G.n6185 G.t1580 132.208
R2100 G.n6239 G.t2560 132.208
R2101 G.n6293 G.t594 132.208
R2102 G.n6347 G.t2080 132.208
R2103 G.n6400 G.t41 132.208
R2104 G.n6451 G.t1534 132.208
R2105 G.n6499 G.t4056 132.208
R2106 G.n6543 G.t1032 132.208
R2107 G.n6584 G.t3572 132.208
R2108 G.n6621 G.t556 132.208
R2109 G.n6654 G.t489 132.208
R2110 G.n6684 G.t1972 132.208
R2111 G.n6711 G.t4431 132.208
R2112 G.n6735 G.t909 132.208
R2113 G.n6756 G.t3929 132.208
R2114 G.n6774 G.t447 132.208
R2115 G.n3452 G.t3460 132.208
R2116 G.n3454 G.t4394 132.208
R2117 G.n3456 G.t2902 132.208
R2118 G.n3463 G.t2781 132.208
R2119 G.n3460 G.t4279 132.208
R2120 G.n6791 G.t3330 132.208
R2121 G.n6773 G.t311 132.208
R2122 G.n6755 G.t3801 132.208
R2123 G.n6734 G.t792 132.208
R2124 G.n6710 G.t4315 132.208
R2125 G.n6683 G.t1841 132.208
R2126 G.n6653 G.t362 132.208
R2127 G.n6620 G.t437 132.208
R2128 G.n6583 G.t3459 132.208
R2129 G.n6542 G.t904 132.208
R2130 G.n6498 G.t3922 132.208
R2131 G.n6450 G.t1404 132.208
R2132 G.n6399 G.t4427 132.208
R2133 G.n6346 G.t1965 132.208
R2134 G.n6292 G.t485 132.208
R2135 G.n6238 G.t2424 132.208
R2136 G.n6184 G.t1447 132.208
R2137 G.n6130 G.t2939 132.208
R2138 G.n6078 G.t2010 132.208
R2139 G.n6027 G.t3508 132.208
R2140 G.n5978 G.t2472 132.208
R2141 G.n5932 G.t3969 132.208
R2142 G.n5887 G.t2983 132.208
R2143 G.n5844 G.t4471 132.208
R2144 G.n5804 G.t3550 132.208
R2145 G.n5765 G.t112 132.208
R2146 G.n5728 G.t3136 132.208
R2147 G.n5694 G.t647 132.208
R2148 G.n5663 G.t3664 132.208
R2149 G.n5632 G.t1141 132.208
R2150 G.n5604 G.t4160 132.208
R2151 G.n5579 G.t1646 132.208
R2152 G.n5554 G.t161 132.208
R2153 G.n5532 G.t2169 132.208
R2154 G.n5513 G.t681 132.208
R2155 G.n5495 G.t2671 132.208
R2156 G.n5479 G.t1695 132.208
R2157 G.n5466 G.t3189 132.208
R2158 G.n5454 G.t2203 132.208
R2159 G.n5444 G.t3701 132.208
R2160 G.n5405 G.t2712 132.208
R2161 G.n5407 G.t4208 132.208
R2162 G.n5410 G.t3596 132.208
R2163 G.n5412 G.t2202 132.208
R2164 G.n6810 G.t1236 132.208
R2165 G.n6805 G.t2728 132.208
R2166 G.n6796 G.t1761 132.208
R2167 G.n6784 G.t3258 132.208
R2168 G.n6769 G.t2247 132.208
R2169 G.n6751 G.t3750 132.208
R2170 G.n6730 G.t2762 132.208
R2171 G.n6706 G.t285 132.208
R2172 G.n6679 G.t3311 132.208
R2173 G.n6649 G.t3391 132.208
R2174 G.n6616 G.t1901 132.208
R2175 G.n6579 G.t3861 132.208
R2176 G.n6538 G.t2363 132.208
R2177 G.n6494 G.t4370 132.208
R2178 G.n6446 G.t2882 132.208
R2179 G.n6395 G.t416 132.208
R2180 G.n6342 G.t3440 132.208
R2181 G.n6288 G.t881 132.208
R2182 G.n6234 G.t4407 132.208
R2183 G.n6180 G.t1389 132.208
R2184 G.n6126 G.t462 132.208
R2185 G.n6074 G.t1946 132.208
R2186 G.n6023 G.t924 132.208
R2187 G.n5974 G.t2407 132.208
R2188 G.n5928 G.t1429 132.208
R2189 G.n5883 G.t2920 132.208
R2190 G.n5840 G.t1993 132.208
R2191 G.n5800 G.t3059 132.208
R2192 G.n5761 G.t1579 132.208
R2193 G.n5724 G.t3610 132.208
R2194 G.n5690 G.t2115 132.208
R2195 G.n5659 G.t4100 132.208
R2196 G.n5628 G.t2606 132.208
R2197 G.n5600 G.t88 132.208
R2198 G.n5575 G.t3111 132.208
R2199 G.n5550 G.t629 132.208
R2200 G.n5528 G.t3650 132.208
R2201 G.n5509 G.t1124 132.208
R2202 G.n5491 G.t140 132.208
R2203 G.n5475 G.t1625 132.208
R2204 G.n5462 G.t664 132.208
R2205 G.n5450 G.t2155 132.208
R2206 G.n5440 G.t1166 132.208
R2207 G.n5433 G.t2654 132.208
R2208 G.n5427 G.t2048 132.208
R2209 G.n5422 G.t663 132.208
R2210 G.n5419 G.t768 132.208
R2211 G.n5417 G.t2152 132.208
R2212 G.n5430 G.t2763 132.208
R2213 G.n5436 G.t1279 132.208
R2214 G.n5443 G.t2249 132.208
R2215 G.n5453 G.t771 132.208
R2216 G.n5465 G.t1767 132.208
R2217 G.n5478 G.t284 132.208
R2218 G.n5494 G.t1238 132.208
R2219 G.n5512 G.t3748 132.208
R2220 G.n5531 G.t730 132.208
R2221 G.n5553 G.t3256 132.208
R2222 G.n5578 G.t236 132.208
R2223 G.n5603 G.t2726 132.208
R2224 G.n5631 G.t4223 132.208
R2225 G.n5662 G.t2214 132.208
R2226 G.n5693 G.t3712 132.208
R2227 G.n5727 G.t1714 132.208
R2228 G.n5764 G.t3206 132.208
R2229 G.n5803 G.t2100 132.208
R2230 G.n5843 G.t3040 132.208
R2231 G.n5886 G.t1557 132.208
R2232 G.n5931 G.t2539 132.208
R2233 G.n5977 G.t1057 132.208
R2234 G.n6026 G.t2066 132.208
R2235 G.n6077 G.t576 132.208
R2236 G.n6129 G.t1511 132.208
R2237 G.n6183 G.t20 132.208
R2238 G.n6237 G.t1009 132.208
R2239 G.n6291 G.t3561 132.208
R2240 G.n6345 G.t539 132.208
R2241 G.n6398 G.t3001 132.208
R2242 G.n6449 G.t4486 132.208
R2243 G.n6497 G.t2492 132.208
R2244 G.n6541 G.t3982 132.208
R2245 G.n6582 G.t2022 132.208
R2246 G.n6619 G.t3520 132.208
R2247 G.n6652 G.t3443 132.208
R2248 G.n6682 G.t424 132.208
R2249 G.n6709 G.t2884 132.208
R2250 G.n6733 G.t3865 132.208
R2251 G.n6754 G.t2368 132.208
R2252 G.n6772 G.t3400 132.208
R2253 G.n6787 G.t1905 132.208
R2254 G.n6799 G.t2845 132.208
R2255 G.n3467 G.t1347 132.208
R2256 G.n3466 G.t2904 120.189
R2257 G.n5416 G.t4336 120.189
R2258 G.n5425 G.t3138 120.189
R2259 G.n5426 G.t1189 120.189
R2260 G.n5429 G.t4478 120.189
R2261 G.n5432 G.t3385 120.189
R2262 G.n5435 G.t2161 120.189
R2263 G.n5439 G.t367 120.189
R2264 G.n5442 G.t3655 120.189
R2265 G.n5449 G.t2835 120.189
R2266 G.n5452 G.t1631 120.189
R2267 G.n5461 G.t4321 120.189
R2268 G.n5464 G.t3121 120.189
R2269 G.n5474 G.t2314 120.189
R2270 G.n5477 G.t1129 120.189
R2271 G.n5490 G.t3806 120.189
R2272 G.n5493 G.t2616 120.189
R2273 G.n5508 G.t1852 120.189
R2274 G.n5511 G.t634 120.189
R2275 G.n5527 G.t3338 120.189
R2276 G.n5530 G.t2123 120.189
R2277 G.n5549 G.t1301 120.189
R2278 G.n5552 G.t95 120.189
R2279 G.n5574 G.t2274 120.189
R2280 G.n5577 G.t1087 120.189
R2281 G.n5599 G.t791 120.189
R2282 G.n5602 G.t4106 120.189
R2283 G.n5627 G.t1799 120.189
R2284 G.n5630 G.t599 120.189
R2285 G.n5658 G.t310 120.189
R2286 G.n5661 G.t3615 120.189
R2287 G.n5689 G.t1263 120.189
R2288 G.n5692 G.t48 120.189
R2289 G.n5723 G.t4283 120.189
R2290 G.n5726 G.t3071 120.189
R2291 G.n5760 G.t752 120.189
R2292 G.n5763 G.t4065 120.189
R2293 G.n5799 G.t3771 120.189
R2294 G.n5802 G.t2564 120.189
R2295 G.n5839 G.t1130 120.189
R2296 G.n5842 G.t4417 120.189
R2297 G.n5882 G.t3656 120.189
R2298 G.n5885 G.t2410 120.189
R2299 G.n5927 G.t635 120.189
R2300 G.n5930 G.t3913 120.189
R2301 G.n5973 G.t3117 120.189
R2302 G.n5976 G.t1949 120.189
R2303 G.n6022 G.t101 120.189
R2304 G.n6025 G.t3449 120.189
R2305 G.n6073 G.t2611 120.189
R2306 G.n6076 G.t1393 120.189
R2307 G.n6125 G.t4107 120.189
R2308 G.n6128 G.t2886 120.189
R2309 G.n6179 G.t2121 120.189
R2310 G.n6182 G.t888 120.189
R2311 G.n6233 G.t3616 120.189
R2312 G.n6236 G.t2371 120.189
R2313 G.n6287 G.t1586 120.189
R2314 G.n6290 G.t423 120.189
R2315 G.n6341 G.t3072 120.189
R2316 G.n6344 G.t1911 120.189
R2317 G.n6394 G.t1086 120.189
R2318 G.n6397 G.t4374 120.189
R2319 G.n6445 G.t2085 120.189
R2320 G.n6448 G.t845 120.189
R2321 G.n6493 G.t596 120.189
R2322 G.n6496 G.t3864 120.189
R2323 G.n6537 G.t1539 120.189
R2324 G.n6540 G.t376 120.189
R2325 G.n6578 G.t45 120.189
R2326 G.n6581 G.t3397 120.189
R2327 G.n6615 G.t1035 120.189
R2328 G.n6618 G.t4334 120.189
R2329 G.n6648 G.t4058 120.189
R2330 G.n6651 G.t2841 120.189
R2331 G.n6678 G.t2439 120.189
R2332 G.n6681 G.t1247 120.189
R2333 G.n6705 G.t955 120.189
R2334 G.n6708 G.t4266 120.189
R2335 G.n6729 G.t1981 120.189
R2336 G.n6732 G.t739 120.189
R2337 G.n6750 G.t4437 120.189
R2338 G.n6753 G.t3263 120.189
R2339 G.n6768 G.t1416 120.189
R2340 G.n6771 G.t246 120.189
R2341 G.n6783 G.t3934 120.189
R2342 G.n6786 G.t2730 120.189
R2343 G.n6795 G.t914 120.189
R2344 G.n6798 G.t4227 120.189
R2345 G.n6804 G.t3471 120.189
R2346 G.n6807 G.t2221 120.189
R2347 G.n6809 G.t449 120.189
R2348 G.n6812 G.t3716 120.189
R2349 G.n5413 G.t188 120.189
R2350 G.n5404 G.t1525 120.189
R2351 G.n5408 G.t3708 120.189
R2352 G.n5437 G.t692 120.189
R2353 G.n5447 G.t3199 120.189
R2354 G.n5459 G.t173 120.189
R2355 G.n5472 G.t2677 120.189
R2356 G.n5488 G.t4171 120.189
R2357 G.n5506 G.t2173 120.189
R2358 G.n5525 G.t3671 120.189
R2359 G.n5547 G.t1652 120.189
R2360 G.n5572 G.t2636 120.189
R2361 G.n5597 G.t1147 120.189
R2362 G.n5625 G.t2140 120.189
R2363 G.n5656 G.t653 120.189
R2364 G.n5687 G.t1606 120.189
R2365 G.n5721 G.t121 120.189
R2366 G.n5758 G.t1107 120.189
R2367 G.n5797 G.t4126 120.189
R2368 G.n5837 G.t1458 120.189
R2369 G.n5880 G.t3971 120.189
R2370 G.n5925 G.t956 120.189
R2371 G.n5971 G.t3511 120.189
R2372 G.n6020 G.t493 120.189
R2373 G.n6071 G.t2942 120.189
R2374 G.n6123 G.t4433 120.189
R2375 G.n6177 G.t2433 120.189
R2376 G.n6231 G.t3933 120.189
R2377 G.n6285 G.t1971 120.189
R2378 G.n6339 G.t3470 120.189
R2379 G.n6392 G.t1408 120.189
R2380 G.n6443 G.t2385 120.189
R2381 G.n6491 G.t907 120.189
R2382 G.n6535 G.t1928 120.189
R2383 G.n6576 G.t444 120.189
R2384 G.n6613 G.t1368 120.189
R2385 G.n6646 G.t4390 120.189
R2386 G.n6676 G.t2793 120.189
R2387 G.n6703 G.t1306 120.189
R2388 G.n6727 G.t2277 120.189
R2389 G.n6748 G.t315 120.189
R2390 G.n6766 G.t1800 120.189
R2391 G.n6781 G.t4285 120.189
R2392 G.n6793 G.t1265 120.189
R2393 G.n6802 G.t3777 120.189
R2394 G.n3461 G.t755 120.189
R2395 G.n3459 G.t3287 120.189
R2396 G.n3450 G.t4452 120.189
R2397 G.n3451 G.t1999 120.189
R2398 G.n6800 G.t515 120.189
R2399 G.n6790 G.t2459 120.189
R2400 G.n6779 G.t973 120.189
R2401 G.n6764 G.t2967 120.189
R2402 G.n6746 G.t1477 120.189
R2403 G.n6725 G.t3535 120.189
R2404 G.n6701 G.t2504 120.189
R2405 G.n6674 G.t4003 120.189
R2406 G.n6644 G.t1102 120.189
R2407 G.n6611 G.t2585 120.189
R2408 G.n6574 G.t1602 120.189
R2409 G.n6533 G.t3087 120.189
R2410 G.n6489 G.t2136 120.189
R2411 G.n6441 G.t3633 120.189
R2412 G.n6390 G.t2632 120.189
R2413 G.n6337 G.t125 120.189
R2414 G.n6283 G.t3145 120.189
R2415 G.n6229 G.t654 120.189
R2416 G.n6175 G.t3670 120.189
R2417 G.n6121 G.t1148 120.189
R2418 G.n6069 G.t4165 120.189
R2419 G.n6018 G.t1653 120.189
R2420 G.n5969 G.t168 120.189
R2421 G.n5923 G.t2177 120.189
R2422 G.n5878 G.t686 120.189
R2423 G.n5835 G.t2678 120.189
R2424 G.n5795 G.t807 120.189
R2425 G.n5756 G.t2289 120.189
R2426 G.n5719 G.t1322 120.189
R2427 G.n5685 G.t2810 120.189
R2428 G.n5654 G.t1869 120.189
R2429 G.n5623 G.t3361 120.189
R2430 G.n5595 G.t2332 120.189
R2431 G.n5570 G.t3828 120.189
R2432 G.n5545 G.t2851 120.189
R2433 G.n5523 G.t387 120.189
R2434 G.n5504 G.t3408 120.189
R2435 G.n5486 G.t852 120.189
R2436 G.n5470 G.t3876 120.189
R2437 G.n5457 G.t1356 120.189
R2438 G.n5445 G.t4383 120.189
R2439 G.n5392 G.t1916 120.189
R2440 G.n5395 G.t435 120.189
R2441 G.n5398 G.t2734 120.189
R2442 G.n5401 G.t1371 120.189
R2443 G.n5368 G.t1742 120.189
R2444 G.n5369 G.t3075 120.189
R2445 G.n5370 G.t743 120.189
R2446 G.n5371 G.t2228 120.189
R2447 G.n5372 G.t250 120.189
R2448 G.n5373 G.t1730 120.189
R2449 G.n5468 G.t4230 120.189
R2450 G.n5484 G.t1213 120.189
R2451 G.n5502 G.t3721 120.189
R2452 G.n5521 G.t704 120.189
R2453 G.n5543 G.t3218 120.189
R2454 G.n5568 G.t4190 120.189
R2455 G.n5593 G.t2693 120.189
R2456 G.n5621 G.t3685 120.189
R2457 G.n5652 G.t2191 120.189
R2458 G.n5683 G.t3168 120.189
R2459 G.n5717 G.t1675 120.189
R2460 G.n5754 G.t2655 120.189
R2461 G.n5793 G.t1167 120.189
R2462 G.n5833 G.t3013 120.189
R2463 G.n5876 G.t1020 120.189
R2464 G.n5921 G.t2505 120.189
R2465 G.n5967 G.t547 120.189
R2466 G.n6016 G.t2036 120.189
R2467 G.n6067 G.t4497 120.189
R2468 G.n6119 G.t1472 120.189
R2469 G.n6173 G.t3991 120.189
R2470 G.n6227 G.t971 120.189
R2471 G.n6281 G.t3526 120.189
R2472 G.n6335 G.t513 120.189
R2473 G.n6388 G.t2957 120.189
R2474 G.n6439 G.t3946 120.189
R2475 G.n6487 G.t2453 120.189
R2476 G.n6531 G.t3485 120.189
R2477 G.n6572 G.t1994 120.189
R2478 G.n6609 G.t2921 120.189
R2479 G.n6642 G.t1428 120.189
R2480 G.n6672 G.t4349 120.189
R2481 G.n6699 G.t2855 120.189
R2482 G.n6723 G.t3829 120.189
R2483 G.n6744 G.t1874 120.189
R2484 G.n6762 G.t3364 120.189
R2485 G.n6777 G.t1325 120.189
R2486 G.n6788 G.t2814 120.189
R2487 G.n3440 G.t813 120.189
R2488 G.n3439 G.t2291 120.189
R2489 G.n3438 G.t339 120.189
R2490 G.n3423 G.t1496 120.189
R2491 G.n3424 G.t3553 120.189
R2492 G.n3425 G.t2056 120.189
R2493 G.n3426 G.t4023 120.189
R2494 G.n6775 G.t2527 120.189
R2495 G.n6759 G.t11 120.189
R2496 G.n6741 G.t3030 120.189
R2497 G.n6720 G.t569 120.189
R2498 G.n6696 G.t4072 120.189
R2499 G.n6669 G.t1049 120.189
R2500 G.n6639 G.t2648 120.189
R2501 G.n6606 G.t4144 120.189
R2502 G.n6569 G.t3162 120.189
R2503 G.n6528 G.t142 120.189
R2504 G.n6484 G.t3680 120.189
R2505 G.n6436 G.t665 120.189
R2506 G.n6385 G.t4184 120.189
R2507 G.n6332 G.t1679 120.189
R2508 G.n6278 G.t195 120.189
R2509 G.n6224 G.t2192 120.189
R2510 G.n6170 G.t705 120.189
R2511 G.n6116 G.t2694 120.189
R2512 G.n6064 G.t1211 120.189
R2513 G.n6013 G.t3219 120.189
R2514 G.n5964 G.t1725 120.189
R2515 G.n5918 G.t3724 120.189
R2516 G.n5873 G.t2226 120.189
R2517 G.n5830 G.t4233 120.189
R2518 G.n5790 G.t2350 120.189
R2519 G.n5751 G.t3849 120.189
R2520 G.n5714 G.t2868 120.189
R2521 G.n5680 G.t4362 120.189
R2522 G.n5649 G.t3428 120.189
R2523 G.n5618 G.t406 120.189
R2524 G.n5590 G.t3897 120.189
R2525 G.n5565 G.t872 120.189
R2526 G.n5540 G.t4400 120.189
R2527 G.n5518 G.t1938 120.189
R2528 G.n5499 G.t454 120.189
R2529 G.n5481 G.t2394 120.189
R2530 G.n5350 G.t919 120.189
R2531 G.n5349 G.t2911 120.189
R2532 G.n5348 G.t1422 120.189
R2533 G.n5347 G.t3477 120.189
R2534 G.n5346 G.t1986 120.189
R2535 G.n5345 G.t4289 120.189
R2536 G.n5344 G.t2922 120.189
R2537 G.n5314 G.t3312 120.189
R2538 G.n5315 G.t131 120.189
R2539 G.n5316 G.t2281 120.189
R2540 G.n5317 G.t3784 120.189
R2541 G.n5318 G.t1805 120.189
R2542 G.n5319 G.t3297 120.189
R2543 G.n5320 G.t1272 120.189
R2544 G.n5321 G.t2755 120.189
R2545 G.n5322 G.t760 120.189
R2546 G.n5516 G.t2238 120.189
R2547 G.n5538 G.t271 120.189
R2548 G.n5563 G.t1227 120.189
R2549 G.n5588 G.t4246 120.189
R2550 G.n5616 G.t720 120.189
R2551 G.n5647 G.t3736 120.189
R2552 G.n5678 G.t220 120.189
R2553 G.n5712 G.t3239 120.189
R2554 G.n5749 G.t4204 120.189
R2555 G.n5788 G.t2713 120.189
R2556 G.n5828 G.t57 120.189
R2557 G.n5871 G.t2574 120.189
R2558 G.n5916 G.t4073 120.189
R2559 G.n5962 G.t2089 120.189
R2560 G.n6011 G.t3585 120.189
R2561 G.n6062 G.t1541 120.189
R2562 G.n6114 G.t3027 120.189
R2563 G.n6168 G.t1041 120.189
R2564 G.n6222 G.t2524 120.189
R2565 G.n6276 G.t561 120.189
R2566 G.n6330 G.t2051 120.189
R2567 G.n6383 G.t3 120.189
R2568 G.n6434 G.t990 120.189
R2569 G.n6482 G.t4018 120.189
R2570 G.n6526 G.t527 120.189
R2571 G.n6567 G.t3547 120.189
R2572 G.n6604 G.t4472 120.189
R2573 G.n6637 G.t2980 120.189
R2574 G.n6667 G.t1381 120.189
R2575 G.n6694 G.t4402 120.189
R2576 G.n6718 G.t876 120.189
R2577 G.n6739 G.t3434 120.189
R2578 G.n6757 G.t411 120.189
R2579 G.n3409 G.t2877 120.189
R2580 G.n3408 G.t4366 120.189
R2581 G.n3407 G.t2355 120.189
R2582 G.n3406 G.t3852 120.189
R2583 G.n3405 G.t1892 120.189
R2584 G.n3384 G.t3048 120.189
R2585 G.n3385 G.t586 120.189
R2586 G.n3386 G.t3602 120.189
R2587 G.n3387 G.t1071 120.189
R2588 G.n3388 G.t4091 120.189
R2589 G.n3389 G.t1571 120.189
R2590 G.n6737 G.t76 120.189
R2591 G.n6715 G.t2110 120.189
R2592 G.n6691 G.t1117 120.189
R2593 G.n6664 G.t2599 120.189
R2594 G.n6634 G.t4199 120.189
R2595 G.n6601 G.t1186 120.189
R2596 G.n6564 G.t214 120.189
R2597 G.n6523 G.t1698 120.189
R2598 G.n6479 G.t714 120.189
R2599 G.n6431 G.t2204 120.189
R2600 G.n6380 G.t1221 120.189
R2601 G.n6327 G.t3245 120.189
R2602 G.n6273 G.t1747 120.189
R2603 G.n6219 G.t3739 120.189
R2604 G.n6165 G.t2236 120.189
R2605 G.n6111 G.t4247 120.189
R2606 G.n6059 G.t2756 120.189
R2607 G.n6008 G.t272 120.189
R2608 G.n5959 G.t3293 120.189
R2609 G.n5913 G.t761 120.189
R2610 G.n5868 G.t3781 120.189
R2611 G.n5825 G.t1273 120.189
R2612 G.n5785 G.t3910 120.189
R2613 G.n5746 G.t894 120.189
R2614 G.n5709 G.t4411 120.189
R2615 G.n5675 G.t1398 120.189
R2616 G.n5644 G.t473 120.189
R2617 G.n5613 G.t1956 120.189
R2618 G.n5585 G.t939 120.189
R2619 G.n5560 G.t2419 120.189
R2620 G.n5535 G.t1439 120.189
R2621 G.n5290 G.t3494 120.189
R2622 G.n5289 G.t2004 120.189
R2623 G.n5288 G.t3956 120.189
R2624 G.n5287 G.t2464 120.189
R2625 G.n5286 G.t4460 120.189
R2626 G.n5285 G.t2973 120.189
R2627 G.n5284 G.t520 120.189
R2628 G.n5283 G.t3541 120.189
R2629 G.n5282 G.t1328 120.189
R2630 G.n5281 G.t4473 120.189
R2631 G.n5243 G.t91 120.189
R2632 G.n5244 G.t1441 120.189
R2633 G.n5245 G.t3641 120.189
R2634 G.n5246 G.t624 120.189
R2635 G.n5247 G.t3100 120.189
R2636 G.n5248 G.t77 120.189
R2637 G.n5249 G.t2596 120.189
R2638 G.n5250 G.t4092 120.189
R2639 G.n5251 G.t2107 120.189
R2640 G.n5252 G.t3604 120.189
R2641 G.n5253 G.t1566 120.189
R2642 G.n5558 G.t2551 120.189
R2643 G.n5583 G.t1068 120.189
R2644 G.n5611 G.t2071 120.189
R2645 G.n5642 G.t584 120.189
R2646 G.n5673 G.t1521 120.189
R2647 G.n5707 G.t30 120.189
R2648 G.n5744 G.t1016 120.189
R2649 G.n5783 G.t4040 120.189
R2650 G.n5823 G.t1382 120.189
R2651 G.n5866 G.t3898 120.189
R2652 G.n5911 G.t877 120.189
R2653 G.n5957 G.t3429 120.189
R2654 G.n6006 G.t407 120.189
R2655 G.n6057 G.t2874 120.189
R2656 G.n6109 G.t4363 120.189
R2657 G.n6163 G.t2356 120.189
R2658 G.n6217 G.t3850 120.189
R2659 G.n6271 G.t1893 120.189
R2660 G.n6325 G.t3382 120.189
R2661 G.n6378 G.t1337 120.189
R2662 G.n6429 G.t2308 120.189
R2663 G.n6477 G.t827 120.189
R2664 G.n6521 G.t1842 120.189
R2665 G.n6562 G.t361 120.189
R2666 G.n6599 G.t1297 120.189
R2667 G.n6632 G.t4313 120.189
R2668 G.n6662 G.t2720 120.189
R2669 G.n6689 G.t1228 120.189
R2670 G.n6713 G.t2209 120.189
R2671 G.n3366 G.t225 120.189
R2672 G.n3365 G.t1703 120.189
R2673 G.n3364 G.t4210 120.189
R2674 G.n3363 G.t1190 120.189
R2675 G.n3362 G.t3702 120.189
R2676 G.n3361 G.t687 120.189
R2677 G.n3360 G.t3195 120.189
R2678 G.n3333 G.t103 120.189
R2679 G.n3334 G.t2127 120.189
R2680 G.n3335 G.t639 120.189
R2681 G.n3336 G.t2621 120.189
R2682 G.n3337 G.t1134 120.189
R2683 G.n3338 G.t3128 120.189
R2684 G.n3339 G.t1638 120.189
R2685 G.n3340 G.t3661 120.189
R2686 G.n6687 G.t2664 120.189
R2687 G.n6659 G.t4154 120.189
R2688 G.n6629 G.t1239 120.189
R2689 G.n6596 G.t2731 120.189
R2690 G.n6559 G.t1768 120.189
R2691 G.n6518 G.t3264 120.189
R2692 G.n6474 G.t2251 120.189
R2693 G.n6426 G.t3756 120.189
R2694 G.n6375 G.t2768 120.189
R2695 G.n6322 G.t291 120.189
R2696 G.n6268 G.t3315 120.189
R2697 G.n6214 G.t778 120.189
R2698 G.n6160 G.t3792 120.189
R2699 G.n6106 G.t1285 120.189
R2700 G.n6054 G.t4303 120.189
R2701 G.n6003 G.t1826 120.189
R2702 G.n5954 G.t346 120.189
R2703 G.n5908 G.t2298 120.189
R2704 G.n5863 G.t819 120.189
R2705 G.n5820 G.t2819 120.189
R2706 G.n5780 G.t953 120.189
R2707 G.n5741 G.t2437 120.189
R2708 G.n5704 G.t1452 120.189
R2709 G.n5670 G.t2948 120.189
R2710 G.n5639 G.t2015 120.189
R2711 G.n5608 G.t3517 120.189
R2712 G.n5213 G.t2485 120.189
R2713 G.n5212 G.t3978 120.189
R2714 G.n5211 G.t2993 120.189
R2715 G.n5210 G.t534 120.189
R2716 G.n5209 G.t3558 120.189
R2717 G.n5208 G.t1000 120.189
R2718 G.n5207 G.t4029 120.189
R2719 G.n5206 G.t1506 120.189
R2720 G.n5205 G.t18 120.189
R2721 G.n5204 G.t2063 120.189
R2722 G.n5203 G.t573 120.189
R2723 G.n5202 G.t2879 120.189
R2724 G.n5201 G.t1519 120.189
R2725 G.n5154 G.t3751 120.189
R2726 G.n5155 G.t621 120.189
R2727 G.n5156 G.t2758 120.189
R2728 G.n5157 G.t4252 120.189
R2729 G.n5158 G.t2239 120.189
R2730 G.n5159 G.t3742 120.189
R2731 G.n5160 G.t1753 120.189
R2732 G.n5161 G.t3246 120.189
R2733 G.n5162 G.t1229 120.189
R2734 G.n5163 G.t2716 120.189
R2735 G.n5164 G.t721 120.189
R2736 G.n5165 G.t1704 120.189
R2737 G.n5166 G.t221 120.189
R2738 G.n5167 G.t1191 120.189
R2739 G.n5637 G.t4206 120.189
R2740 G.n5668 G.t688 120.189
R2741 G.n5702 G.t3699 120.189
R2742 G.n5739 G.t165 120.189
R2743 G.n5778 G.t3190 120.189
R2744 G.n5818 G.t566 120.189
R2745 G.n5861 G.t3031 120.189
R2746 G.n5906 G.t12 120.189
R2747 G.n5952 G.t2528 120.189
R2748 G.n6001 G.t4024 120.189
R2749 G.n6052 G.t2054 120.189
R2750 G.n6104 G.t3554 120.189
R2751 G.n6158 G.t1497 120.189
R2752 G.n6212 G.t2987 120.189
R2753 G.n6266 G.t991 120.189
R2754 G.n6320 G.t2475 120.189
R2755 G.n6373 G.t528 120.189
R2756 G.n6424 G.t1450 120.189
R2757 G.n6472 G.t4474 120.189
R2758 G.n6516 G.t947 120.189
R2759 G.n6557 G.t3965 120.189
R2760 G.n6594 G.t490 120.189
R2761 G.n6627 G.t3505 120.189
R2762 G.n6657 G.t1896 120.189
R2763 G.n3311 G.t412 120.189
R2764 G.n3310 G.t1340 120.189
R2765 G.n3309 G.t3857 120.189
R2766 G.n3308 G.t832 120.189
R2767 G.n3307 G.t3386 120.189
R2768 G.n3306 G.t366 120.189
R2769 G.n3305 G.t2831 120.189
R2770 G.n3304 G.t4322 120.189
R2771 G.n3303 G.t2309 120.189
R2772 G.n3271 G.t3760 120.189
R2773 G.n3272 G.t1249 120.189
R2774 G.n3273 G.t4269 120.189
R2775 G.n3274 G.t1777 120.189
R2776 G.n3275 G.t296 120.189
R2777 G.n3276 G.t2258 120.189
R2778 G.n3277 G.t779 120.189
R2779 G.n3278 G.t2776 120.189
R2780 G.n3279 G.t1827 120.189
R2781 G.n3280 G.t3324 120.189
R2782 G.n6625 G.t425 120.189
R2783 G.n6591 G.t1913 120.189
R2784 G.n6554 G.t889 120.189
R2785 G.n6513 G.t2372 120.189
R2786 G.n6469 G.t1394 120.189
R2787 G.n6421 G.t2891 120.189
R2788 G.n6370 G.t1950 120.189
R2789 G.n6317 G.t3914 120.189
R2790 G.n6263 G.t2415 120.189
R2791 G.n6209 G.t4418 120.189
R2792 G.n6155 G.t2928 120.189
R2793 G.n6101 G.t474 120.189
R2794 G.n6049 G.t3495 120.189
R2795 G.n5998 G.t940 120.189
R2796 G.n5949 G.t3955 120.189
R2797 G.n5903 G.t1442 120.189
R2798 G.n5858 G.t4456 120.189
R2799 G.n5815 G.t2007 120.189
R2800 G.n5775 G.t96 120.189
R2801 G.n5736 G.t1589 120.189
R2802 G.n5699 G.t636 120.189
R2803 G.n5118 G.t2125 120.189
R2804 G.n5117 G.t1131 120.189
R2805 G.n5116 G.t2618 120.189
R2806 G.n5115 G.t1632 120.189
R2807 G.n5114 G.t3129 120.189
R2808 G.n5113 G.t2162 120.189
R2809 G.n5112 G.t4151 120.189
R2810 G.n5111 G.t2659 120.189
R2811 G.n5110 G.t153 120.189
R2812 G.n5109 G.t3179 120.189
R2813 G.n5108 G.t673 120.189
R2814 G.n5107 G.t3690 120.189
R2815 G.n5106 G.t1176 120.189
R2816 G.n5105 G.t4195 120.189
R2817 G.n5104 G.t2059 120.189
R2818 G.n5103 G.t685 120.189
R2819 G.n5049 G.t793 120.189
R2820 G.n5050 G.t2163 120.189
R2821 G.n5051 G.t4307 120.189
R2822 G.n5052 G.t1290 120.189
R2823 G.n5053 G.t3795 120.189
R2824 G.n5054 G.t780 120.189
R2825 G.n5055 G.t3321 120.189
R2826 G.n5056 G.t297 120.189
R2827 G.n5057 G.t2774 120.189
R2828 G.n5058 G.t4270 120.189
R2829 G.n5059 G.t2256 120.189
R2830 G.n5060 G.t3271 120.189
R2831 G.n5061 G.t1774 120.189
R2832 G.n5062 G.t2735 120.189
R2833 G.n5063 G.t1245 120.189
R2834 G.n5064 G.t2225 120.189
R2835 G.n5065 G.t736 120.189
R2836 G.n5734 G.t1723 120.189
R2837 G.n5773 G.t245 120.189
R2838 G.n5813 G.t2111 120.189
R2839 G.n5856 G.t78 120.189
R2840 G.n5901 G.t1572 120.189
R2841 G.n5947 G.t4089 120.189
R2842 G.n5996 G.t1072 120.189
R2843 G.n6047 G.t3603 120.189
R2844 G.n6099 G.t587 120.189
R2845 G.n6153 G.t3049 120.189
R2846 G.n6207 G.t31 120.189
R2847 G.n6261 G.t2547 120.189
R2848 G.n6315 G.t4042 120.189
R2849 G.n6368 G.t2069 120.189
R2850 G.n6419 G.t3007 120.189
R2851 G.n6467 G.t1517 120.189
R2852 G.n6511 G.t2501 120.189
R2853 G.n6552 G.t1012 120.189
R2854 G.n6589 G.t2033 120.189
R2855 G.n3246 G.t545 120.189
R2856 G.n3245 G.t3455 120.189
R2857 G.n3244 G.t1960 120.189
R2858 G.n3243 G.t2893 120.189
R2859 G.n3242 G.t901 120.189
R2860 G.n3241 G.t2376 120.189
R2861 G.n3240 G.t432 120.189
R2862 G.n3239 G.t1917 120.189
R2863 G.n3238 G.t4380 120.189
R2864 G.n3237 G.t1354 120.189
R2865 G.n3236 G.t3873 120.189
R2866 G.n3199 G.t795 120.189
R2867 G.n3200 G.t2794 120.189
R2868 G.n3201 G.t1310 120.189
R2869 G.n3202 G.t3345 120.189
R2870 G.n3203 G.t1856 120.189
R2871 G.n3204 G.t3813 120.189
R2872 G.n3205 G.t2317 120.189
R2873 G.n3206 G.t4330 120.189
R2874 G.n3207 G.t3389 120.189
R2875 G.n3208 G.t373 120.189
R2876 G.n3209 G.t1975 120.189
R2877 G.n3210 G.t3473 120.189
R2878 G.n6549 G.t2434 120.189
R2879 G.n6508 G.t3935 120.189
R2880 G.n6464 G.t2943 120.189
R2881 G.n6416 G.t4438 120.189
R2882 G.n6365 G.t3512 120.189
R2883 G.n6312 G.t957 120.189
R2884 G.n6258 G.t3972 120.189
R2885 G.n6204 G.t1459 120.189
R2886 G.n6150 G.t4481 120.189
R2887 G.n6096 G.t2019 120.189
R2888 G.n6044 G.t535 120.189
R2889 G.n5993 G.t2486 120.189
R2890 G.n5944 G.t1001 120.189
R2891 G.n5898 G.t2997 120.189
R2892 G.n5853 G.t1503 120.189
R2893 G.n5810 G.t3560 120.189
R2894 G.n5007 G.t1654 120.189
R2895 G.n5006 G.t3151 120.189
R2896 G.n5005 G.t2174 120.189
R2897 G.n5004 G.t3675 120.189
R2898 G.n5003 G.t2679 120.189
R2899 G.n5002 G.t4174 120.189
R2900 G.n5001 G.t3200 120.189
R2901 G.n5000 G.t178 120.189
R2902 G.n4999 G.t3709 120.189
R2903 G.n4998 G.t1196 120.189
R2904 G.n4997 G.t4216 120.189
R2905 G.n4996 G.t1709 120.189
R2906 G.n4995 G.t233 120.189
R2907 G.n4994 G.t2212 120.189
R2908 G.n4993 G.t727 120.189
R2909 G.n4992 G.t2723 120.189
R2910 G.n4991 G.t1235 120.189
R2911 G.n4990 G.t3607 120.189
R2912 G.n4989 G.t2223 120.189
R2913 G.n4926 G.t2334 120.189
R2914 G.n4927 G.t3710 120.189
R2915 G.n4928 G.t1345 120.189
R2916 G.n4929 G.t2840 120.189
R2917 G.n4930 G.t836 120.189
R2918 G.n4931 G.t2318 120.189
R2919 G.n4932 G.t371 120.189
R2920 G.n4933 G.t1857 120.189
R2921 G.n4934 G.t4327 120.189
R2922 G.n4935 G.t1311 120.189
R2923 G.n4936 G.t3810 120.189
R2924 G.n4937 G.t323 120.189
R2925 G.n4938 G.t3342 120.189
R2926 G.n4939 G.t4287 120.189
R2927 G.n4940 G.t2791 120.189
R2928 G.n4941 G.t3780 120.189
R2929 G.n4942 G.t2275 120.189
R2930 G.n4943 G.t3291 120.189
R2931 G.n4944 G.t1802 120.189
R2932 G.n4945 G.t3662 120.189
R2933 G.n5851 G.t1634 120.189
R2934 G.n5896 G.t3130 120.189
R2935 G.n5942 G.t1132 120.189
R2936 G.n5991 G.t2622 120.189
R2937 G.n6042 G.t640 120.189
R2938 G.n6094 G.t2126 120.189
R2939 G.n6148 G.t104 120.189
R2940 G.n6202 G.t1590 120.189
R2941 G.n6256 G.t4112 120.189
R2942 G.n6310 G.t1089 120.189
R2943 G.n6363 G.t3618 120.189
R2944 G.n6414 G.t51 120.189
R2945 G.n6462 G.t3073 120.189
R2946 G.n6506 G.t4068 120.189
R2947 G.n3171 G.t2568 120.189
R2948 G.n3170 G.t3580 120.189
R2949 G.n3169 G.t2087 120.189
R2950 G.n3168 G.t502 120.189
R2951 G.n3167 G.t3521 120.189
R2952 G.n3166 G.t4443 120.189
R2953 G.n3165 G.t2441 120.189
R2954 G.n3164 G.t3939 120.189
R2955 G.n3163 G.t1984 120.189
R2956 G.n3162 G.t3474 120.189
R2957 G.n3161 G.t1419 120.189
R2958 G.n3160 G.t2909 120.189
R2959 G.n3159 G.t916 120.189
R2960 G.n3116 G.t2337 120.189
R2961 G.n3117 G.t4350 120.189
R2962 G.n3118 G.t2857 120.189
R2963 G.n3119 G.t393 120.189
R2964 G.n3120 G.t3415 120.189
R2965 G.n3121 G.t860 120.189
R2966 G.n3122 G.t3881 120.189
R2967 G.n3123 G.t1362 120.189
R2968 G.n3124 G.t438 120.189
R2969 G.n3125 G.t1925 120.189
R2970 G.n3126 G.t3528 120.189
R2971 G.n3127 G.t516 120.189
R2972 G.n3128 G.t3997 120.189
R2973 G.n3129 G.t974 120.189
R2974 G.n6459 G.t4498 120.189
R2975 G.n6411 G.t1478 120.189
R2976 G.n6360 G.t548 120.189
R2977 G.n6307 G.t2506 120.189
R2978 G.n6253 G.t1021 120.189
R2979 G.n6199 G.t3014 120.189
R2980 G.n6145 G.t1526 120.189
R2981 G.n6091 G.t3570 120.189
R2982 G.n6039 G.t2075 120.189
R2983 G.n5988 G.t4052 120.189
R2984 G.n5939 G.t2556 120.189
R2985 G.n4878 G.t35 120.189
R2986 G.n4877 G.t3056 120.189
R2987 G.n4876 G.t592 120.189
R2988 G.n4875 G.t3220 120.189
R2989 G.n4874 G.t202 120.189
R2990 G.n4873 G.t3722 120.189
R2991 G.n4872 G.t707 120.189
R2992 G.n4871 G.t4231 120.189
R2993 G.n4870 G.t1215 120.189
R2994 G.n4869 G.t251 120.189
R2995 G.n4868 G.t1733 120.189
R2996 G.n4867 G.t744 120.189
R2997 G.n4866 G.t2736 120.189
R2998 G.n4865 G.t1255 120.189
R2999 G.n4864 G.t3275 120.189
R3000 G.n4863 G.t1781 120.189
R3001 G.n4862 G.t3765 120.189
R3002 G.n4861 G.t2263 120.189
R3003 G.n4860 G.t4275 120.189
R3004 G.n4859 G.t2780 120.189
R3005 G.n4858 G.t642 120.189
R3006 G.n4857 G.t3778 120.189
R3007 G.n4785 G.t3894 120.189
R3008 G.n4786 G.t745 120.189
R3009 G.n4787 G.t2899 120.189
R3010 G.n4788 G.t4387 120.189
R3011 G.n4789 G.t2380 120.189
R3012 G.n4790 G.t3882 120.189
R3013 G.n4791 G.t1922 120.189
R3014 G.n4792 G.t3416 120.189
R3015 G.n4793 G.t1360 120.189
R3016 G.n4794 G.t2861 120.189
R3017 G.n4795 G.t858 120.189
R3018 G.n4796 G.t1876 120.189
R3019 G.n4797 G.t390 120.189
R3020 G.n4798 G.t1329 120.189
R3021 G.n4799 G.t4347 120.189
R3022 G.n4800 G.t818 120.189
R3023 G.n4801 G.t3830 120.189
R3024 G.n4802 G.t343 120.189
R3025 G.n4803 G.t3362 120.189
R3026 G.n4804 G.t698 120.189
R3027 G.n4805 G.t3202 120.189
R3028 G.n4806 G.t182 120.189
R3029 G.n4807 G.t2681 120.189
R3030 G.n5986 G.t4175 120.189
R3031 G.n6037 G.t2181 120.189
R3032 G.n6089 G.t3676 120.189
R3033 G.n6143 G.t1660 120.189
R3034 G.n6197 G.t3152 120.189
R3035 G.n6251 G.t1152 120.189
R3036 G.n6305 G.t2639 120.189
R3037 G.n6358 G.t656 120.189
R3038 G.n6409 G.t1613 120.189
R3039 G.n6457 G.t126 120.189
R3040 G.n3084 G.t1109 120.189
R3041 G.n3083 G.t4129 120.189
R3042 G.n3082 G.t616 120.189
R3043 G.n3081 G.t3635 120.189
R3044 G.n3080 G.t2045 120.189
R3045 G.n3079 G.t553 120.189
R3046 G.n3078 G.t1486 120.189
R3047 G.n3077 G.t4006 120.189
R3048 G.n3076 G.t978 120.189
R3049 G.n3075 G.t3538 120.189
R3050 G.n3074 G.t517 120.189
R3051 G.n3073 G.t2971 120.189
R3052 G.n3072 G.t4457 120.189
R3053 G.n3071 G.t2465 120.189
R3054 G.n3023 G.t3687 120.189
R3055 G.n3024 G.t1174 120.189
R3056 G.n3025 G.t4193 120.189
R3057 G.n3026 G.t1685 120.189
R3058 G.n3027 G.t205 120.189
R3059 G.n3028 G.t2196 120.189
R3060 G.n3029 G.t709 120.189
R3061 G.n3030 G.t2701 120.189
R3062 G.n3031 G.t1737 120.189
R3063 G.n3032 G.t3228 120.189
R3064 G.n3033 G.t340 120.189
R3065 G.n3034 G.t1823 120.189
R3066 G.n3035 G.t814 120.189
R3067 G.n3036 G.t2295 120.189
R3068 G.n3037 G.t1324 120.189
R3069 G.n6407 G.t2815 120.189
R3070 G.n6355 G.t1870 120.189
R3071 G.n6302 G.t3831 120.189
R3072 G.n6248 G.t2338 120.189
R3073 G.n6194 G.t4348 120.189
R3074 G.n6140 G.t2858 120.189
R3075 G.n6086 G.t391 120.189
R3076 G.n4731 G.t3413 120.189
R3077 G.n4730 G.t861 120.189
R3078 G.n4729 G.t3878 120.189
R3079 G.n4728 G.t1363 120.189
R3080 G.n4727 G.t4385 120.189
R3081 G.n4726 G.t1923 120.189
R3082 G.n4725 G.t13 120.189
R3083 G.n4724 G.t1500 120.189
R3084 G.n4723 G.t567 120.189
R3085 G.n4722 G.t2058 120.189
R3086 G.n4721 G.t1046 120.189
R3087 G.n4720 G.t2531 120.189
R3088 G.n4719 G.t1547 120.189
R3089 G.n4718 G.t3034 120.189
R3090 G.n4717 G.t2093 120.189
R3091 G.n4716 G.t4077 120.189
R3092 G.n4715 G.t2578 120.189
R3093 G.n4714 G.t60 120.189
R3094 G.n4713 G.t3081 120.189
R3095 G.n4712 G.t607 120.189
R3096 G.n4711 G.t3624 120.189
R3097 G.n4710 G.t1099 120.189
R3098 G.n4709 G.t4119 120.189
R3099 G.n4708 G.t1989 120.189
R3100 G.n4707 G.t619 120.189
R3101 G.n4631 G.t936 120.189
R3102 G.n4632 G.t2282 120.189
R3103 G.n4633 G.t4446 120.189
R3104 G.n4634 G.t1425 120.189
R3105 G.n4635 G.t3940 120.189
R3106 G.n4636 G.t923 120.189
R3107 G.n4637 G.t3479 120.189
R3108 G.n4638 G.t460 120.189
R3109 G.n4639 G.t2914 120.189
R3110 G.n4640 G.t4406 120.189
R3111 G.n4641 G.t2398 120.189
R3112 G.n4642 G.t3437 120.189
R3113 G.n4643 G.t1941 120.189
R3114 G.n4644 G.t2880 120.189
R3115 G.n4645 G.t1383 120.189
R3116 G.n4646 G.t2362 120.189
R3117 G.n4647 G.t873 120.189
R3118 G.n4648 G.t1898 120.189
R3119 G.n4649 G.t409 120.189
R3120 G.n4650 G.t2231 120.189
R3121 G.n4651 G.t254 120.189
R3122 G.n4652 G.t1734 120.189
R3123 G.n4653 G.t4236 120.189
R3124 G.n4654 G.t1216 120.189
R3125 G.n4655 G.t3727 120.189
R3126 G.n1087 G.t708 120.189
R3127 G.n1175 G.t3226 120.189
R3128 G.n1263 G.t203 120.189
R3129 G.n1351 G.t2696 120.189
R3130 G.n1439 G.t4191 120.189
R3131 G.n1527 G.t2194 120.189
R3132 G.n2989 G.t3171 120.189
R3133 G.n2988 G.t1680 120.189
R3134 G.n2987 G.t2657 120.189
R3135 G.n2986 G.t1171 120.189
R3136 G.n2985 G.t2157 120.189
R3137 G.n2984 G.t666 120.189
R3138 G.n2983 G.t3592 120.189
R3139 G.n2982 G.t2096 120.189
R3140 G.n2981 G.t3036 120.189
R3141 G.n2980 G.t1051 120.189
R3142 G.n2979 G.t2533 120.189
R3143 G.n2978 G.t572 120.189
R3144 G.n2977 G.t2060 120.189
R3145 G.n2976 G.t19 120.189
R3146 G.n2975 G.t1504 120.189
R3147 G.n2974 G.t4025 120.189
R3148 G.n2928 G.t724 120.189
R3149 G.n2929 G.t2721 120.189
R3150 G.n2930 G.t1232 120.189
R3151 G.n2931 G.t3250 120.189
R3152 G.n2932 G.t1758 120.189
R3153 G.n2933 G.t3743 120.189
R3154 G.n2934 G.t2245 120.189
R3155 G.n2935 G.t4256 120.189
R3156 G.n2936 G.t3300 120.189
R3157 G.n2937 G.t280 120.189
R3158 G.n2938 G.t1894 120.189
R3159 G.n2939 G.t3383 120.189
R3160 G.n2940 G.t2357 120.189
R3161 G.n2941 G.t3854 120.189
R3162 G.n2942 G.t2875 120.189
R3163 G.n1614 G.t4368 120.189
R3164 G.n1529 G.t3430 120.189
R3165 G.n1442 G.t878 120.189
R3166 G.n1354 G.t3899 120.189
R3167 G.n1266 G.t1384 120.189
R3168 G.n1178 G.t4403 120.189
R3169 G.n1090 G.t1942 120.189
R3170 G.n1002 G.t458 120.189
R3171 G.n4581 G.t2399 120.189
R3172 G.n4580 G.t922 120.189
R3173 G.n4579 G.t2915 120.189
R3174 G.n4578 G.t1424 120.189
R3175 G.n4577 G.t3481 120.189
R3176 G.n4576 G.t1567 120.189
R3177 G.n4575 G.t3051 120.189
R3178 G.n4574 G.t2112 120.189
R3179 G.n4573 G.t3605 120.189
R3180 G.n4572 G.t2597 120.189
R3181 G.n4571 G.t4095 120.189
R3182 G.n4570 G.t3101 120.189
R3183 G.n4569 G.t82 120.189
R3184 G.n4568 G.t3642 120.189
R3185 G.n4567 G.t1120 120.189
R3186 G.n4566 G.t4138 120.189
R3187 G.n4565 G.t1619 120.189
R3188 G.n4564 G.t136 120.189
R3189 G.n4563 G.t2150 120.189
R3190 G.n4562 G.t660 120.189
R3191 G.n4561 G.t2647 120.189
R3192 G.n4560 G.t1160 120.189
R3193 G.n4559 G.t3542 120.189
R3194 G.n4558 G.t2158 120.189
R3195 G.n4488 G.t2482 120.189
R3196 G.n4489 G.t3836 120.189
R3197 G.n4490 G.t1490 120.189
R3198 G.n4491 G.t2978 120.189
R3199 G.n4492 G.t982 120.189
R3200 G.n4493 G.t2470 120.189
R3201 G.n4494 G.t521 120.189
R3202 G.n4495 G.t2009 120.189
R3203 G.n4496 G.t4463 120.189
R3204 G.n4497 G.t1446 120.189
R3205 G.n4498 G.t3959 120.189
R3206 G.n4499 G.t481 120.189
R3207 G.n4500 G.t3501 120.189
R3208 G.n4501 G.t4422 120.189
R3209 G.n4502 G.t2932 120.189
R3210 G.n4503 G.t3919 120.189
R3211 G.n4504 G.t2420 120.189
R3212 G.n4505 G.t3454 120.189
R3213 G.n4506 G.t1958 120.189
R3214 G.n4507 G.t3785 120.189
R3215 G.n4508 G.t1811 120.189
R3216 G.n4509 G.t3301 120.189
R3217 G.n4510 G.t1274 120.189
R3218 G.n920 G.t2759 120.189
R3219 G.n1005 G.t764 120.189
R3220 G.n1093 G.t2243 120.189
R3221 G.n1181 G.t274 120.189
R3222 G.n1269 G.t1756 120.189
R3223 G.n1357 G.t4250 120.189
R3224 G.n1445 G.t1230 120.189
R3225 G.n1532 G.t3740 120.189
R3226 G.n1616 G.t226 120.189
R3227 G.n2896 G.t3247 120.189
R3228 G.n2895 G.t4212 120.189
R3229 G.n2894 G.t2714 120.189
R3230 G.n2893 G.t3704 120.189
R3231 G.n2892 G.t2205 120.189
R3232 G.n2891 G.t628 120.189
R3233 G.n2890 G.t3644 120.189
R3234 G.n2889 G.t83 120.189
R3235 G.n2888 G.t2601 120.189
R3236 G.n2887 G.t4097 120.189
R3237 G.n2886 G.t2114 120.189
R3238 G.n2885 G.t3608 120.189
R3239 G.n2884 G.t1575 120.189
R3240 G.n2883 G.t3057 120.189
R3241 G.n2882 G.t1074 120.189
R3242 G.n2839 G.t2259 120.189
R3243 G.n2840 G.t4274 120.189
R3244 G.n2841 G.t2779 120.189
R3245 G.n2842 G.t305 120.189
R3246 G.n2843 G.t3326 120.189
R3247 G.n2844 G.t783 120.189
R3248 G.n2845 G.t3799 120.189
R3249 G.n2846 G.t1292 120.189
R3250 G.n2847 G.t352 120.189
R3251 G.n2848 G.t1836 120.189
R3252 G.n2849 G.t3450 120.189
R3253 G.n2850 G.t433 120.189
R3254 G.n2851 G.t3918 120.189
R3255 G.n2852 G.t897 120.189
R3256 G.n1697 G.t4419 120.189
R3257 G.n1618 G.t1401 120.189
R3258 G.n1535 G.t476 120.189
R3259 G.n1448 G.t2422 120.189
R3260 G.n1360 G.t941 120.189
R3261 G.n1272 G.t2934 120.189
R3262 G.n1184 G.t1443 120.189
R3263 G.n1096 G.t3502 120.189
R3264 G.n1008 G.t2008 120.189
R3265 G.n923 G.t3960 120.189
R3266 G.n4440 G.t2468 120.189
R3267 G.n4439 G.t4464 120.189
R3268 G.n4438 G.t2975 120.189
R3269 G.n4437 G.t523 120.189
R3270 G.n4436 G.t3125 120.189
R3271 G.n4435 G.t107 120.189
R3272 G.n4434 G.t3658 120.189
R3273 G.n4433 G.t643 120.189
R3274 G.n4432 G.t4155 120.189
R3275 G.n4431 G.t1137 120.189
R3276 G.n4430 G.t156 120.189
R3277 G.n4429 G.t1641 120.189
R3278 G.n4428 G.t675 120.189
R3279 G.n4427 G.t2667 120.189
R3280 G.n4426 G.t1179 120.189
R3281 G.n4425 G.t3182 120.189
R3282 G.n4424 G.t1690 120.189
R3283 G.n4423 G.t3694 120.189
R3284 G.n4422 G.t2199 120.189
R3285 G.n4421 G.t4198 120.189
R3286 G.n4420 G.t2704 120.189
R3287 G.n4419 G.t574 120.189
R3288 G.n4418 G.t3705 120.189
R3289 G.n4351 G.t4049 120.189
R3290 G.n4352 G.t882 120.189
R3291 G.n4353 G.t3039 120.189
R3292 G.n4354 G.t24 120.189
R3293 G.n4355 G.t2537 120.189
R3294 G.n4356 G.t4036 120.189
R3295 G.n4357 G.t2064 120.189
R3296 G.n4358 G.t3562 120.189
R3297 G.n4359 G.t1508 120.189
R3298 G.n4360 G.t3002 120.189
R3299 G.n4361 G.t1004 120.189
R3300 G.n4362 G.t2024 120.189
R3301 G.n4363 G.t537 120.189
R3302 G.n4364 G.t1462 120.189
R3303 G.n4365 G.t4485 120.189
R3304 G.n4366 G.t962 120.189
R3305 G.n4367 G.t3979 120.189
R3306 G.n4368 G.t501 120.189
R3307 G.n4369 G.t3519 120.189
R3308 G.n4370 G.t823 120.189
R3309 G.n4371 G.t3373 120.189
R3310 G.n4372 G.t353 120.189
R3311 G.n844 G.t2822 120.189
R3312 G.n926 G.t4309 120.189
R3313 G.n1011 G.t2300 120.189
R3314 G.n1099 G.t3797 120.189
R3315 G.n1187 G.t1831 120.189
R3316 G.n1275 G.t3322 120.189
R3317 G.n1363 G.t1287 120.189
R3318 G.n1451 G.t2775 120.189
R3319 G.n1538 G.t781 120.189
R3320 G.n1621 G.t1778 120.189
R3321 G.n1699 G.t298 120.189
R3322 G.n2810 G.t1252 120.189
R3323 G.n2809 G.t4267 120.189
R3324 G.n2808 G.t741 120.189
R3325 G.n2807 G.t3758 120.189
R3326 G.n2806 G.t2168 120.189
R3327 G.n2805 G.t677 120.189
R3328 G.n2804 G.t1642 120.189
R3329 G.n2803 G.t4156 120.189
R3330 G.n2802 G.t1138 120.189
R3331 G.n2801 G.t3663 120.189
R3332 G.n2800 G.t644 120.189
R3333 G.n2799 G.t3135 120.189
R3334 G.n2798 G.t110 120.189
R3335 G.n2797 G.t2625 120.189
R3336 G.n2757 G.t3814 120.189
R3337 G.n2758 G.t1313 120.189
R3338 G.n2759 G.t4331 120.189
R3339 G.n2760 G.t1862 120.189
R3340 G.n2761 G.t375 120.189
R3341 G.n2762 G.t2322 120.189
R3342 G.n2763 G.t840 120.189
R3343 G.n2764 G.t2842 120.189
R3344 G.n2765 G.t1902 120.189
R3345 G.n2766 G.t3401 120.189
R3346 G.n2767 G.t497 120.189
R3347 G.n2768 G.t1985 120.189
R3348 G.n2769 G.t958 120.189
R3349 G.n1775 G.t2442 120.189
R3350 G.n1702 G.t1460 120.189
R3351 G.n1624 G.t2951 120.189
R3352 G.n1541 G.t2020 120.189
R3353 G.n1454 G.t3980 120.189
R3354 G.n1366 G.t2489 120.189
R3355 G.n1278 G.t4487 120.189
R3356 G.n1190 G.t2998 120.189
R3357 G.n1102 G.t540 120.189
R3358 G.n1014 G.t3563 120.189
R3359 G.n929 G.t1005 120.189
R3360 G.n847 G.t4033 120.189
R3361 G.n771 G.t1509 120.189
R3362 G.n4307 G.t21 120.189
R3363 G.n4306 G.t2065 120.189
R3364 G.n4305 G.t179 120.189
R3365 G.n4304 G.t1662 120.189
R3366 G.n4303 G.t696 120.189
R3367 G.n4302 G.t2182 120.189
R3368 G.n4301 G.t1197 120.189
R3369 G.n4300 G.t2684 120.189
R3370 G.n4299 G.t1715 120.189
R3371 G.n4298 G.t3207 120.189
R3372 G.n4297 G.t2215 120.189
R3373 G.n4296 G.t4222 120.189
R3374 G.n4295 G.t2725 120.189
R3375 G.n4294 G.t237 120.189
R3376 G.n4293 G.t3255 120.189
R3377 G.n4292 G.t731 120.189
R3378 G.n4291 G.t3745 120.189
R3379 G.n4290 G.t1237 120.189
R3380 G.n4289 G.t4260 120.189
R3381 G.n4288 G.t2117 120.189
R3382 G.n4287 G.t742 120.189
R3383 G.n4226 G.t1094 120.189
R3384 G.n4227 G.t2425 120.189
R3385 G.n4228 G.t89 120.189
R3386 G.n4229 G.t1584 120.189
R3387 G.n4230 G.t4101 120.189
R3388 G.n4231 G.t1081 120.189
R3389 G.n4232 G.t3611 120.189
R3390 G.n4233 G.t595 120.189
R3391 G.n4234 G.t3061 120.189
R3392 G.n4235 G.t42 120.189
R3393 G.n4236 G.t2558 120.189
R3394 G.n4237 G.t3575 120.189
R3395 G.n4238 G.t2079 120.189
R3396 G.n4239 G.t3021 120.189
R3397 G.n4240 G.t1531 120.189
R3398 G.n4241 G.t2513 120.189
R3399 G.n4242 G.t1028 120.189
R3400 G.n4243 G.t2044 120.189
R3401 G.n4244 G.t555 120.189
R3402 G.n4245 G.t2366 120.189
R3403 G.n701 G.t420 120.189
R3404 G.n774 G.t1903 120.189
R3405 G.n850 G.t4371 120.189
R3406 G.n932 G.t1349 120.189
R3407 G.n1017 G.t3862 120.189
R3408 G.n1105 G.t837 120.189
R3409 G.n1193 G.t3392 120.189
R3410 G.n1281 G.t372 120.189
R3411 G.n1369 G.t2838 120.189
R3412 G.n1457 G.t4328 120.189
R3413 G.n1544 G.t2319 120.189
R3414 G.n1627 G.t3346 120.189
R3415 G.n1705 G.t1854 120.189
R3416 G.n1777 G.t2797 120.189
R3417 G.n1847 G.t1308 120.189
R3418 G.n2731 G.t2278 120.189
R3419 G.n2730 G.t797 120.189
R3420 G.n2729 G.t3714 120.189
R3421 G.n2728 G.t2217 120.189
R3422 G.n2727 G.t3209 120.189
R3423 G.n2726 G.t1201 120.189
R3424 G.n2725 G.t2686 120.189
R3425 G.n2724 G.t699 120.189
R3426 G.n2723 G.t2184 120.189
R3427 G.n2722 G.t185 120.189
R3428 G.n2721 G.t1664 120.189
R3429 G.n2720 G.t4179 120.189
R3430 G.n2683 G.t862 120.189
R3431 G.n2684 G.t2863 120.189
R3432 G.n2685 G.t1367 120.189
R3433 G.n2686 G.t3422 120.189
R3434 G.n2687 G.t1926 120.189
R3435 G.n2688 G.t3885 120.189
R3436 G.n2689 G.t2383 120.189
R3437 G.n2690 G.t4391 120.189
R3438 G.n2691 G.t3462 120.189
R3439 G.n2692 G.t445 120.189
R3440 G.n2693 G.t2039 120.189
R3441 G.n2694 G.t3539 120.189
R3442 G.n1849 G.t2509 120.189
R3443 G.n1780 G.t4007 120.189
R3444 G.n1708 G.t3016 120.189
R3445 G.n1630 G.t4509 120.189
R3446 G.n1547 G.t3573 120.189
R3447 G.n1460 G.t1029 120.189
R3448 G.n1372 G.t4054 120.189
R3449 G.n1284 G.t1532 120.189
R3450 G.n1196 G.t38 120.189
R3451 G.n1108 G.t2081 120.189
R3452 G.n1020 G.t593 120.189
R3453 G.n935 G.t2561 120.189
R3454 G.n853 G.t1082 120.189
R3455 G.n777 G.t3062 120.189
R3456 G.n704 G.t1581 120.189
R3457 G.n634 G.t3612 120.189
R3458 G.n4186 G.t1735 120.189
R3459 G.n4185 G.t3227 120.189
R3460 G.n4184 G.t2230 120.189
R3461 G.n4183 G.t3728 120.189
R3462 G.n4182 G.t2740 120.189
R3463 G.n4181 G.t4238 120.189
R3464 G.n4180 G.t3276 120.189
R3465 G.n4179 G.t257 120.189
R3466 G.n4178 G.t3768 120.189
R3467 G.n4177 G.t1259 120.189
R3468 G.n4176 G.t4278 120.189
R3469 G.n4175 G.t1787 120.189
R3470 G.n4174 G.t307 120.189
R3471 G.n4173 G.t2267 120.189
R3472 G.n4172 G.t786 120.189
R3473 G.n4171 G.t2784 120.189
R3474 G.n4170 G.t1296 120.189
R3475 G.n4169 G.t3666 120.189
R3476 G.n4168 G.t2280 120.189
R3477 G.n4113 G.t2643 120.189
R3478 G.n4114 G.t3987 120.189
R3479 G.n4115 G.t1647 120.189
R3480 G.n4116 G.t3140 120.189
R3481 G.n4117 G.t1142 120.189
R3482 G.n4118 G.t2629 120.189
R3483 G.n4119 G.t648 120.189
R3484 G.n4120 G.t2132 120.189
R3485 G.n4121 G.t114 120.189
R3486 G.n4122 G.t1600 120.189
R3487 G.n4123 G.t4120 120.189
R3488 G.n4124 G.t612 120.189
R3489 G.n4125 G.t3625 120.189
R3490 G.n4126 G.t63 120.189
R3491 G.n4127 G.t3082 120.189
R3492 G.n4128 G.t4078 120.189
R3493 G.n4129 G.t2579 120.189
R3494 G.n4130 G.t3591 120.189
R3495 G.n570 G.t2094 120.189
R3496 G.n637 G.t3927 120.189
R3497 G.n707 G.t1966 120.189
R3498 G.n780 G.t3463 120.189
R3499 G.n856 G.t1405 120.189
R3500 G.n938 G.t2900 120.189
R3501 G.n1023 G.t905 120.189
R3502 G.n1111 G.t2381 120.189
R3503 G.n1199 G.t441 120.189
R3504 G.n1287 G.t1924 120.189
R3505 G.n1375 G.t4388 120.189
R3506 G.n1463 G.t1364 120.189
R3507 G.n1550 G.t3879 120.189
R3508 G.n1633 G.t394 120.189
R3509 G.n1711 G.t3414 120.189
R3510 G.n1783 G.t4351 120.189
R3511 G.n1851 G.t2860 120.189
R3512 G.n1915 G.t3833 120.189
R3513 G.n2659 G.t2340 120.189
R3514 G.n2658 G.t751 120.189
R3515 G.n2657 G.t3769 120.189
R3516 G.n2656 G.t260 120.189
R3517 G.n2655 G.t2743 120.189
R3518 G.n2654 G.t4240 120.189
R3519 G.n2653 G.t2232 120.189
R3520 G.n2652 G.t3729 120.189
R3521 G.n2651 G.t1740 120.189
R3522 G.n2650 G.t3229 120.189
R3523 G.n2649 G.t1218 120.189
R3524 G.n2615 G.t2401 120.189
R3525 G.n2616 G.t4408 120.189
R3526 G.n2617 G.t2918 120.189
R3527 G.n2618 G.t467 120.189
R3528 G.n2619 G.t3482 120.189
R3529 G.n2620 G.t928 120.189
R3530 G.n2621 G.t3941 120.189
R3531 G.n2622 G.t1430 120.189
R3532 G.n2623 G.t509 120.189
R3533 G.n2624 G.t1995 120.189
R3534 G.n2625 G.t3588 120.189
R3535 G.n1917 G.t570 120.189
R3536 G.n1854 G.t4075 120.189
R3537 G.n1786 G.t1052 120.189
R3538 G.n1714 G.t59 120.189
R3539 G.n1636 G.t1553 120.189
R3540 G.n1553 G.t608 120.189
R3541 G.n1466 G.t2580 120.189
R3542 G.n1378 G.t1098 120.189
R3543 G.n1290 G.t3083 120.189
R3544 G.n1202 G.t1596 120.189
R3545 G.n1114 G.t3626 120.189
R3546 G.n1026 G.t2130 120.189
R3547 G.n941 G.t4124 120.189
R3548 G.n859 G.t2627 120.189
R3549 G.n783 G.t115 120.189
R3550 G.n710 G.t3141 120.189
R3551 G.n640 G.t649 120.189
R3552 G.n573 G.t3302 120.189
R3553 G.n509 G.t279 120.189
R3554 G.n4077 G.t3786 120.189
R3555 G.n4076 G.t765 120.189
R3556 G.n4075 G.t4292 120.189
R3557 G.n4074 G.t1277 120.189
R3558 G.n4073 G.t327 120.189
R3559 G.n4072 G.t1817 120.189
R3560 G.n4071 G.t803 120.189
R3561 G.n4070 G.t2805 120.189
R3562 G.n4069 G.t1316 120.189
R3563 G.n4068 G.t3352 120.189
R3564 G.n4067 G.t1865 120.189
R3565 G.n4066 G.t3819 120.189
R3566 G.n4065 G.t2325 120.189
R3567 G.n4064 G.t4341 120.189
R3568 G.n4063 G.t2847 120.189
R3569 G.n4062 G.t702 120.189
R3570 G.n4061 G.t3835 120.189
R3571 G.n4012 G.t4376 120.189
R3572 G.n4013 G.t1073 120.189
R3573 G.n4014 G.t1121 120.189
R3574 G.n4015 G.t2400 120.189
R3575 G.n4016 G.t4127 120.189
R3576 G.n4017 G.t906 120.189
R3577 G.n4018 G.t2613 120.189
R3578 G.n4019 G.t3908 120.189
R3579 G.n4020 G.t1114 120.189
R3580 G.n4021 G.t2390 120.189
R3581 G.n4022 G.t4115 120.189
R3582 G.n4023 G.t2418 120.189
R3583 G.n4024 G.t2602 120.189
R3584 G.n4025 G.t920 120.189
R3585 G.n4026 G.t1103 120.189
R3586 G.n4027 G.t3923 120.189
R3587 G.n451 G.t4108 120.189
R3588 G.n512 G.t2403 120.189
R3589 G.n576 G.t2592 120.189
R3590 G.n643 G.t53 120.189
R3591 G.n713 G.t1782 120.189
R3592 G.n786 G.t3053 120.189
R3593 G.n862 G.t281 120.189
R3594 G.n944 G.t1554 120.189
R3595 G.n1029 G.t3284 120.189
R3596 G.n1117 G.t46 120.189
R3597 G.n1205 G.t1776 120.189
R3598 G.n1293 G.t3045 120.189
R3599 G.n1381 G.t275 120.189
R3600 G.n1469 G.t1546 120.189
R3601 G.n1556 G.t3277 120.189
R3602 G.n1639 G.t1573 120.189
R3603 G.n1717 G.t1762 120.189
R3604 G.n1789 G.t61 120.189
R3605 G.n1857 G.t263 120.189
R3606 G.n1919 G.t3063 120.189
R3607 G.n1977 G.t3266 120.189
R3608 G.n2593 G.t1064 120.189
R3609 G.n2592 G.t1231 120.189
R3610 G.n2591 G.t4070 120.189
R3611 G.n2590 G.t1256 120.189
R3612 G.n2589 G.t2553 120.189
R3613 G.n2588 G.t4257 120.189
R3614 G.n2587 G.t1053 120.189
R3615 G.n2586 G.t2747 120.189
R3616 G.n2585 G.t4059 120.189
R3617 G.n2584 G.t1242 120.189
R3618 G.n2554 G.t2676 120.189
R3619 G.n2555 G.t969 120.189
R3620 G.n2556 G.t4185 120.189
R3621 G.n2557 G.t2471 120.189
R3622 G.n2558 G.t1183 120.189
R3623 G.n2559 G.t3983 120.189
R3624 G.n2560 G.t2685 120.189
R3625 G.n2561 G.t976 120.189
R3626 G.n2562 G.t2666 120.189
R3627 G.n2563 G.t2476 120.189
R3628 G.n1979 G.t170 120.189
R3629 G.n1922 G.t4492 120.189
R3630 G.n1860 G.t1676 120.189
R3631 G.n1792 G.t1487 120.189
R3632 G.n1720 G.t3185 120.189
R3633 G.n1642 G.t2994 120.189
R3634 G.n1559 G.t186 120.189
R3635 G.n1472 G.t2969 120.189
R3636 G.n1384 G.t1688 120.189
R3637 G.n1296 G.t4476 120.189
R3638 G.n1208 G.t3198 120.189
R3639 G.n1120 G.t1468 120.189
R3640 G.n1032 G.t197 120.189
R3641 G.n947 G.t2979 120.189
R3642 G.n865 G.t1694 120.189
R3643 G.n789 G.t4488 120.189
R3644 G.n716 G.t3208 120.189
R3645 G.n646 G.t1481 120.189
R3646 G.n579 G.t4028 120.189
R3647 G.n515 G.t3845 120.189
R3648 G.n454 G.t1019 120.189
R3649 G.n396 G.t841 120.189
R3650 G.n3980 G.t2520 120.189
R3651 G.n3979 G.t2344 120.189
R3652 G.n3978 G.t4037 120.189
R3653 G.n3977 G.t3859 120.189
R3654 G.n3976 G.t1030 120.189
R3655 G.n3975 G.t3827 120.189
R3656 G.n3974 G.t2529 120.189
R3657 G.n3973 G.t828 120.189
R3658 G.n3972 G.t4043 120.189
R3659 G.n3971 G.t2324 120.189
R3660 G.n3970 G.t1037 120.189
R3661 G.n3969 G.t3837 120.189
R3662 G.n3968 G.t2538 120.189
R3663 G.n3967 G.t2487 120.189
R3664 G.n3966 G.t1304 120.189
R3665 G.n3920 G.t1412 120.189
R3666 G.n3921 G.t2619 120.189
R3667 G.n3922 G.t2669 120.189
R3668 G.n3923 G.t3961 120.189
R3669 G.n3924 G.t1168 120.189
R3670 G.n3925 G.t2452 120.189
R3671 G.n3926 G.t4168 120.189
R3672 G.n3927 G.t951 120.189
R3673 G.n3928 G.t2661 120.189
R3674 G.n3929 G.t3951 120.189
R3675 G.n3930 G.t1157 120.189
R3676 G.n3931 G.t3977 120.189
R3677 G.n3932 G.t4157 120.189
R3678 G.n3933 G.t2467 120.189
R3679 G.n3934 G.t2649 120.189
R3680 G.n399 G.t966 120.189
R3681 G.n457 G.t1150 120.189
R3682 G.n518 G.t3967 120.189
R3683 G.n582 G.t4149 120.189
R3684 G.n649 G.t1615 120.189
R3685 G.n719 G.t3348 120.189
R3686 G.n792 G.t108 120.189
R3687 G.n868 G.t1837 120.189
R3688 G.n950 G.t3107 120.189
R3689 G.n1035 G.t336 120.189
R3690 G.n1123 G.t1603 120.189
R3691 G.n1211 G.t3340 120.189
R3692 G.n1299 G.t97 120.189
R3693 G.n1387 G.t1828 120.189
R3694 G.n1475 G.t3095 120.189
R3695 G.n1562 G.t324 120.189
R3696 G.n1645 G.t3132 120.189
R3697 G.n1723 G.t3331 120.189
R3698 G.n1795 G.t1621 120.189
R3699 G.n1863 G.t1821 120.189
R3700 G.n1925 G.t117 120.189
R3701 G.n1982 G.t317 120.189
R3702 G.n2034 G.t2614 120.189
R3703 G.n2534 G.t2778 120.189
R3704 G.n2533 G.t1115 120.189
R3705 G.n2532 G.t2801 120.189
R3706 G.n2531 G.t4116 120.189
R3707 G.n2530 G.t1295 120.189
R3708 G.n2529 G.t2603 120.189
R3709 G.n2528 G.t4298 120.189
R3710 G.n2527 G.t1104 120.189
R3711 G.n2526 G.t2789 120.189
R3712 G.n2499 G.t4232 120.189
R3713 G.n2500 G.t2521 120.189
R3714 G.n2501 G.t1224 120.189
R3715 G.n2502 G.t4034 120.189
R3716 G.n2503 G.t2729 120.189
R3717 G.n2504 G.t1031 120.189
R3718 G.n2505 G.t4237 120.189
R3719 G.n2506 G.t2530 120.189
R3720 G.n2507 G.t4221 120.189
R3721 G.n2036 G.t4044 120.189
R3722 G.n1985 G.t1729 120.189
R3723 G.n1928 G.t1538 120.189
R3724 G.n1866 G.t3244 120.189
R3725 G.n1798 G.t3038 120.189
R3726 G.n1726 G.t242 120.189
R3727 G.n1648 G.t37 120.189
R3728 G.n1565 G.t1741 120.189
R3729 G.n1478 G.t16 120.189
R3730 G.n1390 G.t3253 120.189
R3731 G.n1302 G.t1524 120.189
R3732 G.n1214 G.t249 120.189
R3733 G.n1126 G.t3025 120.189
R3734 G.n1038 G.t1750 120.189
R3735 G.n953 G.t25 120.189
R3736 G.n871 G.t3259 120.189
R3737 G.n795 G.t1535 120.189
R3738 G.n722 G.t258 120.189
R3739 G.n652 G.t3033 120.189
R3740 G.n585 G.t1077 120.189
R3741 G.n521 G.t890 120.189
R3742 G.n460 G.t2571 120.189
R3743 G.n402 G.t2384 120.189
R3744 G.n347 G.t4083 120.189
R3745 G.n3890 G.t3902 120.189
R3746 G.n3889 G.t1083 120.189
R3747 G.n3888 G.t898 120.189
R3748 G.n3887 G.t2581 120.189
R3749 G.n3886 G.t874 120.189
R3750 G.n3885 G.t4093 120.189
R3751 G.n3884 G.t2373 120.189
R3752 G.n3883 G.t1090 120.189
R3753 G.n3882 G.t3888 120.189
R3754 G.n3881 G.t2587 120.189
R3755 G.n3880 G.t883 120.189
R3756 G.n3879 G.t4102 120.189
R3757 G.n3878 G.t4053 120.189
R3758 G.n3877 G.t2852 120.189
R3759 G.n3837 G.t2965 120.189
R3760 G.n3838 G.t4176 120.189
R3761 G.n3839 G.t4225 120.189
R3762 G.n3840 G.t1008 120.189
R3763 G.n3841 G.t2711 120.189
R3764 G.n3842 G.t4014 120.189
R3765 G.n3843 G.t1210 120.189
R3766 G.n3844 G.t2499 120.189
R3767 G.n3845 G.t4219 120.189
R3768 G.n3846 G.t994 120.189
R3769 G.n3847 G.t2703 120.189
R3770 G.n3848 G.t1027 120.189
R3771 G.n3849 G.t1204 120.189
R3772 G.n301 G.t4031 120.189
R3773 G.n350 G.t4203 120.189
R3774 G.n405 G.t2515 120.189
R3775 G.n463 G.t2695 120.189
R3776 G.n524 G.t1013 120.189
R3777 G.n588 G.t1195 120.189
R3778 G.n655 G.t3178 120.189
R3779 G.n725 G.t398 120.189
R3780 G.n798 G.t1666 120.189
R3781 G.n874 G.t3402 120.189
R3782 G.n956 G.t160 120.189
R3783 G.n1041 G.t1891 120.189
R3784 G.n1129 G.t3165 120.189
R3785 G.n1217 G.t389 120.189
R3786 G.n1305 G.t1657 120.189
R3787 G.n1393 G.t3390 120.189
R3788 G.n1481 G.t152 120.189
R3789 G.n1568 G.t1881 120.189
R3790 G.n1651 G.t181 120.189
R3791 G.n1729 G.t380 120.189
R3792 G.n1801 G.t3181 120.189
R3793 G.n1869 G.t3381 120.189
R3794 G.n1931 G.t1673 120.189
R3795 G.n1988 G.t1873 120.189
R3796 G.n2039 G.t4170 120.189
R3797 G.n2085 G.t4333 120.189
R3798 G.n2481 G.t2663 120.189
R3799 G.n2480 G.t4355 120.189
R3800 G.n2479 G.t1159 120.189
R3801 G.n2478 G.t2846 120.189
R3802 G.n2477 G.t4159 120.189
R3803 G.n2476 G.t1338 120.189
R3804 G.n2475 G.t2651 120.189
R3805 G.n2474 G.t4346 120.189
R3806 G.n2452 G.t1271 120.189
R3807 G.n2453 G.t4084 120.189
R3808 G.n2454 G.t2767 120.189
R3809 G.n2455 G.t1084 120.189
R3810 G.n2456 G.t4282 120.189
R3811 G.n2457 G.t2582 120.189
R3812 G.n2458 G.t1276 120.189
R3813 G.n2130 G.t4094 120.189
R3814 G.n2087 G.t1258 120.189
R3815 G.n2042 G.t1092 120.189
R3816 G.n1991 G.t3296 120.189
R3817 G.n1934 G.t3089 120.189
R3818 G.n1872 G.t295 120.189
R3819 G.n1804 G.t87 120.189
R3820 G.n1732 G.t1795 120.189
R3821 G.n1654 G.t1595 120.189
R3822 G.n1571 G.t3310 120.189
R3823 G.n1484 G.t1578 120.189
R3824 G.n1396 G.t306 120.189
R3825 G.n1308 G.t3078 120.189
R3826 G.n1220 G.t1808 120.189
R3827 G.n1132 G.t72 120.189
R3828 G.n1044 G.t3317 120.189
R3829 G.n959 G.t1585 120.189
R3830 G.n877 G.t312 120.189
R3831 G.n801 G.t3084 120.189
R3832 G.n728 G.t1816 120.189
R3833 G.n658 G.t81 120.189
R3834 G.n591 G.t2624 120.189
R3835 G.n527 G.t2432 120.189
R3836 G.n466 G.t4133 120.189
R3837 G.n408 G.t3943 120.189
R3838 G.n353 G.t1127 120.189
R3839 G.n304 G.t945 120.189
R3840 G.n258 G.t2631 120.189
R3841 G.n3811 G.t2448 120.189
R3842 G.n3810 G.t4143 120.189
R3843 G.n3809 G.t2421 120.189
R3844 G.n3808 G.t1136 120.189
R3845 G.n3807 G.t3936 120.189
R3846 G.n3806 G.t2641 120.189
R3847 G.n3805 G.t930 120.189
R3848 G.n3804 G.t4146 120.189
R3849 G.n3803 G.t2427 120.189
R3850 G.n3802 G.t1143 120.189
R3851 G.n3801 G.t1096 120.189
R3852 G.n3800 G.t4399 120.189
R3853 G.n3766 G.t9 120.189
R3854 G.n3767 G.t1217 120.189
R3855 G.n3768 G.t1261 120.189
R3856 G.n3769 G.t2563 120.189
R3857 G.n3770 G.t4264 120.189
R3858 G.n3771 G.t1060 120.189
R3859 G.n3772 G.t2754 120.189
R3860 G.n3773 G.t4066 120.189
R3861 G.n3774 G.t1254 120.189
R3862 G.n3775 G.t2549 120.189
R3863 G.n3776 G.t4255 120.189
R3864 G.n218 G.t2577 120.189
R3865 G.n261 G.t2746 120.189
R3866 G.n307 G.t1079 120.189
R3867 G.n356 G.t1244 120.189
R3868 G.n411 G.t4080 120.189
R3869 G.n469 G.t4249 120.189
R3870 G.n530 G.t2569 120.189
R3871 G.n594 G.t2739 120.189
R3872 G.n661 G.t232 120.189
R3873 G.n731 G.t1945 120.189
R3874 G.n804 G.t3231 120.189
R3875 G.n880 G.t448 120.189
R3876 G.n962 G.t1717 120.189
R3877 G.n1047 G.t3452 120.189
R3878 G.n1135 G.t216 120.189
R3879 G.n1223 G.t1940 120.189
R3880 G.n1311 G.t3222 120.189
R3881 G.n1399 G.t440 120.189
R3882 G.n1487 G.t1708 120.189
R3883 G.n1574 G.t3441 120.189
R3884 G.n1657 G.t1736 120.189
R3885 G.n1735 G.t1932 120.189
R3886 G.n1807 G.t235 120.189
R3887 G.n1875 G.t430 120.189
R3888 G.n1937 G.t3233 120.189
R3889 G.n1994 G.t3433 120.189
R3890 G.n2045 G.t1209 120.189
R3891 G.n2090 G.t1365 120.189
R3892 G.n2132 G.t4215 120.189
R3893 G.n2436 G.t1388 120.189
R3894 G.n2435 G.t2702 120.189
R3895 G.n2434 G.t4395 120.189
R3896 G.n2433 G.t1203 120.189
R3897 G.n2432 G.t2890 120.189
R3898 G.n2431 G.t4202 120.189
R3899 G.n2430 G.t1380 120.189
R3900 G.n2411 G.t2818 120.189
R3901 G.n2412 G.t1126 120.189
R3902 G.n2413 G.t4320 120.189
R3903 G.n2414 G.t2630 120.189
R3904 G.n2415 G.t1321 120.189
R3905 G.n2416 G.t4142 120.189
R3906 G.n2171 G.t2825 120.189
R3907 G.n2134 G.t1135 120.189
R3908 G.n2093 G.t2803 120.189
R3909 G.n2048 G.t2640 120.189
R3910 G.n1997 G.t348 120.189
R3911 G.n1940 G.t145 120.189
R3912 G.n1878 G.t1853 120.189
R3913 G.n1810 G.t1645 120.189
R3914 G.n1738 G.t3360 120.189
R3915 G.n1660 G.t3157 120.189
R3916 G.n1577 G.t360 120.189
R3917 G.n1490 G.t3134 120.189
R3918 G.n1402 G.t1863 120.189
R3919 G.n1314 G.t130 120.189
R3920 G.n1226 G.t3369 120.189
R3921 G.n1138 G.t1628 120.189
R3922 G.n1050 G.t365 120.189
R3923 G.n965 G.t3143 120.189
R3924 G.n883 G.t1868 120.189
R3925 G.n807 G.t138 120.189
R3926 G.n734 G.t3376 120.189
R3927 G.n664 G.t1640 120.189
R3928 G.n597 G.t4178 120.189
R3929 G.n533 G.t3996 120.189
R3930 G.n472 G.t1173 120.189
R3931 G.n414 G.t987 120.189
R3932 G.n359 G.t2673 120.189
R3933 G.n310 G.t2496 120.189
R3934 G.n264 G.t4183 120.189
R3935 G.n221 G.t4010 120.189
R3936 G.n181 G.t1182 120.189
R3937 G.n3744 G.t3981 120.189
R3938 G.n3743 G.t2683 120.189
R3939 G.n3742 G.t975 120.189
R3940 G.n3741 G.t4192 120.189
R3941 G.n3740 G.t2477 120.189
R3942 G.n3739 G.t1188 120.189
R3943 G.n3738 G.t3988 120.189
R3944 G.n3737 G.t2689 120.189
R3945 G.n3736 G.t2645 120.189
R3946 G.n3735 G.t1438 120.189
R3947 G.n3707 G.t1569 120.189
R3948 G.n3708 G.t2760 120.189
R3949 G.n3709 G.t2807 120.189
R3950 G.n3710 G.t4125 120.189
R3951 G.n3711 G.t1305 120.189
R3952 G.n3712 G.t2609 120.189
R3953 G.n3713 G.t4306 120.189
R3954 G.n3714 G.t1111 120.189
R3955 G.n3715 G.t2800 120.189
R3956 G.n147 G.t4113 120.189
R3957 G.n184 G.t1294 120.189
R3958 G.n224 G.t4137 120.189
R3959 G.n267 G.t4297 120.189
R3960 G.n313 G.t2626 120.189
R3961 G.n362 G.t2787 120.189
R3962 G.n417 G.t1122 120.189
R3963 G.n475 G.t1284 120.189
R3964 G.n536 G.t4130 120.189
R3965 G.n600 G.t4290 120.189
R3966 G.n667 G.t1779 120.189
R3967 G.n737 G.t3507 120.189
R3968 G.n810 G.t283 120.189
R3969 G.n886 G.t1998 120.189
R3970 G.n968 G.t3286 120.189
R3971 G.n1053 G.t499 120.189
R3972 G.n1141 G.t1773 120.189
R3973 G.n1229 G.t3499 120.189
R3974 G.n1317 G.t273 120.189
R3975 G.n1405 G.t1990 120.189
R3976 G.n1493 G.t3274 120.189
R3977 G.n1580 G.t486 120.189
R3978 G.n1663 G.t3303 120.189
R3979 G.n1741 G.t3488 120.189
R3980 G.n1813 G.t1788 120.189
R3981 G.n1881 G.t1980 120.189
R3982 G.n1943 G.t286 120.189
R3983 G.n2000 G.t479 120.189
R3984 G.n2051 G.t2753 120.189
R3985 G.n2096 G.t2916 120.189
R3986 G.n2137 G.t1253 120.189
R3987 G.n2173 G.t2938 120.189
R3988 G.n2397 G.t4254 120.189
R3989 G.n2396 G.t1433 120.189
R3990 G.n2395 G.t2745 120.189
R3991 G.n2394 G.t4439 120.189
R3992 G.n2393 G.t1241 120.189
R3993 G.n2392 G.t2933 120.189
R3994 G.n2376 G.t4153 120.189
R3995 G.n2377 G.t2436 120.189
R3996 G.n2378 G.t1155 120.189
R3997 G.n2379 G.t3945 120.189
R3998 G.n2380 G.t2653 120.189
R3999 G.n2206 G.t946 120.189
R4000 G.n2175 G.t4162 120.189
R4001 G.n2140 G.t2447 120.189
R4002 G.n2099 G.t4141 120.189
R4003 G.n2054 G.t3954 120.189
R4004 G.n2003 G.t1637 120.189
R4005 G.n1946 G.t1449 120.189
R4006 G.n1884 G.t3150 120.189
R4007 G.n1816 G.t2955 120.189
R4008 G.n1744 G.t144 120.189
R4009 G.n1666 G.t4465 120.189
R4010 G.n1583 G.t1644 120.189
R4011 G.n1496 G.t4445 120.189
R4012 G.n1408 G.t3156 120.189
R4013 G.n1320 G.t1440 120.189
R4014 G.n1232 G.t155 120.189
R4015 G.n1144 G.t2944 120.189
R4016 G.n1056 G.t1659 120.189
R4017 G.n971 G.t4449 120.189
R4018 G.n889 G.t3167 120.189
R4019 G.n813 G.t1448 120.189
R4020 G.n740 G.t163 120.189
R4021 G.n670 G.t2953 120.189
R4022 G.n603 G.t981 120.189
R4023 G.n539 G.t816 120.189
R4024 G.n478 G.t2488 120.189
R4025 G.n420 G.t2306 120.189
R4026 G.n365 G.t3995 120.189
R4027 G.n316 G.t3818 120.189
R4028 G.n270 G.t986 120.189
R4029 G.n227 G.t822 120.189
R4030 G.n187 G.t2495 120.189
R4031 G.n150 G.t800 120.189
R4032 G.n116 G.t4009 120.189
R4033 G.n3689 G.t2292 120.189
R4034 G.n3688 G.t999 120.189
R4035 G.n3687 G.t3802 120.189
R4036 G.n3686 G.t2503 120.189
R4037 G.n3685 G.t806 120.189
R4038 G.n3684 G.t4017 120.189
R4039 G.n3683 G.t3962 120.189
R4040 G.n3682 G.t2773 120.189
R4041 G.n3657 G.t3124 120.189
R4042 G.n3658 G.t4311 120.189
R4043 G.n3659 G.t4359 120.189
R4044 G.n3660 G.t1165 120.189
R4045 G.n3661 G.t2854 120.189
R4046 G.n3662 G.t4164 120.189
R4047 G.n3663 G.t1343 120.189
R4048 G.n3664 G.t2658 120.189
R4049 G.n119 G.t4354 120.189
R4050 G.n153 G.t1156 120.189
R4051 G.n190 G.t2844 120.189
R4052 G.n230 G.t1178 120.189
R4053 G.n273 G.t1336 120.189
R4054 G.n319 G.t4181 120.189
R4055 G.n368 G.t4343 120.189
R4056 G.n423 G.t2670 120.189
R4057 G.n481 G.t2837 120.189
R4058 G.n542 G.t1169 120.189
R4059 G.n606 G.t1330 120.189
R4060 G.n673 G.t3347 120.189
R4061 G.n743 G.t543 120.189
R4062 G.n816 G.t1835 120.189
R4063 G.n892 G.t3551 120.189
R4064 G.n974 G.t335 120.189
R4065 G.n1059 G.t2041 120.189
R4066 G.n1147 G.t3337 120.189
R4067 G.n1235 G.t538 120.189
R4068 G.n1323 G.t1830 120.189
R4069 G.n1411 G.t3544 120.189
R4070 G.n1499 G.t326 120.189
R4071 G.n1586 G.t2029 120.189
R4072 G.n1669 G.t354 120.189
R4073 G.n1747 G.t530 120.189
R4074 G.n1819 G.t3353 120.189
R4075 G.n1887 G.t3534 120.189
R4076 G.n1949 G.t1844 120.189
R4077 G.n2006 G.t2021 120.189
R4078 G.n2057 G.t4305 120.189
R4079 G.n2102 G.t4467 120.189
R4080 G.n2143 G.t2799 120.189
R4081 G.n2178 G.t4493 120.189
R4082 G.n2208 G.t1293 120.189
R4083 G.n2365 G.t2986 120.189
R4084 G.n2364 G.t4296 120.189
R4085 G.n2363 G.t1476 120.189
R4086 G.n2362 G.t2786 120.189
R4087 G.n2361 G.t4484 120.189
R4088 G.n2348 G.t1199 120.189
R4089 G.n2349 G.t3994 120.189
R4090 G.n2350 G.t2699 120.189
R4091 G.n2351 G.t985 120.189
R4092 G.n2236 G.t4201 120.189
R4093 G.n2211 G.t2494 120.189
R4094 G.n2181 G.t1202 120.189
R4095 G.n2146 G.t4008 120.189
R4096 G.n2105 G.t1181 120.189
R4097 G.n2060 G.t998 120.189
R4098 G.n2009 G.t3205 120.189
R4099 G.n1952 G.t3006 120.189
R4100 G.n1890 G.t201 120.189
R4101 G.n1822 G.t0 120.189
R4102 G.n1750 G.t1700 120.189
R4103 G.n1672 G.t1510 120.189
R4104 G.n1589 G.t3212 120.189
R4105 G.n1502 G.t1488 120.189
R4106 G.n1414 G.t209 120.189
R4107 G.n1326 G.t2996 120.189
R4108 G.n1238 G.t1712 120.189
R4109 G.n1150 G.t4502 120.189
R4110 G.n1062 G.t3224 120.189
R4111 G.n977 G.t1495 120.189
R4112 G.n895 G.t219 120.189
R4113 G.n819 G.t3005 120.189
R4114 G.n746 G.t1720 120.189
R4115 G.n676 G.t4510 120.189
R4116 G.n609 G.t2536 120.189
R4117 G.n545 G.t2359 120.189
R4118 G.n484 G.t4051 120.189
R4119 G.n426 G.t3866 120.189
R4120 G.n371 G.t1044 120.189
R4121 G.n322 G.t863 120.189
R4122 G.n276 G.t2545 120.189
R4123 G.n233 G.t2364 120.189
R4124 G.n193 G.t4062 120.189
R4125 G.n156 G.t2342 120.189
R4126 G.n122 G.t1055 120.189
R4127 G.n91 G.t3855 120.189
R4128 G.n3641 G.t2555 120.189
R4129 G.n3640 G.t848 120.189
R4130 G.n3639 G.t4071 120.189
R4131 G.n3638 G.t2349 120.189
R4132 G.n3637 G.t1066 120.189
R4133 G.n3636 G.t1007 120.189
R4134 G.n3635 G.t4326 120.189
R4135 G.n3616 G.t176 120.189
R4136 G.n3617 G.t1346 120.189
R4137 G.n3618 G.t1395 120.189
R4138 G.n3619 G.t2710 120.189
R4139 G.n3620 G.t4401 120.189
R4140 G.n3621 G.t1208 120.189
R4141 G.n69 G.t2897 120.189
R4142 G.n94 G.t4214 120.189
R4143 G.n125 G.t1387 120.189
R4144 G.n159 G.t2700 120.189
R4145 G.n196 G.t4393 120.189
R4146 G.n236 G.t2724 120.189
R4147 G.n279 G.t2889 120.189
R4148 G.n325 G.t1219 120.189
R4149 G.n374 G.t1377 120.189
R4150 G.n429 G.t4226 120.189
R4151 G.n487 G.t4384 120.189
R4152 G.n548 G.t2715 120.189
R4153 G.n612 G.t2881 120.189
R4154 G.n679 G.t397 120.189
R4155 G.n749 G.t2083 120.189
R4156 G.n822 G.t3399 120.189
R4157 G.n898 G.t583 120.189
R4158 G.n980 G.t1889 120.189
R4159 G.n1065 G.t3587 120.189
R4160 G.n1153 G.t386 120.189
R4161 G.n1241 G.t2078 120.189
R4162 G.n1329 G.t3388 120.189
R4163 G.n1417 G.t575 120.189
R4164 G.n1505 G.t1880 120.189
R4165 G.n1592 G.t3578 120.189
R4166 G.n1675 G.t1904 120.189
R4167 G.n1753 G.t2070 120.189
R4168 G.n1825 G.t400 120.189
R4169 G.n1893 G.t568 120.189
R4170 G.n1955 G.t3407 120.189
R4171 G.n2012 G.t3574 120.189
R4172 G.n2063 G.t1342 120.189
R4173 G.n2108 G.t1513 120.189
R4174 G.n2149 G.t4353 120.189
R4175 G.n2184 G.t1537 120.189
R4176 G.n2214 G.t2843 120.189
R4177 G.n2238 G.t29 120.189
R4178 G.n2260 G.t1335 120.189
R4179 G.n2340 G.t3029 120.189
R4180 G.n2339 G.t4342 120.189
R4181 G.n2338 G.t1530 120.189
R4182 G.n2328 G.t2738 120.189
R4183 G.n2329 G.t1043 120.189
R4184 G.n2330 G.t4248 120.189
R4185 G.n2262 G.t2544 120.189
R4186 G.n2241 G.t1243 120.189
R4187 G.n2217 G.t4061 120.189
R4188 G.n2187 G.t2748 120.189
R4189 G.n2152 G.t1054 120.189
R4190 G.n2111 G.t2727 120.189
R4191 G.n2066 G.t2554 120.189
R4192 G.n2015 G.t255 120.189
R4193 G.n1958 G.t50 120.189
R4194 G.n1896 G.t1754 120.189
R4195 G.n1828 G.t1558 120.189
R4196 G.n1756 G.t3267 120.189
R4197 G.n1678 G.t3064 120.189
R4198 G.n1595 G.t264 120.189
R4199 G.n1508 G.t3037 120.189
R4200 G.n1420 G.t1764 120.189
R4201 G.n1332 G.t36 120.189
R4202 G.n1244 G.t3278 120.189
R4203 G.n1156 G.t1544 120.189
R4204 G.n1068 G.t277 120.189
R4205 G.n983 G.t3046 120.189
R4206 G.n901 G.t1772 120.189
R4207 G.n825 G.t47 120.189
R4208 G.n752 G.t3285 120.189
R4209 G.n682 G.t1555 120.189
R4210 G.n615 G.t4099 120.189
R4211 G.n551 G.t3915 120.189
R4212 G.n490 G.t1095 120.189
R4213 G.n432 G.t910 120.189
R4214 G.n377 G.t2594 120.189
R4215 G.n328 G.t2405 120.189
R4216 G.n282 G.t4110 120.189
R4217 G.n239 G.t3925 120.189
R4218 G.n199 G.t1106 120.189
R4219 G.n162 G.t3904 120.189
R4220 G.n128 G.t2605 120.189
R4221 G.n97 G.t899 120.189
R4222 G.n72 G.t4118 120.189
R4223 G.n50 G.t2391 120.189
R4224 G.n3604 G.t1116 120.189
R4225 G.n3603 G.t3909 120.189
R4226 G.n3602 G.t2615 120.189
R4227 G.n3601 G.t2562 120.189
R4228 G.n3600 G.t1359 120.189
R4229 G.n3587 G.t1731 120.189
R4230 G.n3588 G.t2901 120.189
R4231 G.n3589 G.t2941 120.189
R4232 G.n3590 G.t4261 120.189
R4233 G.n34 G.t1437 120.189
R4234 G.n53 G.t2751 120.189
R4235 G.n75 G.t4444 120.189
R4236 G.n100 G.t1250 120.189
R4237 G.n131 G.t2937 120.189
R4238 G.n165 G.t4253 120.189
R4239 G.n202 G.t1432 120.189
R4240 G.n242 G.t4276 120.189
R4241 G.n285 G.t4436 120.189
R4242 G.n331 G.t2761 120.189
R4243 G.n380 G.t2931 120.189
R4244 G.n435 G.t1264 120.189
R4245 G.n493 G.t1423 120.189
R4246 G.n554 G.t4268 120.189
R4247 G.n618 G.t4428 120.189
R4248 G.n685 G.t1944 120.189
R4249 G.n755 G.t3631 120.189
R4250 G.n828 G.t446 120.189
R4251 G.n904 G.t2124 120.189
R4252 G.n986 G.t3448 120.189
R4253 G.n1071 G.t623 120.189
R4254 G.n1159 G.t1937 120.189
R4255 G.n1247 G.t3623 120.189
R4256 G.n1335 G.t436 120.189
R4257 G.n1423 G.t2118 120.189
R4258 G.n1511 G.t3439 120.189
R4259 G.n1598 G.t613 120.189
R4260 G.n1681 G.t3465 120.189
R4261 G.n1759 G.t3619 120.189
R4262 G.n1831 G.t1948 120.189
R4263 G.n1899 G.t2109 120.189
R4264 G.n1961 G.t453 120.189
R4265 G.n2018 G.t609 120.189
R4266 G.n2069 G.t2896 120.189
R4267 G.n2114 G.t3068 120.189
R4268 G.n2155 G.t1386 120.189
R4269 G.n2190 G.t3088 120.189
R4270 G.n2220 G.t4392 120.189
R4271 G.n2244 G.t1588 120.189
R4272 G.n2264 G.t2888 120.189
R4273 G.n2280 G.t75 120.189
R4274 G.n2322 G.t1376 120.189
R4275 G.n2321 G.t3080 120.189
R4276 G.n2314 G.t4291 120.189
R4277 G.n2315 G.t2593 120.189
R4278 G.n2282 G.t1286 120.189
R4279 G.n2267 G.t4109 120.189
R4280 G.n2247 G.t2790 120.189
R4281 G.n2223 G.t1105 120.189
R4282 G.n2193 G.t4299 120.189
R4283 G.n2158 G.t2604 120.189
R4284 G.n2117 G.t4281 120.189
R4285 G.n2072 G.t4117 120.189
R4286 G.n2021 G.t1813 120.189
R4287 G.n1964 G.t1611 120.189
R4288 G.n1902 G.t3323 120.189
R4289 G.n1834 G.t3115 120.189
R4290 G.n1762 G.t318 120.189
R4291 G.n1684 G.t119 120.189
R4292 G.n1601 G.t1822 120.189
R4293 G.n1514 G.t85 120.189
R4294 G.n1426 G.t3327 120.189
R4295 G.n1338 G.t1593 120.189
R4296 G.n1250 G.t325 120.189
R4297 G.n1162 G.t3097 120.189
R4298 G.n1074 G.t1829 120.189
R4299 G.n989 G.t99 120.189
R4300 G.n907 G.t3341 120.189
R4301 G.n831 G.t1604 120.189
R4302 G.n758 G.t337 120.189
R4303 G.n688 G.t3108 120.189
R4304 G.n621 G.t1140 120.189
R4305 G.n557 G.t960 120.189
R4306 G.n496 G.t2644 120.189
R4307 G.n438 G.t2457 120.189
R4308 G.n383 G.t4150 120.189
R4309 G.n334 G.t3968 120.189
R4310 G.n288 G.t1151 120.189
R4311 G.n245 G.t967 120.189
R4312 G.n205 G.t2650 120.189
R4313 G.n168 G.t943 120.189
R4314 G.n134 G.t4158 120.189
R4315 G.n103 G.t2445 120.189
R4316 G.n78 G.t1158 120.189
R4317 G.n56 G.t3952 120.189
R4318 G.n37 G.t2662 120.189
R4319 G.n21 G.t952 120.189
R4320 G.n3579 G.t4169 120.189
R4321 G.n3578 G.t4121 120.189
R4322 G.n3577 G.t2913 120.189
R4323 G.n3570 G.t3298 120.189
R4324 G.n3571 G.t4447 120.189
R4325 G.n11 G.t4496 120.189
R4326 G.n24 G.t1300 120.189
R4327 G.n40 G.t2990 120.189
R4328 G.n59 G.t4302 120.189
R4329 G.n81 G.t1484 120.189
R4330 G.n106 G.t2795 120.189
R4331 G.n137 G.t4490 120.189
R4332 G.n171 G.t1291 120.189
R4333 G.n208 G.t2981 120.189
R4334 G.n248 G.t1314 120.189
R4335 G.n291 G.t1475 120.189
R4336 G.n337 G.t4314 120.189
R4337 G.n386 G.t4483 120.189
R4338 G.n441 G.t2813 120.189
R4339 G.n499 G.t2974 120.189
R4340 G.n560 G.t1309 120.189
R4341 G.n624 G.t1466 120.189
R4342 G.n691 G.t3504 120.189
R4343 G.n761 G.t667 120.189
R4344 G.n834 G.t1996 120.189
R4345 G.n910 G.t3674 120.189
R4346 G.n992 G.t495 120.189
R4347 G.n1077 G.t2165 120.189
R4348 G.n1165 G.t3496 120.189
R4349 G.n1253 G.t659 120.189
R4350 G.n1341 G.t1987 120.189
R4351 G.n1429 G.t3667 120.189
R4352 G.n1517 G.t484 120.189
R4353 G.n1604 G.t2154 120.189
R4354 G.n1687 G.t507 120.189
R4355 G.n1765 G.t657 120.189
R4356 G.n1837 G.t3509 120.189
R4357 G.n1905 G.t3660 120.189
R4358 G.n1967 G.t2001 120.189
R4359 G.n2024 G.t2148 120.189
R4360 G.n2075 G.t4442 120.189
R4361 G.n2120 G.t118 120.189
R4362 G.n2161 G.t2936 120.189
R4363 G.n2196 G.t143 120.189
R4364 G.n2226 G.t1431 120.189
R4365 G.n2250 G.t3149 120.189
R4366 G.n2270 G.t4435 120.189
R4367 G.n2284 G.t1636 120.189
R4368 G.n2294 G.t2930 120.189
R4369 G.n2310 G.t135 120.189
R4370 G.n2307 G.t4063 120.189
R4371 G.n2296 G.t2995 120.189
R4372 G.n2287 G.t2026 120.189
R4373 G.n2273 G.t938 120.189
R4374 G.n2253 G.t4426 120.189
R4375 G.n2229 G.t3427 120.189
R4376 G.n2199 G.t2361 120.189
R4377 G.n2164 G.t1317 120.189
R4378 G.n2123 G.t1426 120.189
R4379 G.n2078 G.t3766 120.189
R4380 G.n2027 G.t2345 120.189
R4381 G.n1970 G.t187 120.189
R4382 G.n1908 G.t320 120.189
R4383 G.n1840 G.t2623 120.189
R4384 G.n1768 G.t2733 120.189
R4385 G.n1690 G.t585 120.189
R4386 G.n1607 G.t684 120.189
R4387 G.n1520 G.t4139 120.189
R4388 G.n1432 G.t3113 120.189
R4389 G.n1344 G.t2091 120.189
R4390 G.n1256 G.t1056 120.189
R4391 G.n1168 G.t4501 120.189
R4392 G.n1080 G.t3540 120.189
R4393 G.n995 G.t2430 120.189
R4394 G.n913 G.t1421 120.189
R4395 G.n837 G.t422 120.189
R4396 G.n764 G.t3872 120.189
R4397 G.n694 G.t2824 120.189
R4398 G.n627 G.t3054 120.189
R4399 G.n563 G.t880 120.189
R4400 G.n502 G.t997 120.189
R4401 G.n444 G.t3366 120.189
R4402 G.n389 G.t3490 120.189
R4403 G.n340 G.t1268 120.189
R4404 G.n294 G.t1372 120.189
R4405 G.n251 G.t3715 120.189
R4406 G.n211 G.t3817 120.189
R4407 G.n174 G.t2772 120.189
R4408 G.n140 G.t1783 120.189
R4409 G.n109 G.t715 120.189
R4410 G.n84 G.t4218 120.189
R4411 G.n62 G.t3163 120.189
R4412 G.n43 G.t2160 120.189
R4413 G.n27 G.t1100 120.189
R4414 G.n14 G.t71 120.189
R4415 G.n4 G.t2057 120.189
R4416 G.n3566 G.t3903 120.189
R4417 G.n3 G.t2809 120.189
R4418 G.n0 G.t3305 120.189
R4419 G.n10 G.t4001 120.189
R4420 G.n7 G.t2798 120.189
R4421 G.n20 G.t4060 120.189
R4422 G.n17 G.t459 120.189
R4423 G.n33 G.t838 120.189
R4424 G.n30 G.t3188 120.189
R4425 G.n49 G.t2543 120.189
R4426 G.n46 G.t2404 120.189
R4427 G.n68 G.t3843 120.189
R4428 G.n65 G.t690 120.189
R4429 G.n90 G.t1042 120.189
R4430 G.n87 G.t4416 120.189
R4431 G.n115 G.t2331 120.189
R4432 G.n112 G.t2682 120.189
R4433 G.n146 G.t4050 120.189
R4434 G.n143 G.t1963 120.189
R4435 G.n180 G.t831 120.189
R4436 G.n177 G.t193 120.189
R4437 G.n217 G.t2535 120.189
R4438 G.n214 G.t3928 120.189
R4439 G.n257 G.t856 120.189
R4440 G.n254 G.t3394 120.189
R4441 G.n300 G.t1034 120.189
R4442 G.n297 G.t1415 120.189
R4443 G.n346 G.t3860 120.189
R4444 G.n343 G.t842 120.189
R4445 G.n395 G.t4039 120.189
R4446 G.n392 G.t3478 120.189
R4447 G.n450 G.t2346 120.189
R4448 G.n447 G.t2853 120.189
R4449 G.n508 G.t2522 120.189
R4450 G.n505 G.t929 120.189
R4451 G.n569 G.t843 120.189
R4452 G.n566 G.t396 120.189
R4453 G.n633 G.t1023 120.189
R4454 G.n630 G.t2927 120.189
R4455 G.n700 G.t2992 120.189
R4456 G.n697 G.t2744 120.189
R4457 G.n770 G.t206 120.189
R4458 G.n767 G.t2027 120.189
R4459 G.n843 G.t1485 120.189
R4460 G.n840 G.t265 120.189
R4461 G.n919 G.t3210 120.189
R4462 G.n916 G.t3989 120.189
R4463 G.n1001 G.t4491 120.189
R4464 G.n998 G.t2241 120.189
R4465 G.n1086 G.t1696 120.189
R4466 G.n1083 G.t1482 120.189
R4467 G.n1174 G.t2982 120.189
R4468 G.n1171 G.t4258 120.189
R4469 G.n1262 G.t198 120.189
R4470 G.n1259 G.t3543 120.189
R4471 G.n1350 G.t1471 120.189
R4472 G.n1347 G.t1771 120.189
R4473 G.n1438 G.t3204 120.189
R4474 G.n1435 G.t989 120.189
R4475 G.n1526 G.t4480 120.189
R4476 G.n1523 G.t3763 120.189
R4477 G.n1613 G.t1691 120.189
R4478 G.n1610 G.t2991 120.189
R4479 G.n1696 G.t4508 120.189
R4480 G.n1693 G.t2409 120.189
R4481 G.n1774 G.t191 120.189
R4482 G.n1771 G.t542 120.189
R4483 G.n1846 G.t3003 120.189
R4484 G.n1843 G.t4420 120.189
R4485 G.n1914 G.t3192 120.189
R4486 G.n1911 G.t2498 120.189
R4487 G.n1976 G.t1491 120.189
R4488 G.n1973 G.t1969 120.189
R4489 G.n2033 G.t1681 120.189
R4490 G.n2030 G.t4505 120.189
R4491 G.n2084 G.t3993 120.189
R4492 G.n2081 G.t2802 120.189
R4493 G.n2129 G.t4177 120.189
R4494 G.n2126 G.t871 120.189
R4495 G.n2170 G.t2484 120.189
R4496 G.n2167 G.t334 120.189
R4497 G.n2205 G.t4196 120.189
R4498 G.n2202 G.t4064 120.189
R4499 G.n2235 G.t980 120.189
R4500 G.n2232 G.t2297 120.189
R4501 G.n2259 G.t2687 120.189
R4502 G.n2256 G.t1543 120.189
R4503 G.n2279 G.t3985 120.189
R4504 G.n2276 G.t4310 120.189
R4505 G.n2293 G.t1185 120.189
R4506 G.n2290 G.t3589 120.189
R4507 G.n2302 G.t2473 120.189
R4508 G.n2299 G.t1840 120.189
R4509 G.n2305 G.t4189 120.189
R4510 G.n2303 G.t1058 120.189
R4511 G.n6814 G.t1722 120.189
R4512 G.n3456 G.n3455 0.686
R4513 G.n3454 G.n3453 0.686
R4514 G.n6778 G.n6774 0.686
R4515 G.n6763 G.n6756 0.686
R4516 G.n6745 G.n6735 0.686
R4517 G.n6724 G.n6711 0.686
R4518 G.n6700 G.n6684 0.686
R4519 G.n6673 G.n6654 0.686
R4520 G.n6643 G.n6621 0.686
R4521 G.n6610 G.n6584 0.686
R4522 G.n6573 G.n6543 0.686
R4523 G.n6532 G.n6499 0.686
R4524 G.n6488 G.n6451 0.686
R4525 G.n6440 G.n6400 0.686
R4526 G.n6389 G.n6347 0.686
R4527 G.n6336 G.n6293 0.686
R4528 G.n6282 G.n6239 0.686
R4529 G.n6228 G.n6185 0.686
R4530 G.n6174 G.n6131 0.686
R4531 G.n6120 G.n6079 0.686
R4532 G.n6068 G.n6028 0.686
R4533 G.n6017 G.n5979 0.686
R4534 G.n5968 G.n5933 0.686
R4535 G.n5922 G.n5888 0.686
R4536 G.n5877 G.n5845 0.686
R4537 G.n5834 G.n5805 0.686
R4538 G.n5794 G.n5766 0.686
R4539 G.n5755 G.n5729 0.686
R4540 G.n5718 G.n5695 0.686
R4541 G.n5684 G.n5664 0.686
R4542 G.n5653 G.n5633 0.686
R4543 G.n5622 G.n5605 0.686
R4544 G.n5594 G.n5580 0.686
R4545 G.n5569 G.n5555 0.686
R4546 G.n5544 G.n5533 0.686
R4547 G.n5522 G.n5514 0.686
R4548 G.n5503 G.n5496 0.686
R4549 G.n5485 G.n5480 0.686
R4550 G.n5469 G.n5467 0.686
R4551 G.n5456 G.n5455 0.686
R4552 G.n5390 G.n5389 0.686
R4553 G.n5393 G.n5391 0.686
R4554 G.n5396 G.n5394 0.686
R4555 G.n5399 G.n5397 0.686
R4556 G.n5402 G.n5400 0.686
R4557 G.n3448 G.n3447 0.686
R4558 G.n3446 G.n3445 0.686
R4559 G.n3444 G.n3443 0.686
R4560 G.n3442 G.n3441 0.686
R4561 G.n5376 G.n5375 0.686
R4562 G.n5378 G.n5377 0.686
R4563 G.n5380 G.n5379 0.686
R4564 G.n5382 G.n5381 0.686
R4565 G.n5384 G.n5383 0.686
R4566 G.n5386 G.n5385 0.686
R4567 G.n3435 G.n3434 0.686
R4568 G.n3433 G.n3432 0.686
R4569 G.n3431 G.n3430 0.686
R4570 G.n3429 G.n3428 0.686
R4571 G.n6740 G.n6736 0.686
R4572 G.n6719 G.n6712 0.686
R4573 G.n6695 G.n6685 0.686
R4574 G.n6668 G.n6655 0.686
R4575 G.n6638 G.n6622 0.686
R4576 G.n6605 G.n6585 0.686
R4577 G.n6568 G.n6544 0.686
R4578 G.n6527 G.n6500 0.686
R4579 G.n6483 G.n6452 0.686
R4580 G.n6435 G.n6401 0.686
R4581 G.n6384 G.n6348 0.686
R4582 G.n6331 G.n6294 0.686
R4583 G.n6277 G.n6240 0.686
R4584 G.n6223 G.n6186 0.686
R4585 G.n6169 G.n6132 0.686
R4586 G.n6115 G.n6080 0.686
R4587 G.n6063 G.n6029 0.686
R4588 G.n6012 G.n5980 0.686
R4589 G.n5963 G.n5934 0.686
R4590 G.n5917 G.n5889 0.686
R4591 G.n5872 G.n5846 0.686
R4592 G.n5829 G.n5806 0.686
R4593 G.n5789 G.n5767 0.686
R4594 G.n5750 G.n5730 0.686
R4595 G.n5713 G.n5696 0.686
R4596 G.n5679 G.n5665 0.686
R4597 G.n5648 G.n5634 0.686
R4598 G.n5617 G.n5606 0.686
R4599 G.n5589 G.n5581 0.686
R4600 G.n5564 G.n5556 0.686
R4601 G.n5539 G.n5534 0.686
R4602 G.n5517 G.n5515 0.686
R4603 G.n5498 G.n5497 0.686
R4604 G.n5352 G.n5351 0.686
R4605 G.n5354 G.n5353 0.686
R4606 G.n5356 G.n5355 0.686
R4607 G.n5358 G.n5357 0.686
R4608 G.n5360 G.n5359 0.686
R4609 G.n5362 G.n5361 0.686
R4610 G.n5364 G.n5363 0.686
R4611 G.n5366 G.n5365 0.686
R4612 G.n3421 G.n3420 0.686
R4613 G.n3419 G.n3418 0.686
R4614 G.n3417 G.n3416 0.686
R4615 G.n3415 G.n3414 0.686
R4616 G.n3413 G.n3412 0.686
R4617 G.n3411 G.n3410 0.686
R4618 G.n5325 G.n5324 0.686
R4619 G.n5327 G.n5326 0.686
R4620 G.n5329 G.n5328 0.686
R4621 G.n5331 G.n5330 0.686
R4622 G.n5333 G.n5332 0.686
R4623 G.n5335 G.n5334 0.686
R4624 G.n5337 G.n5336 0.686
R4625 G.n5339 G.n5338 0.686
R4626 G.n5341 G.n5340 0.686
R4627 G.n3402 G.n3401 0.686
R4628 G.n3400 G.n3399 0.686
R4629 G.n3398 G.n3397 0.686
R4630 G.n3396 G.n3395 0.686
R4631 G.n3394 G.n3393 0.686
R4632 G.n3392 G.n3391 0.686
R4633 G.n6690 G.n6686 0.686
R4634 G.n6663 G.n6656 0.686
R4635 G.n6633 G.n6623 0.686
R4636 G.n6600 G.n6586 0.686
R4637 G.n6563 G.n6545 0.686
R4638 G.n6522 G.n6501 0.686
R4639 G.n6478 G.n6453 0.686
R4640 G.n6430 G.n6402 0.686
R4641 G.n6379 G.n6349 0.686
R4642 G.n6326 G.n6295 0.686
R4643 G.n6272 G.n6241 0.686
R4644 G.n6218 G.n6187 0.686
R4645 G.n6164 G.n6133 0.686
R4646 G.n6110 G.n6081 0.686
R4647 G.n6058 G.n6030 0.686
R4648 G.n6007 G.n5981 0.686
R4649 G.n5958 G.n5935 0.686
R4650 G.n5912 G.n5890 0.686
R4651 G.n5867 G.n5847 0.686
R4652 G.n5824 G.n5807 0.686
R4653 G.n5784 G.n5768 0.686
R4654 G.n5745 G.n5731 0.686
R4655 G.n5708 G.n5697 0.686
R4656 G.n5674 G.n5666 0.686
R4657 G.n5643 G.n5635 0.686
R4658 G.n5612 G.n5607 0.686
R4659 G.n5584 G.n5582 0.686
R4660 G.n5559 G.n5557 0.686
R4661 G.n5292 G.n5291 0.686
R4662 G.n5294 G.n5293 0.686
R4663 G.n5296 G.n5295 0.686
R4664 G.n5298 G.n5297 0.686
R4665 G.n5300 G.n5299 0.686
R4666 G.n5302 G.n5301 0.686
R4667 G.n5304 G.n5303 0.686
R4668 G.n5306 G.n5305 0.686
R4669 G.n5308 G.n5307 0.686
R4670 G.n5310 G.n5309 0.686
R4671 G.n5312 G.n5311 0.686
R4672 G.n3382 G.n3381 0.686
R4673 G.n3380 G.n3379 0.686
R4674 G.n3378 G.n3377 0.686
R4675 G.n3376 G.n3375 0.686
R4676 G.n3374 G.n3373 0.686
R4677 G.n3372 G.n3371 0.686
R4678 G.n3370 G.n3369 0.686
R4679 G.n3368 G.n3367 0.686
R4680 G.n5256 G.n5255 0.686
R4681 G.n5258 G.n5257 0.686
R4682 G.n5260 G.n5259 0.686
R4683 G.n5262 G.n5261 0.686
R4684 G.n5264 G.n5263 0.686
R4685 G.n5266 G.n5265 0.686
R4686 G.n5268 G.n5267 0.686
R4687 G.n5270 G.n5269 0.686
R4688 G.n5272 G.n5271 0.686
R4689 G.n5274 G.n5273 0.686
R4690 G.n5276 G.n5275 0.686
R4691 G.n5278 G.n5277 0.686
R4692 G.n3357 G.n3356 0.686
R4693 G.n3355 G.n3354 0.686
R4694 G.n3353 G.n3352 0.686
R4695 G.n3351 G.n3350 0.686
R4696 G.n3349 G.n3348 0.686
R4697 G.n3347 G.n3346 0.686
R4698 G.n3345 G.n3344 0.686
R4699 G.n3343 G.n3342 0.686
R4700 G.n6628 G.n6624 0.686
R4701 G.n6595 G.n6587 0.686
R4702 G.n6558 G.n6546 0.686
R4703 G.n6517 G.n6502 0.686
R4704 G.n6473 G.n6454 0.686
R4705 G.n6425 G.n6403 0.686
R4706 G.n6374 G.n6350 0.686
R4707 G.n6321 G.n6296 0.686
R4708 G.n6267 G.n6242 0.686
R4709 G.n6213 G.n6188 0.686
R4710 G.n6159 G.n6134 0.686
R4711 G.n6105 G.n6082 0.686
R4712 G.n6053 G.n6031 0.686
R4713 G.n6002 G.n5982 0.686
R4714 G.n5953 G.n5936 0.686
R4715 G.n5907 G.n5891 0.686
R4716 G.n5862 G.n5848 0.686
R4717 G.n5819 G.n5808 0.686
R4718 G.n5779 G.n5769 0.686
R4719 G.n5740 G.n5732 0.686
R4720 G.n5703 G.n5698 0.686
R4721 G.n5669 G.n5667 0.686
R4722 G.n5638 G.n5636 0.686
R4723 G.n5215 G.n5214 0.686
R4724 G.n5217 G.n5216 0.686
R4725 G.n5219 G.n5218 0.686
R4726 G.n5221 G.n5220 0.686
R4727 G.n5223 G.n5222 0.686
R4728 G.n5225 G.n5224 0.686
R4729 G.n5227 G.n5226 0.686
R4730 G.n5229 G.n5228 0.686
R4731 G.n5231 G.n5230 0.686
R4732 G.n5233 G.n5232 0.686
R4733 G.n5235 G.n5234 0.686
R4734 G.n5237 G.n5236 0.686
R4735 G.n5239 G.n5238 0.686
R4736 G.n5241 G.n5240 0.686
R4737 G.n3331 G.n3330 0.686
R4738 G.n3329 G.n3328 0.686
R4739 G.n3327 G.n3326 0.686
R4740 G.n3325 G.n3324 0.686
R4741 G.n3323 G.n3322 0.686
R4742 G.n3321 G.n3320 0.686
R4743 G.n3319 G.n3318 0.686
R4744 G.n3317 G.n3316 0.686
R4745 G.n3315 G.n3314 0.686
R4746 G.n3313 G.n3312 0.686
R4747 G.n5170 G.n5169 0.686
R4748 G.n5172 G.n5171 0.686
R4749 G.n5174 G.n5173 0.686
R4750 G.n5176 G.n5175 0.686
R4751 G.n5178 G.n5177 0.686
R4752 G.n5180 G.n5179 0.686
R4753 G.n5182 G.n5181 0.686
R4754 G.n5184 G.n5183 0.686
R4755 G.n5186 G.n5185 0.686
R4756 G.n5188 G.n5187 0.686
R4757 G.n5190 G.n5189 0.686
R4758 G.n5192 G.n5191 0.686
R4759 G.n5194 G.n5193 0.686
R4760 G.n5196 G.n5195 0.686
R4761 G.n5198 G.n5197 0.686
R4762 G.n3300 G.n3299 0.686
R4763 G.n3298 G.n3297 0.686
R4764 G.n3296 G.n3295 0.686
R4765 G.n3294 G.n3293 0.686
R4766 G.n3292 G.n3291 0.686
R4767 G.n3290 G.n3289 0.686
R4768 G.n3288 G.n3287 0.686
R4769 G.n3286 G.n3285 0.686
R4770 G.n3284 G.n3283 0.686
R4771 G.n3282 G.n3281 0.686
R4772 G.n6590 G.n6588 0.686
R4773 G.n6553 G.n6547 0.686
R4774 G.n6512 G.n6503 0.686
R4775 G.n6468 G.n6455 0.686
R4776 G.n6420 G.n6404 0.686
R4777 G.n6369 G.n6351 0.686
R4778 G.n6316 G.n6297 0.686
R4779 G.n6262 G.n6243 0.686
R4780 G.n6208 G.n6189 0.686
R4781 G.n6154 G.n6135 0.686
R4782 G.n6100 G.n6083 0.686
R4783 G.n6048 G.n6032 0.686
R4784 G.n5997 G.n5983 0.686
R4785 G.n5948 G.n5937 0.686
R4786 G.n5902 G.n5892 0.686
R4787 G.n5857 G.n5849 0.686
R4788 G.n5814 G.n5809 0.686
R4789 G.n5774 G.n5770 0.686
R4790 G.n5735 G.n5733 0.686
R4791 G.n5120 G.n5119 0.686
R4792 G.n5122 G.n5121 0.686
R4793 G.n5124 G.n5123 0.686
R4794 G.n5126 G.n5125 0.686
R4795 G.n5128 G.n5127 0.686
R4796 G.n5130 G.n5129 0.686
R4797 G.n5132 G.n5131 0.686
R4798 G.n5134 G.n5133 0.686
R4799 G.n5136 G.n5135 0.686
R4800 G.n5138 G.n5137 0.686
R4801 G.n5140 G.n5139 0.686
R4802 G.n5142 G.n5141 0.686
R4803 G.n5144 G.n5143 0.686
R4804 G.n5146 G.n5145 0.686
R4805 G.n5148 G.n5147 0.686
R4806 G.n5150 G.n5149 0.686
R4807 G.n5152 G.n5151 0.686
R4808 G.n3269 G.n3268 0.686
R4809 G.n3267 G.n3266 0.686
R4810 G.n3265 G.n3264 0.686
R4811 G.n3263 G.n3262 0.686
R4812 G.n3261 G.n3260 0.686
R4813 G.n3259 G.n3258 0.686
R4814 G.n3257 G.n3256 0.686
R4815 G.n3255 G.n3254 0.686
R4816 G.n3253 G.n3252 0.686
R4817 G.n3251 G.n3250 0.686
R4818 G.n3249 G.n3248 0.686
R4819 G.n5068 G.n5067 0.686
R4820 G.n5070 G.n5069 0.686
R4821 G.n5072 G.n5071 0.686
R4822 G.n5074 G.n5073 0.686
R4823 G.n5076 G.n5075 0.686
R4824 G.n5078 G.n5077 0.686
R4825 G.n5080 G.n5079 0.686
R4826 G.n5082 G.n5081 0.686
R4827 G.n5084 G.n5083 0.686
R4828 G.n5086 G.n5085 0.686
R4829 G.n5088 G.n5087 0.686
R4830 G.n5090 G.n5089 0.686
R4831 G.n5092 G.n5091 0.686
R4832 G.n5094 G.n5093 0.686
R4833 G.n5096 G.n5095 0.686
R4834 G.n5098 G.n5097 0.686
R4835 G.n5100 G.n5099 0.686
R4836 G.n3233 G.n3232 0.686
R4837 G.n3231 G.n3230 0.686
R4838 G.n3229 G.n3228 0.686
R4839 G.n3227 G.n3226 0.686
R4840 G.n3225 G.n3224 0.686
R4841 G.n3223 G.n3222 0.686
R4842 G.n3221 G.n3220 0.686
R4843 G.n3219 G.n3218 0.686
R4844 G.n3217 G.n3216 0.686
R4845 G.n3215 G.n3214 0.686
R4846 G.n3213 G.n3212 0.686
R4847 G.n6507 G.n6504 0.686
R4848 G.n6463 G.n6456 0.686
R4849 G.n6415 G.n6405 0.686
R4850 G.n6364 G.n6352 0.686
R4851 G.n6311 G.n6298 0.686
R4852 G.n6257 G.n6244 0.686
R4853 G.n6203 G.n6190 0.686
R4854 G.n6149 G.n6136 0.686
R4855 G.n6095 G.n6084 0.686
R4856 G.n6043 G.n6033 0.686
R4857 G.n5992 G.n5984 0.686
R4858 G.n5943 G.n5938 0.686
R4859 G.n5897 G.n5893 0.686
R4860 G.n5852 G.n5850 0.686
R4861 G.n5009 G.n5008 0.686
R4862 G.n5011 G.n5010 0.686
R4863 G.n5013 G.n5012 0.686
R4864 G.n5015 G.n5014 0.686
R4865 G.n5017 G.n5016 0.686
R4866 G.n5019 G.n5018 0.686
R4867 G.n5021 G.n5020 0.686
R4868 G.n5023 G.n5022 0.686
R4869 G.n5025 G.n5024 0.686
R4870 G.n5027 G.n5026 0.686
R4871 G.n5029 G.n5028 0.686
R4872 G.n5031 G.n5030 0.686
R4873 G.n5033 G.n5032 0.686
R4874 G.n5035 G.n5034 0.686
R4875 G.n5037 G.n5036 0.686
R4876 G.n5039 G.n5038 0.686
R4877 G.n5041 G.n5040 0.686
R4878 G.n5043 G.n5042 0.686
R4879 G.n5045 G.n5044 0.686
R4880 G.n5047 G.n5046 0.686
R4881 G.n3197 G.n3196 0.686
R4882 G.n3195 G.n3194 0.686
R4883 G.n3193 G.n3192 0.686
R4884 G.n3191 G.n3190 0.686
R4885 G.n3189 G.n3188 0.686
R4886 G.n3187 G.n3186 0.686
R4887 G.n3185 G.n3184 0.686
R4888 G.n3183 G.n3182 0.686
R4889 G.n3181 G.n3180 0.686
R4890 G.n3179 G.n3178 0.686
R4891 G.n3177 G.n3176 0.686
R4892 G.n3175 G.n3174 0.686
R4893 G.n3173 G.n3172 0.686
R4894 G.n4948 G.n4947 0.686
R4895 G.n4950 G.n4949 0.686
R4896 G.n4952 G.n4951 0.686
R4897 G.n4954 G.n4953 0.686
R4898 G.n4956 G.n4955 0.686
R4899 G.n4958 G.n4957 0.686
R4900 G.n4960 G.n4959 0.686
R4901 G.n4962 G.n4961 0.686
R4902 G.n4964 G.n4963 0.686
R4903 G.n4966 G.n4965 0.686
R4904 G.n4968 G.n4967 0.686
R4905 G.n4970 G.n4969 0.686
R4906 G.n4972 G.n4971 0.686
R4907 G.n4974 G.n4973 0.686
R4908 G.n4976 G.n4975 0.686
R4909 G.n4978 G.n4977 0.686
R4910 G.n4980 G.n4979 0.686
R4911 G.n4982 G.n4981 0.686
R4912 G.n4984 G.n4983 0.686
R4913 G.n4986 G.n4985 0.686
R4914 G.n3156 G.n3155 0.686
R4915 G.n3154 G.n3153 0.686
R4916 G.n3152 G.n3151 0.686
R4917 G.n3150 G.n3149 0.686
R4918 G.n3148 G.n3147 0.686
R4919 G.n3146 G.n3145 0.686
R4920 G.n3144 G.n3143 0.686
R4921 G.n3142 G.n3141 0.686
R4922 G.n3140 G.n3139 0.686
R4923 G.n3138 G.n3137 0.686
R4924 G.n3136 G.n3135 0.686
R4925 G.n3134 G.n3133 0.686
R4926 G.n3132 G.n3131 0.686
R4927 G.n6410 G.n6406 0.686
R4928 G.n6359 G.n6353 0.686
R4929 G.n6306 G.n6299 0.686
R4930 G.n6252 G.n6245 0.686
R4931 G.n6198 G.n6191 0.686
R4932 G.n6144 G.n6137 0.686
R4933 G.n6090 G.n6085 0.686
R4934 G.n6038 G.n6034 0.686
R4935 G.n5987 G.n5985 0.686
R4936 G.n4880 G.n4879 0.686
R4937 G.n4882 G.n4881 0.686
R4938 G.n4884 G.n4883 0.686
R4939 G.n4886 G.n4885 0.686
R4940 G.n4888 G.n4887 0.686
R4941 G.n4890 G.n4889 0.686
R4942 G.n4892 G.n4891 0.686
R4943 G.n4894 G.n4893 0.686
R4944 G.n4896 G.n4895 0.686
R4945 G.n4898 G.n4897 0.686
R4946 G.n4900 G.n4899 0.686
R4947 G.n4902 G.n4901 0.686
R4948 G.n4904 G.n4903 0.686
R4949 G.n4906 G.n4905 0.686
R4950 G.n4908 G.n4907 0.686
R4951 G.n4910 G.n4909 0.686
R4952 G.n4912 G.n4911 0.686
R4953 G.n4914 G.n4913 0.686
R4954 G.n4916 G.n4915 0.686
R4955 G.n4918 G.n4917 0.686
R4956 G.n4920 G.n4919 0.686
R4957 G.n4922 G.n4921 0.686
R4958 G.n4924 G.n4923 0.686
R4959 G.n3114 G.n3113 0.686
R4960 G.n3112 G.n3111 0.686
R4961 G.n3110 G.n3109 0.686
R4962 G.n3108 G.n3107 0.686
R4963 G.n3106 G.n3105 0.686
R4964 G.n3104 G.n3103 0.686
R4965 G.n3102 G.n3101 0.686
R4966 G.n3100 G.n3099 0.686
R4967 G.n3098 G.n3097 0.686
R4968 G.n3096 G.n3095 0.686
R4969 G.n3094 G.n3093 0.686
R4970 G.n3092 G.n3091 0.686
R4971 G.n3090 G.n3089 0.686
R4972 G.n3088 G.n3087 0.686
R4973 G.n3086 G.n3085 0.686
R4974 G.n4810 G.n4809 0.686
R4975 G.n4812 G.n4811 0.686
R4976 G.n4814 G.n4813 0.686
R4977 G.n4816 G.n4815 0.686
R4978 G.n4818 G.n4817 0.686
R4979 G.n4820 G.n4819 0.686
R4980 G.n4822 G.n4821 0.686
R4981 G.n4824 G.n4823 0.686
R4982 G.n4826 G.n4825 0.686
R4983 G.n4828 G.n4827 0.686
R4984 G.n4830 G.n4829 0.686
R4985 G.n4832 G.n4831 0.686
R4986 G.n4834 G.n4833 0.686
R4987 G.n4836 G.n4835 0.686
R4988 G.n4838 G.n4837 0.686
R4989 G.n4840 G.n4839 0.686
R4990 G.n4842 G.n4841 0.686
R4991 G.n4844 G.n4843 0.686
R4992 G.n4846 G.n4845 0.686
R4993 G.n4848 G.n4847 0.686
R4994 G.n4850 G.n4849 0.686
R4995 G.n4852 G.n4851 0.686
R4996 G.n4854 G.n4853 0.686
R4997 G.n3068 G.n3067 0.686
R4998 G.n3066 G.n3065 0.686
R4999 G.n3064 G.n3063 0.686
R5000 G.n3062 G.n3061 0.686
R5001 G.n3060 G.n3059 0.686
R5002 G.n3058 G.n3057 0.686
R5003 G.n3056 G.n3055 0.686
R5004 G.n3054 G.n3053 0.686
R5005 G.n3052 G.n3051 0.686
R5006 G.n3050 G.n3049 0.686
R5007 G.n3048 G.n3047 0.686
R5008 G.n3046 G.n3045 0.686
R5009 G.n3044 G.n3043 0.686
R5010 G.n3042 G.n3041 0.686
R5011 G.n3040 G.n3039 0.686
R5012 G.n6301 G.n6300 0.686
R5013 G.n6247 G.n6246 0.686
R5014 G.n6193 G.n6192 0.686
R5015 G.n6139 G.n6138 0.686
R5016 G.n4733 G.n4732 0.686
R5017 G.n4735 G.n4734 0.686
R5018 G.n4737 G.n4736 0.686
R5019 G.n4739 G.n4738 0.686
R5020 G.n4741 G.n4740 0.686
R5021 G.n4743 G.n4742 0.686
R5022 G.n4745 G.n4744 0.686
R5023 G.n4747 G.n4746 0.686
R5024 G.n4749 G.n4748 0.686
R5025 G.n4751 G.n4750 0.686
R5026 G.n4753 G.n4752 0.686
R5027 G.n4755 G.n4754 0.686
R5028 G.n4757 G.n4756 0.686
R5029 G.n4759 G.n4758 0.686
R5030 G.n4761 G.n4760 0.686
R5031 G.n4763 G.n4762 0.686
R5032 G.n4765 G.n4764 0.686
R5033 G.n4767 G.n4766 0.686
R5034 G.n4769 G.n4768 0.686
R5035 G.n4771 G.n4770 0.686
R5036 G.n4773 G.n4772 0.686
R5037 G.n4775 G.n4774 0.686
R5038 G.n4777 G.n4776 0.686
R5039 G.n4779 G.n4778 0.686
R5040 G.n4781 G.n4780 0.686
R5041 G.n4783 G.n4782 0.686
R5042 G.n3021 G.n3020 0.686
R5043 G.n3019 G.n3018 0.686
R5044 G.n3017 G.n3016 0.686
R5045 G.n3015 G.n3014 0.686
R5046 G.n3013 G.n3012 0.686
R5047 G.n3011 G.n3010 0.686
R5048 G.n3009 G.n3008 0.686
R5049 G.n3007 G.n3006 0.686
R5050 G.n3005 G.n3004 0.686
R5051 G.n3003 G.n3002 0.686
R5052 G.n3001 G.n3000 0.686
R5053 G.n2999 G.n2998 0.686
R5054 G.n2997 G.n2996 0.686
R5055 G.n2995 G.n2994 0.686
R5056 G.n2993 G.n2992 0.686
R5057 G.n2991 G.n2990 0.686
R5058 G.n4658 G.n4657 0.686
R5059 G.n4660 G.n4659 0.686
R5060 G.n4662 G.n4661 0.686
R5061 G.n4664 G.n4663 0.686
R5062 G.n4666 G.n4665 0.686
R5063 G.n4668 G.n4667 0.686
R5064 G.n4670 G.n4669 0.686
R5065 G.n4672 G.n4671 0.686
R5066 G.n4674 G.n4673 0.686
R5067 G.n4676 G.n4675 0.686
R5068 G.n4678 G.n4677 0.686
R5069 G.n4680 G.n4679 0.686
R5070 G.n4682 G.n4681 0.686
R5071 G.n4684 G.n4683 0.686
R5072 G.n4686 G.n4685 0.686
R5073 G.n4688 G.n4687 0.686
R5074 G.n4690 G.n4689 0.686
R5075 G.n4692 G.n4691 0.686
R5076 G.n4694 G.n4693 0.686
R5077 G.n4696 G.n4695 0.686
R5078 G.n4698 G.n4697 0.686
R5079 G.n4700 G.n4699 0.686
R5080 G.n4702 G.n4701 0.686
R5081 G.n4704 G.n4703 0.686
R5082 G.n2971 G.n2970 0.686
R5083 G.n2969 G.n2968 0.686
R5084 G.n2967 G.n2966 0.686
R5085 G.n2965 G.n2964 0.686
R5086 G.n2963 G.n2962 0.686
R5087 G.n2961 G.n2960 0.686
R5088 G.n2959 G.n2958 0.686
R5089 G.n2957 G.n2956 0.686
R5090 G.n2955 G.n2954 0.686
R5091 G.n2953 G.n2952 0.686
R5092 G.n2951 G.n2950 0.686
R5093 G.n2949 G.n2948 0.686
R5094 G.n2947 G.n2946 0.686
R5095 G.n2945 G.n2944 0.686
R5096 G.n1531 G.n1530 0.686
R5097 G.n1444 G.n1443 0.686
R5098 G.n1356 G.n1355 0.686
R5099 G.n1268 G.n1267 0.686
R5100 G.n1180 G.n1179 0.686
R5101 G.n1092 G.n1091 0.686
R5102 G.n1004 G.n1003 0.686
R5103 G.n4583 G.n4582 0.686
R5104 G.n4585 G.n4584 0.686
R5105 G.n4587 G.n4586 0.686
R5106 G.n4589 G.n4588 0.686
R5107 G.n4591 G.n4590 0.686
R5108 G.n4593 G.n4592 0.686
R5109 G.n4595 G.n4594 0.686
R5110 G.n4597 G.n4596 0.686
R5111 G.n4599 G.n4598 0.686
R5112 G.n4601 G.n4600 0.686
R5113 G.n4603 G.n4602 0.686
R5114 G.n4605 G.n4604 0.686
R5115 G.n4607 G.n4606 0.686
R5116 G.n4609 G.n4608 0.686
R5117 G.n4611 G.n4610 0.686
R5118 G.n4613 G.n4612 0.686
R5119 G.n4615 G.n4614 0.686
R5120 G.n4617 G.n4616 0.686
R5121 G.n4619 G.n4618 0.686
R5122 G.n4621 G.n4620 0.686
R5123 G.n4623 G.n4622 0.686
R5124 G.n4625 G.n4624 0.686
R5125 G.n4627 G.n4626 0.686
R5126 G.n4629 G.n4628 0.686
R5127 G.n2926 G.n2925 0.686
R5128 G.n2924 G.n2923 0.686
R5129 G.n2922 G.n2921 0.686
R5130 G.n2920 G.n2919 0.686
R5131 G.n2918 G.n2917 0.686
R5132 G.n2916 G.n2915 0.686
R5133 G.n2914 G.n2913 0.686
R5134 G.n2912 G.n2911 0.686
R5135 G.n2910 G.n2909 0.686
R5136 G.n2908 G.n2907 0.686
R5137 G.n2906 G.n2905 0.686
R5138 G.n2904 G.n2903 0.686
R5139 G.n2902 G.n2901 0.686
R5140 G.n2900 G.n2899 0.686
R5141 G.n2898 G.n2897 0.686
R5142 G.n4513 G.n4512 0.686
R5143 G.n4515 G.n4514 0.686
R5144 G.n4517 G.n4516 0.686
R5145 G.n4519 G.n4518 0.686
R5146 G.n4521 G.n4520 0.686
R5147 G.n4523 G.n4522 0.686
R5148 G.n4525 G.n4524 0.686
R5149 G.n4527 G.n4526 0.686
R5150 G.n4529 G.n4528 0.686
R5151 G.n4531 G.n4530 0.686
R5152 G.n4533 G.n4532 0.686
R5153 G.n4535 G.n4534 0.686
R5154 G.n4537 G.n4536 0.686
R5155 G.n4539 G.n4538 0.686
R5156 G.n4541 G.n4540 0.686
R5157 G.n4543 G.n4542 0.686
R5158 G.n4545 G.n4544 0.686
R5159 G.n4547 G.n4546 0.686
R5160 G.n4549 G.n4548 0.686
R5161 G.n4551 G.n4550 0.686
R5162 G.n4553 G.n4552 0.686
R5163 G.n4555 G.n4554 0.686
R5164 G.n2879 G.n2878 0.686
R5165 G.n2877 G.n2876 0.686
R5166 G.n2875 G.n2874 0.686
R5167 G.n2873 G.n2872 0.686
R5168 G.n2871 G.n2870 0.686
R5169 G.n2869 G.n2868 0.686
R5170 G.n2867 G.n2866 0.686
R5171 G.n2865 G.n2864 0.686
R5172 G.n2863 G.n2862 0.686
R5173 G.n2861 G.n2860 0.686
R5174 G.n2859 G.n2858 0.686
R5175 G.n2857 G.n2856 0.686
R5176 G.n2855 G.n2854 0.686
R5177 G.n1620 G.n1619 0.686
R5178 G.n1537 G.n1536 0.686
R5179 G.n1450 G.n1449 0.686
R5180 G.n1362 G.n1361 0.686
R5181 G.n1274 G.n1273 0.686
R5182 G.n1186 G.n1185 0.686
R5183 G.n1098 G.n1097 0.686
R5184 G.n1010 G.n1009 0.686
R5185 G.n925 G.n924 0.686
R5186 G.n4442 G.n4441 0.686
R5187 G.n4444 G.n4443 0.686
R5188 G.n4446 G.n4445 0.686
R5189 G.n4448 G.n4447 0.686
R5190 G.n4450 G.n4449 0.686
R5191 G.n4452 G.n4451 0.686
R5192 G.n4454 G.n4453 0.686
R5193 G.n4456 G.n4455 0.686
R5194 G.n4458 G.n4457 0.686
R5195 G.n4460 G.n4459 0.686
R5196 G.n4462 G.n4461 0.686
R5197 G.n4464 G.n4463 0.686
R5198 G.n4466 G.n4465 0.686
R5199 G.n4468 G.n4467 0.686
R5200 G.n4470 G.n4469 0.686
R5201 G.n4472 G.n4471 0.686
R5202 G.n4474 G.n4473 0.686
R5203 G.n4476 G.n4475 0.686
R5204 G.n4478 G.n4477 0.686
R5205 G.n4480 G.n4479 0.686
R5206 G.n4482 G.n4481 0.686
R5207 G.n4484 G.n4483 0.686
R5208 G.n4486 G.n4485 0.686
R5209 G.n2837 G.n2836 0.686
R5210 G.n2835 G.n2834 0.686
R5211 G.n2833 G.n2832 0.686
R5212 G.n2831 G.n2830 0.686
R5213 G.n2829 G.n2828 0.686
R5214 G.n2827 G.n2826 0.686
R5215 G.n2825 G.n2824 0.686
R5216 G.n2823 G.n2822 0.686
R5217 G.n2821 G.n2820 0.686
R5218 G.n2819 G.n2818 0.686
R5219 G.n2817 G.n2816 0.686
R5220 G.n2815 G.n2814 0.686
R5221 G.n2813 G.n2812 0.686
R5222 G.n4375 G.n4374 0.686
R5223 G.n4377 G.n4376 0.686
R5224 G.n4379 G.n4378 0.686
R5225 G.n4381 G.n4380 0.686
R5226 G.n4383 G.n4382 0.686
R5227 G.n4385 G.n4384 0.686
R5228 G.n4387 G.n4386 0.686
R5229 G.n4389 G.n4388 0.686
R5230 G.n4391 G.n4390 0.686
R5231 G.n4393 G.n4392 0.686
R5232 G.n4395 G.n4394 0.686
R5233 G.n4397 G.n4396 0.686
R5234 G.n4399 G.n4398 0.686
R5235 G.n4401 G.n4400 0.686
R5236 G.n4403 G.n4402 0.686
R5237 G.n4405 G.n4404 0.686
R5238 G.n4407 G.n4406 0.686
R5239 G.n4409 G.n4408 0.686
R5240 G.n4411 G.n4410 0.686
R5241 G.n4413 G.n4412 0.686
R5242 G.n4415 G.n4414 0.686
R5243 G.n2794 G.n2793 0.686
R5244 G.n2792 G.n2791 0.686
R5245 G.n2790 G.n2789 0.686
R5246 G.n2788 G.n2787 0.686
R5247 G.n2786 G.n2785 0.686
R5248 G.n2784 G.n2783 0.686
R5249 G.n2782 G.n2781 0.686
R5250 G.n2780 G.n2779 0.686
R5251 G.n2778 G.n2777 0.686
R5252 G.n2776 G.n2775 0.686
R5253 G.n2774 G.n2773 0.686
R5254 G.n2772 G.n2771 0.686
R5255 G.n1704 G.n1703 0.686
R5256 G.n1626 G.n1625 0.686
R5257 G.n1543 G.n1542 0.686
R5258 G.n1456 G.n1455 0.686
R5259 G.n1368 G.n1367 0.686
R5260 G.n1280 G.n1279 0.686
R5261 G.n1192 G.n1191 0.686
R5262 G.n1104 G.n1103 0.686
R5263 G.n1016 G.n1015 0.686
R5264 G.n931 G.n930 0.686
R5265 G.n849 G.n848 0.686
R5266 G.n773 G.n772 0.686
R5267 G.n4309 G.n4308 0.686
R5268 G.n4311 G.n4310 0.686
R5269 G.n4313 G.n4312 0.686
R5270 G.n4315 G.n4314 0.686
R5271 G.n4317 G.n4316 0.686
R5272 G.n4319 G.n4318 0.686
R5273 G.n4321 G.n4320 0.686
R5274 G.n4323 G.n4322 0.686
R5275 G.n4325 G.n4324 0.686
R5276 G.n4327 G.n4326 0.686
R5277 G.n4329 G.n4328 0.686
R5278 G.n4331 G.n4330 0.686
R5279 G.n4333 G.n4332 0.686
R5280 G.n4335 G.n4334 0.686
R5281 G.n4337 G.n4336 0.686
R5282 G.n4339 G.n4338 0.686
R5283 G.n4341 G.n4340 0.686
R5284 G.n4343 G.n4342 0.686
R5285 G.n4345 G.n4344 0.686
R5286 G.n4347 G.n4346 0.686
R5287 G.n4349 G.n4348 0.686
R5288 G.n2755 G.n2754 0.686
R5289 G.n2753 G.n2752 0.686
R5290 G.n2751 G.n2750 0.686
R5291 G.n2749 G.n2748 0.686
R5292 G.n2747 G.n2746 0.686
R5293 G.n2745 G.n2744 0.686
R5294 G.n2743 G.n2742 0.686
R5295 G.n2741 G.n2740 0.686
R5296 G.n2739 G.n2738 0.686
R5297 G.n2737 G.n2736 0.686
R5298 G.n2735 G.n2734 0.686
R5299 G.n2733 G.n2732 0.686
R5300 G.n4248 G.n4247 0.686
R5301 G.n4250 G.n4249 0.686
R5302 G.n4252 G.n4251 0.686
R5303 G.n4254 G.n4253 0.686
R5304 G.n4256 G.n4255 0.686
R5305 G.n4258 G.n4257 0.686
R5306 G.n4260 G.n4259 0.686
R5307 G.n4262 G.n4261 0.686
R5308 G.n4264 G.n4263 0.686
R5309 G.n4266 G.n4265 0.686
R5310 G.n4268 G.n4267 0.686
R5311 G.n4270 G.n4269 0.686
R5312 G.n4272 G.n4271 0.686
R5313 G.n4274 G.n4273 0.686
R5314 G.n4276 G.n4275 0.686
R5315 G.n4278 G.n4277 0.686
R5316 G.n4280 G.n4279 0.686
R5317 G.n4282 G.n4281 0.686
R5318 G.n4284 G.n4283 0.686
R5319 G.n2717 G.n2716 0.686
R5320 G.n2715 G.n2714 0.686
R5321 G.n2713 G.n2712 0.686
R5322 G.n2711 G.n2710 0.686
R5323 G.n2709 G.n2708 0.686
R5324 G.n2707 G.n2706 0.686
R5325 G.n2705 G.n2704 0.686
R5326 G.n2703 G.n2702 0.686
R5327 G.n2701 G.n2700 0.686
R5328 G.n2699 G.n2698 0.686
R5329 G.n2697 G.n2696 0.686
R5330 G.n1782 G.n1781 0.686
R5331 G.n1710 G.n1709 0.686
R5332 G.n1632 G.n1631 0.686
R5333 G.n1549 G.n1548 0.686
R5334 G.n1462 G.n1461 0.686
R5335 G.n1374 G.n1373 0.686
R5336 G.n1286 G.n1285 0.686
R5337 G.n1198 G.n1197 0.686
R5338 G.n1110 G.n1109 0.686
R5339 G.n1022 G.n1021 0.686
R5340 G.n937 G.n936 0.686
R5341 G.n855 G.n854 0.686
R5342 G.n779 G.n778 0.686
R5343 G.n706 G.n705 0.686
R5344 G.n636 G.n635 0.686
R5345 G.n4188 G.n4187 0.686
R5346 G.n4190 G.n4189 0.686
R5347 G.n4192 G.n4191 0.686
R5348 G.n4194 G.n4193 0.686
R5349 G.n4196 G.n4195 0.686
R5350 G.n4198 G.n4197 0.686
R5351 G.n4200 G.n4199 0.686
R5352 G.n4202 G.n4201 0.686
R5353 G.n4204 G.n4203 0.686
R5354 G.n4206 G.n4205 0.686
R5355 G.n4208 G.n4207 0.686
R5356 G.n4210 G.n4209 0.686
R5357 G.n4212 G.n4211 0.686
R5358 G.n4214 G.n4213 0.686
R5359 G.n4216 G.n4215 0.686
R5360 G.n4218 G.n4217 0.686
R5361 G.n4220 G.n4219 0.686
R5362 G.n4222 G.n4221 0.686
R5363 G.n4224 G.n4223 0.686
R5364 G.n2681 G.n2680 0.686
R5365 G.n2679 G.n2678 0.686
R5366 G.n2677 G.n2676 0.686
R5367 G.n2675 G.n2674 0.686
R5368 G.n2673 G.n2672 0.686
R5369 G.n2671 G.n2670 0.686
R5370 G.n2669 G.n2668 0.686
R5371 G.n2667 G.n2666 0.686
R5372 G.n2665 G.n2664 0.686
R5373 G.n2663 G.n2662 0.686
R5374 G.n2661 G.n2660 0.686
R5375 G.n4133 G.n4132 0.686
R5376 G.n4135 G.n4134 0.686
R5377 G.n4137 G.n4136 0.686
R5378 G.n4139 G.n4138 0.686
R5379 G.n4141 G.n4140 0.686
R5380 G.n4143 G.n4142 0.686
R5381 G.n4145 G.n4144 0.686
R5382 G.n4147 G.n4146 0.686
R5383 G.n4149 G.n4148 0.686
R5384 G.n4151 G.n4150 0.686
R5385 G.n4153 G.n4152 0.686
R5386 G.n4155 G.n4154 0.686
R5387 G.n4157 G.n4156 0.686
R5388 G.n4159 G.n4158 0.686
R5389 G.n4161 G.n4160 0.686
R5390 G.n4163 G.n4162 0.686
R5391 G.n4165 G.n4164 0.686
R5392 G.n2646 G.n2645 0.686
R5393 G.n2644 G.n2643 0.686
R5394 G.n2642 G.n2641 0.686
R5395 G.n2640 G.n2639 0.686
R5396 G.n2638 G.n2637 0.686
R5397 G.n2636 G.n2635 0.686
R5398 G.n2634 G.n2633 0.686
R5399 G.n2632 G.n2631 0.686
R5400 G.n2630 G.n2629 0.686
R5401 G.n2628 G.n2627 0.686
R5402 G.n1856 G.n1855 0.686
R5403 G.n1788 G.n1787 0.686
R5404 G.n1716 G.n1715 0.686
R5405 G.n1638 G.n1637 0.686
R5406 G.n1555 G.n1554 0.686
R5407 G.n1468 G.n1467 0.686
R5408 G.n1380 G.n1379 0.686
R5409 G.n1292 G.n1291 0.686
R5410 G.n1204 G.n1203 0.686
R5411 G.n1116 G.n1115 0.686
R5412 G.n1028 G.n1027 0.686
R5413 G.n943 G.n942 0.686
R5414 G.n861 G.n860 0.686
R5415 G.n785 G.n784 0.686
R5416 G.n712 G.n711 0.686
R5417 G.n642 G.n641 0.686
R5418 G.n575 G.n574 0.686
R5419 G.n511 G.n510 0.686
R5420 G.n4079 G.n4078 0.686
R5421 G.n4081 G.n4080 0.686
R5422 G.n4083 G.n4082 0.686
R5423 G.n4085 G.n4084 0.686
R5424 G.n4087 G.n4086 0.686
R5425 G.n4089 G.n4088 0.686
R5426 G.n4091 G.n4090 0.686
R5427 G.n4093 G.n4092 0.686
R5428 G.n4095 G.n4094 0.686
R5429 G.n4097 G.n4096 0.686
R5430 G.n4099 G.n4098 0.686
R5431 G.n4101 G.n4100 0.686
R5432 G.n4103 G.n4102 0.686
R5433 G.n4105 G.n4104 0.686
R5434 G.n4107 G.n4106 0.686
R5435 G.n4109 G.n4108 0.686
R5436 G.n4111 G.n4110 0.686
R5437 G.n2613 G.n2612 0.686
R5438 G.n2611 G.n2610 0.686
R5439 G.n2609 G.n2608 0.686
R5440 G.n2607 G.n2606 0.686
R5441 G.n2605 G.n2604 0.686
R5442 G.n2603 G.n2602 0.686
R5443 G.n2601 G.n2600 0.686
R5444 G.n2599 G.n2598 0.686
R5445 G.n2597 G.n2596 0.686
R5446 G.n2595 G.n2594 0.686
R5447 G.n4030 G.n4029 0.686
R5448 G.n4032 G.n4031 0.686
R5449 G.n4034 G.n4033 0.686
R5450 G.n4036 G.n4035 0.686
R5451 G.n4038 G.n4037 0.686
R5452 G.n4040 G.n4039 0.686
R5453 G.n4042 G.n4041 0.686
R5454 G.n4044 G.n4043 0.686
R5455 G.n4046 G.n4045 0.686
R5456 G.n4048 G.n4047 0.686
R5457 G.n4050 G.n4049 0.686
R5458 G.n4052 G.n4051 0.686
R5459 G.n4054 G.n4053 0.686
R5460 G.n4056 G.n4055 0.686
R5461 G.n4058 G.n4057 0.686
R5462 G.n2581 G.n2580 0.686
R5463 G.n2579 G.n2578 0.686
R5464 G.n2577 G.n2576 0.686
R5465 G.n2575 G.n2574 0.686
R5466 G.n2573 G.n2572 0.686
R5467 G.n2571 G.n2570 0.686
R5468 G.n2569 G.n2568 0.686
R5469 G.n2567 G.n2566 0.686
R5470 G.n2565 G.n2564 0.686
R5471 G.n1981 G.n1980 0.686
R5472 G.n1924 G.n1923 0.686
R5473 G.n1862 G.n1861 0.686
R5474 G.n1794 G.n1793 0.686
R5475 G.n1722 G.n1721 0.686
R5476 G.n1644 G.n1643 0.686
R5477 G.n1561 G.n1560 0.686
R5478 G.n1474 G.n1473 0.686
R5479 G.n1386 G.n1385 0.686
R5480 G.n1298 G.n1297 0.686
R5481 G.n1210 G.n1209 0.686
R5482 G.n1122 G.n1121 0.686
R5483 G.n1034 G.n1033 0.686
R5484 G.n949 G.n948 0.686
R5485 G.n867 G.n866 0.686
R5486 G.n791 G.n790 0.686
R5487 G.n718 G.n717 0.686
R5488 G.n648 G.n647 0.686
R5489 G.n581 G.n580 0.686
R5490 G.n517 G.n516 0.686
R5491 G.n456 G.n455 0.686
R5492 G.n398 G.n397 0.686
R5493 G.n3982 G.n3981 0.686
R5494 G.n3984 G.n3983 0.686
R5495 G.n3986 G.n3985 0.686
R5496 G.n3988 G.n3987 0.686
R5497 G.n3990 G.n3989 0.686
R5498 G.n3992 G.n3991 0.686
R5499 G.n3994 G.n3993 0.686
R5500 G.n3996 G.n3995 0.686
R5501 G.n3998 G.n3997 0.686
R5502 G.n4000 G.n3999 0.686
R5503 G.n4002 G.n4001 0.686
R5504 G.n4004 G.n4003 0.686
R5505 G.n4006 G.n4005 0.686
R5506 G.n4008 G.n4007 0.686
R5507 G.n4010 G.n4009 0.686
R5508 G.n2552 G.n2551 0.686
R5509 G.n2550 G.n2549 0.686
R5510 G.n2548 G.n2547 0.686
R5511 G.n2546 G.n2545 0.686
R5512 G.n2544 G.n2543 0.686
R5513 G.n2542 G.n2541 0.686
R5514 G.n2540 G.n2539 0.686
R5515 G.n2538 G.n2537 0.686
R5516 G.n2536 G.n2535 0.686
R5517 G.n3937 G.n3936 0.686
R5518 G.n3939 G.n3938 0.686
R5519 G.n3941 G.n3940 0.686
R5520 G.n3943 G.n3942 0.686
R5521 G.n3945 G.n3944 0.686
R5522 G.n3947 G.n3946 0.686
R5523 G.n3949 G.n3948 0.686
R5524 G.n3951 G.n3950 0.686
R5525 G.n3953 G.n3952 0.686
R5526 G.n3955 G.n3954 0.686
R5527 G.n3957 G.n3956 0.686
R5528 G.n3959 G.n3958 0.686
R5529 G.n3961 G.n3960 0.686
R5530 G.n3963 G.n3962 0.686
R5531 G.n2523 G.n2522 0.686
R5532 G.n2521 G.n2520 0.686
R5533 G.n2519 G.n2518 0.686
R5534 G.n2517 G.n2516 0.686
R5535 G.n2515 G.n2514 0.686
R5536 G.n2513 G.n2512 0.686
R5537 G.n2511 G.n2510 0.686
R5538 G.n2509 G.n2508 0.686
R5539 G.n2038 G.n2037 0.686
R5540 G.n1987 G.n1986 0.686
R5541 G.n1930 G.n1929 0.686
R5542 G.n1868 G.n1867 0.686
R5543 G.n1800 G.n1799 0.686
R5544 G.n1728 G.n1727 0.686
R5545 G.n1650 G.n1649 0.686
R5546 G.n1567 G.n1566 0.686
R5547 G.n1480 G.n1479 0.686
R5548 G.n1392 G.n1391 0.686
R5549 G.n1304 G.n1303 0.686
R5550 G.n1216 G.n1215 0.686
R5551 G.n1128 G.n1127 0.686
R5552 G.n1040 G.n1039 0.686
R5553 G.n955 G.n954 0.686
R5554 G.n873 G.n872 0.686
R5555 G.n797 G.n796 0.686
R5556 G.n724 G.n723 0.686
R5557 G.n654 G.n653 0.686
R5558 G.n587 G.n586 0.686
R5559 G.n523 G.n522 0.686
R5560 G.n462 G.n461 0.686
R5561 G.n404 G.n403 0.686
R5562 G.n349 G.n348 0.686
R5563 G.n3892 G.n3891 0.686
R5564 G.n3894 G.n3893 0.686
R5565 G.n3896 G.n3895 0.686
R5566 G.n3898 G.n3897 0.686
R5567 G.n3900 G.n3899 0.686
R5568 G.n3902 G.n3901 0.686
R5569 G.n3904 G.n3903 0.686
R5570 G.n3906 G.n3905 0.686
R5571 G.n3908 G.n3907 0.686
R5572 G.n3910 G.n3909 0.686
R5573 G.n3912 G.n3911 0.686
R5574 G.n3914 G.n3913 0.686
R5575 G.n3916 G.n3915 0.686
R5576 G.n3918 G.n3917 0.686
R5577 G.n2497 G.n2496 0.686
R5578 G.n2495 G.n2494 0.686
R5579 G.n2493 G.n2492 0.686
R5580 G.n2491 G.n2490 0.686
R5581 G.n2489 G.n2488 0.686
R5582 G.n2487 G.n2486 0.686
R5583 G.n2485 G.n2484 0.686
R5584 G.n2483 G.n2482 0.686
R5585 G.n3852 G.n3851 0.686
R5586 G.n3854 G.n3853 0.686
R5587 G.n3856 G.n3855 0.686
R5588 G.n3858 G.n3857 0.686
R5589 G.n3860 G.n3859 0.686
R5590 G.n3862 G.n3861 0.686
R5591 G.n3864 G.n3863 0.686
R5592 G.n3866 G.n3865 0.686
R5593 G.n3868 G.n3867 0.686
R5594 G.n3870 G.n3869 0.686
R5595 G.n3872 G.n3871 0.686
R5596 G.n3874 G.n3873 0.686
R5597 G.n2471 G.n2470 0.686
R5598 G.n2469 G.n2468 0.686
R5599 G.n2467 G.n2466 0.686
R5600 G.n2465 G.n2464 0.686
R5601 G.n2463 G.n2462 0.686
R5602 G.n2461 G.n2460 0.686
R5603 G.n2089 G.n2088 0.686
R5604 G.n2044 G.n2043 0.686
R5605 G.n1993 G.n1992 0.686
R5606 G.n1936 G.n1935 0.686
R5607 G.n1874 G.n1873 0.686
R5608 G.n1806 G.n1805 0.686
R5609 G.n1734 G.n1733 0.686
R5610 G.n1656 G.n1655 0.686
R5611 G.n1573 G.n1572 0.686
R5612 G.n1486 G.n1485 0.686
R5613 G.n1398 G.n1397 0.686
R5614 G.n1310 G.n1309 0.686
R5615 G.n1222 G.n1221 0.686
R5616 G.n1134 G.n1133 0.686
R5617 G.n1046 G.n1045 0.686
R5618 G.n961 G.n960 0.686
R5619 G.n879 G.n878 0.686
R5620 G.n803 G.n802 0.686
R5621 G.n730 G.n729 0.686
R5622 G.n660 G.n659 0.686
R5623 G.n593 G.n592 0.686
R5624 G.n529 G.n528 0.686
R5625 G.n468 G.n467 0.686
R5626 G.n410 G.n409 0.686
R5627 G.n355 G.n354 0.686
R5628 G.n306 G.n305 0.686
R5629 G.n260 G.n259 0.686
R5630 G.n3813 G.n3812 0.686
R5631 G.n3815 G.n3814 0.686
R5632 G.n3817 G.n3816 0.686
R5633 G.n3819 G.n3818 0.686
R5634 G.n3821 G.n3820 0.686
R5635 G.n3823 G.n3822 0.686
R5636 G.n3825 G.n3824 0.686
R5637 G.n3827 G.n3826 0.686
R5638 G.n3829 G.n3828 0.686
R5639 G.n3831 G.n3830 0.686
R5640 G.n3833 G.n3832 0.686
R5641 G.n3835 G.n3834 0.686
R5642 G.n2450 G.n2449 0.686
R5643 G.n2448 G.n2447 0.686
R5644 G.n2446 G.n2445 0.686
R5645 G.n2444 G.n2443 0.686
R5646 G.n2442 G.n2441 0.686
R5647 G.n2440 G.n2439 0.686
R5648 G.n2438 G.n2437 0.686
R5649 G.n3779 G.n3778 0.686
R5650 G.n3781 G.n3780 0.686
R5651 G.n3783 G.n3782 0.686
R5652 G.n3785 G.n3784 0.686
R5653 G.n3787 G.n3786 0.686
R5654 G.n3789 G.n3788 0.686
R5655 G.n3791 G.n3790 0.686
R5656 G.n3793 G.n3792 0.686
R5657 G.n3795 G.n3794 0.686
R5658 G.n3797 G.n3796 0.686
R5659 G.n2427 G.n2426 0.686
R5660 G.n2425 G.n2424 0.686
R5661 G.n2423 G.n2422 0.686
R5662 G.n2421 G.n2420 0.686
R5663 G.n2419 G.n2418 0.686
R5664 G.n2136 G.n2135 0.686
R5665 G.n2095 G.n2094 0.686
R5666 G.n2050 G.n2049 0.686
R5667 G.n1999 G.n1998 0.686
R5668 G.n1942 G.n1941 0.686
R5669 G.n1880 G.n1879 0.686
R5670 G.n1812 G.n1811 0.686
R5671 G.n1740 G.n1739 0.686
R5672 G.n1662 G.n1661 0.686
R5673 G.n1579 G.n1578 0.686
R5674 G.n1492 G.n1491 0.686
R5675 G.n1404 G.n1403 0.686
R5676 G.n1316 G.n1315 0.686
R5677 G.n1228 G.n1227 0.686
R5678 G.n1140 G.n1139 0.686
R5679 G.n1052 G.n1051 0.686
R5680 G.n967 G.n966 0.686
R5681 G.n885 G.n884 0.686
R5682 G.n809 G.n808 0.686
R5683 G.n736 G.n735 0.686
R5684 G.n666 G.n665 0.686
R5685 G.n599 G.n598 0.686
R5686 G.n535 G.n534 0.686
R5687 G.n474 G.n473 0.686
R5688 G.n416 G.n415 0.686
R5689 G.n361 G.n360 0.686
R5690 G.n312 G.n311 0.686
R5691 G.n266 G.n265 0.686
R5692 G.n223 G.n222 0.686
R5693 G.n183 G.n182 0.686
R5694 G.n3746 G.n3745 0.686
R5695 G.n3748 G.n3747 0.686
R5696 G.n3750 G.n3749 0.686
R5697 G.n3752 G.n3751 0.686
R5698 G.n3754 G.n3753 0.686
R5699 G.n3756 G.n3755 0.686
R5700 G.n3758 G.n3757 0.686
R5701 G.n3760 G.n3759 0.686
R5702 G.n3762 G.n3761 0.686
R5703 G.n3764 G.n3763 0.686
R5704 G.n2409 G.n2408 0.686
R5705 G.n2407 G.n2406 0.686
R5706 G.n2405 G.n2404 0.686
R5707 G.n2403 G.n2402 0.686
R5708 G.n2401 G.n2400 0.686
R5709 G.n2399 G.n2398 0.686
R5710 G.n3718 G.n3717 0.686
R5711 G.n3720 G.n3719 0.686
R5712 G.n3722 G.n3721 0.686
R5713 G.n3724 G.n3723 0.686
R5714 G.n3726 G.n3725 0.686
R5715 G.n3728 G.n3727 0.686
R5716 G.n3730 G.n3729 0.686
R5717 G.n3732 G.n3731 0.686
R5718 G.n2389 G.n2388 0.686
R5719 G.n2387 G.n2386 0.686
R5720 G.n2385 G.n2384 0.686
R5721 G.n2383 G.n2382 0.686
R5722 G.n2177 G.n2176 0.686
R5723 G.n2142 G.n2141 0.686
R5724 G.n2101 G.n2100 0.686
R5725 G.n2056 G.n2055 0.686
R5726 G.n2005 G.n2004 0.686
R5727 G.n1948 G.n1947 0.686
R5728 G.n1886 G.n1885 0.686
R5729 G.n1818 G.n1817 0.686
R5730 G.n1746 G.n1745 0.686
R5731 G.n1668 G.n1667 0.686
R5732 G.n1585 G.n1584 0.686
R5733 G.n1498 G.n1497 0.686
R5734 G.n1410 G.n1409 0.686
R5735 G.n1322 G.n1321 0.686
R5736 G.n1234 G.n1233 0.686
R5737 G.n1146 G.n1145 0.686
R5738 G.n1058 G.n1057 0.686
R5739 G.n973 G.n972 0.686
R5740 G.n891 G.n890 0.686
R5741 G.n815 G.n814 0.686
R5742 G.n742 G.n741 0.686
R5743 G.n672 G.n671 0.686
R5744 G.n605 G.n604 0.686
R5745 G.n541 G.n540 0.686
R5746 G.n480 G.n479 0.686
R5747 G.n422 G.n421 0.686
R5748 G.n367 G.n366 0.686
R5749 G.n318 G.n317 0.686
R5750 G.n272 G.n271 0.686
R5751 G.n229 G.n228 0.686
R5752 G.n189 G.n188 0.686
R5753 G.n152 G.n151 0.686
R5754 G.n118 G.n117 0.686
R5755 G.n3691 G.n3690 0.686
R5756 G.n3693 G.n3692 0.686
R5757 G.n3695 G.n3694 0.686
R5758 G.n3697 G.n3696 0.686
R5759 G.n3699 G.n3698 0.686
R5760 G.n3701 G.n3700 0.686
R5761 G.n3703 G.n3702 0.686
R5762 G.n3705 G.n3704 0.686
R5763 G.n2374 G.n2373 0.686
R5764 G.n2372 G.n2371 0.686
R5765 G.n2370 G.n2369 0.686
R5766 G.n2368 G.n2367 0.686
R5767 G.n3667 G.n3666 0.686
R5768 G.n3669 G.n3668 0.686
R5769 G.n3671 G.n3670 0.686
R5770 G.n3673 G.n3672 0.686
R5771 G.n3675 G.n3674 0.686
R5772 G.n3677 G.n3676 0.686
R5773 G.n3679 G.n3678 0.686
R5774 G.n2358 G.n2357 0.686
R5775 G.n2356 G.n2355 0.686
R5776 G.n2354 G.n2353 0.686
R5777 G.n2213 G.n2212 0.686
R5778 G.n2183 G.n2182 0.686
R5779 G.n2148 G.n2147 0.686
R5780 G.n2107 G.n2106 0.686
R5781 G.n2062 G.n2061 0.686
R5782 G.n2011 G.n2010 0.686
R5783 G.n1954 G.n1953 0.686
R5784 G.n1892 G.n1891 0.686
R5785 G.n1824 G.n1823 0.686
R5786 G.n1752 G.n1751 0.686
R5787 G.n1674 G.n1673 0.686
R5788 G.n1591 G.n1590 0.686
R5789 G.n1504 G.n1503 0.686
R5790 G.n1416 G.n1415 0.686
R5791 G.n1328 G.n1327 0.686
R5792 G.n1240 G.n1239 0.686
R5793 G.n1152 G.n1151 0.686
R5794 G.n1064 G.n1063 0.686
R5795 G.n979 G.n978 0.686
R5796 G.n897 G.n896 0.686
R5797 G.n821 G.n820 0.686
R5798 G.n748 G.n747 0.686
R5799 G.n678 G.n677 0.686
R5800 G.n611 G.n610 0.686
R5801 G.n547 G.n546 0.686
R5802 G.n486 G.n485 0.686
R5803 G.n428 G.n427 0.686
R5804 G.n373 G.n372 0.686
R5805 G.n324 G.n323 0.686
R5806 G.n278 G.n277 0.686
R5807 G.n235 G.n234 0.686
R5808 G.n195 G.n194 0.686
R5809 G.n158 G.n157 0.686
R5810 G.n124 G.n123 0.686
R5811 G.n93 G.n92 0.686
R5812 G.n3643 G.n3642 0.686
R5813 G.n3645 G.n3644 0.686
R5814 G.n3647 G.n3646 0.686
R5815 G.n3649 G.n3648 0.686
R5816 G.n3651 G.n3650 0.686
R5817 G.n3653 G.n3652 0.686
R5818 G.n3655 G.n3654 0.686
R5819 G.n2346 G.n2345 0.686
R5820 G.n2344 G.n2343 0.686
R5821 G.n2342 G.n2341 0.686
R5822 G.n3624 G.n3623 0.686
R5823 G.n3626 G.n3625 0.686
R5824 G.n3628 G.n3627 0.686
R5825 G.n3630 G.n3629 0.686
R5826 G.n3632 G.n3631 0.686
R5827 G.n2335 G.n2334 0.686
R5828 G.n2333 G.n2332 0.686
R5829 G.n2243 G.n2242 0.686
R5830 G.n2219 G.n2218 0.686
R5831 G.n2189 G.n2188 0.686
R5832 G.n2154 G.n2153 0.686
R5833 G.n2113 G.n2112 0.686
R5834 G.n2068 G.n2067 0.686
R5835 G.n2017 G.n2016 0.686
R5836 G.n1960 G.n1959 0.686
R5837 G.n1898 G.n1897 0.686
R5838 G.n1830 G.n1829 0.686
R5839 G.n1758 G.n1757 0.686
R5840 G.n1680 G.n1679 0.686
R5841 G.n1597 G.n1596 0.686
R5842 G.n1510 G.n1509 0.686
R5843 G.n1422 G.n1421 0.686
R5844 G.n1334 G.n1333 0.686
R5845 G.n1246 G.n1245 0.686
R5846 G.n1158 G.n1157 0.686
R5847 G.n1070 G.n1069 0.686
R5848 G.n985 G.n984 0.686
R5849 G.n903 G.n902 0.686
R5850 G.n827 G.n826 0.686
R5851 G.n754 G.n753 0.686
R5852 G.n684 G.n683 0.686
R5853 G.n617 G.n616 0.686
R5854 G.n553 G.n552 0.686
R5855 G.n492 G.n491 0.686
R5856 G.n434 G.n433 0.686
R5857 G.n379 G.n378 0.686
R5858 G.n330 G.n329 0.686
R5859 G.n284 G.n283 0.686
R5860 G.n241 G.n240 0.686
R5861 G.n201 G.n200 0.686
R5862 G.n164 G.n163 0.686
R5863 G.n130 G.n129 0.686
R5864 G.n99 G.n98 0.686
R5865 G.n74 G.n73 0.686
R5866 G.n52 G.n51 0.686
R5867 G.n3606 G.n3605 0.686
R5868 G.n3608 G.n3607 0.686
R5869 G.n3610 G.n3609 0.686
R5870 G.n3612 G.n3611 0.686
R5871 G.n3614 G.n3613 0.686
R5872 G.n2326 G.n2325 0.686
R5873 G.n2324 G.n2323 0.686
R5874 G.n3593 G.n3592 0.686
R5875 G.n3595 G.n3594 0.686
R5876 G.n3597 G.n3596 0.686
R5877 G.n2318 G.n2317 0.686
R5878 G.n2269 G.n2268 0.686
R5879 G.n2249 G.n2248 0.686
R5880 G.n2225 G.n2224 0.686
R5881 G.n2195 G.n2194 0.686
R5882 G.n2160 G.n2159 0.686
R5883 G.n2119 G.n2118 0.686
R5884 G.n2074 G.n2073 0.686
R5885 G.n2023 G.n2022 0.686
R5886 G.n1966 G.n1965 0.686
R5887 G.n1904 G.n1903 0.686
R5888 G.n1836 G.n1835 0.686
R5889 G.n1764 G.n1763 0.686
R5890 G.n1686 G.n1685 0.686
R5891 G.n1603 G.n1602 0.686
R5892 G.n1516 G.n1515 0.686
R5893 G.n1428 G.n1427 0.686
R5894 G.n1340 G.n1339 0.686
R5895 G.n1252 G.n1251 0.686
R5896 G.n1164 G.n1163 0.686
R5897 G.n1076 G.n1075 0.686
R5898 G.n991 G.n990 0.686
R5899 G.n909 G.n908 0.686
R5900 G.n833 G.n832 0.686
R5901 G.n760 G.n759 0.686
R5902 G.n690 G.n689 0.686
R5903 G.n623 G.n622 0.686
R5904 G.n559 G.n558 0.686
R5905 G.n498 G.n497 0.686
R5906 G.n440 G.n439 0.686
R5907 G.n385 G.n384 0.686
R5908 G.n336 G.n335 0.686
R5909 G.n290 G.n289 0.686
R5910 G.n247 G.n246 0.686
R5911 G.n207 G.n206 0.686
R5912 G.n170 G.n169 0.686
R5913 G.n136 G.n135 0.686
R5914 G.n105 G.n104 0.686
R5915 G.n80 G.n79 0.686
R5916 G.n58 G.n57 0.686
R5917 G.n39 G.n38 0.686
R5918 G.n23 G.n22 0.686
R5919 G.n3581 G.n3580 0.686
R5920 G.n3583 G.n3582 0.686
R5921 G.n3585 G.n3584 0.686
R5922 G.n2312 G.n2311 0.686
R5923 G.n3574 G.n3573 0.686
R5924 G.n2298 G.n2297 0.686
R5925 G.n2289 G.n2288 0.686
R5926 G.n2275 G.n2274 0.686
R5927 G.n2255 G.n2254 0.686
R5928 G.n2231 G.n2230 0.686
R5929 G.n2201 G.n2200 0.686
R5930 G.n2166 G.n2165 0.686
R5931 G.n2125 G.n2124 0.686
R5932 G.n2080 G.n2079 0.686
R5933 G.n2029 G.n2028 0.686
R5934 G.n1972 G.n1971 0.686
R5935 G.n1910 G.n1909 0.686
R5936 G.n1842 G.n1841 0.686
R5937 G.n1770 G.n1769 0.686
R5938 G.n1692 G.n1691 0.686
R5939 G.n1609 G.n1608 0.686
R5940 G.n1522 G.n1521 0.686
R5941 G.n1434 G.n1433 0.686
R5942 G.n1346 G.n1345 0.686
R5943 G.n1258 G.n1257 0.686
R5944 G.n1170 G.n1169 0.686
R5945 G.n1082 G.n1081 0.686
R5946 G.n997 G.n996 0.686
R5947 G.n915 G.n914 0.686
R5948 G.n839 G.n838 0.686
R5949 G.n766 G.n765 0.686
R5950 G.n696 G.n695 0.686
R5951 G.n629 G.n628 0.686
R5952 G.n565 G.n564 0.686
R5953 G.n504 G.n503 0.686
R5954 G.n446 G.n445 0.686
R5955 G.n391 G.n390 0.686
R5956 G.n342 G.n341 0.686
R5957 G.n296 G.n295 0.686
R5958 G.n253 G.n252 0.686
R5959 G.n213 G.n212 0.686
R5960 G.n176 G.n175 0.686
R5961 G.n142 G.n141 0.686
R5962 G.n111 G.n110 0.686
R5963 G.n86 G.n85 0.686
R5964 G.n64 G.n63 0.686
R5965 G.n45 G.n44 0.686
R5966 G.n29 G.n28 0.686
R5967 G.n16 G.n15 0.686
R5968 G.n6 G.n5 0.686
R5969 G.n3568 G.n3567 0.686
R5970 G.n2301 G.n2300 0.686
R5971 G.n2292 G.n2291 0.686
R5972 G.n2278 G.n2277 0.686
R5973 G.n2258 G.n2257 0.686
R5974 G.n2234 G.n2233 0.686
R5975 G.n2204 G.n2203 0.686
R5976 G.n2169 G.n2168 0.686
R5977 G.n2128 G.n2127 0.686
R5978 G.n2083 G.n2082 0.686
R5979 G.n2032 G.n2031 0.686
R5980 G.n1975 G.n1974 0.686
R5981 G.n1913 G.n1912 0.686
R5982 G.n1845 G.n1844 0.686
R5983 G.n1773 G.n1772 0.686
R5984 G.n1695 G.n1694 0.686
R5985 G.n1612 G.n1611 0.686
R5986 G.n1525 G.n1524 0.686
R5987 G.n1437 G.n1436 0.686
R5988 G.n1349 G.n1348 0.686
R5989 G.n1261 G.n1260 0.686
R5990 G.n1173 G.n1172 0.686
R5991 G.n1085 G.n1084 0.686
R5992 G.n1000 G.n999 0.686
R5993 G.n918 G.n917 0.686
R5994 G.n842 G.n841 0.686
R5995 G.n769 G.n768 0.686
R5996 G.n699 G.n698 0.686
R5997 G.n632 G.n631 0.686
R5998 G.n568 G.n567 0.686
R5999 G.n507 G.n506 0.686
R6000 G.n449 G.n448 0.686
R6001 G.n394 G.n393 0.686
R6002 G.n345 G.n344 0.686
R6003 G.n299 G.n298 0.686
R6004 G.n256 G.n255 0.686
R6005 G.n216 G.n215 0.686
R6006 G.n179 G.n178 0.686
R6007 G.n145 G.n144 0.686
R6008 G.n114 G.n113 0.686
R6009 G.n89 G.n88 0.686
R6010 G.n67 G.n66 0.686
R6011 G.n48 G.n47 0.686
R6012 G.n32 G.n31 0.686
R6013 G.n19 G.n18 0.686
R6014 G.n9 G.n8 0.686
R6015 G.n2 G.n1 0.686
R6016 G.n2286 G.n2285 0.686
R6017 G.n2272 G.n2271 0.686
R6018 G.n2252 G.n2251 0.686
R6019 G.n2228 G.n2227 0.686
R6020 G.n2198 G.n2197 0.686
R6021 G.n2163 G.n2162 0.686
R6022 G.n2122 G.n2121 0.686
R6023 G.n2077 G.n2076 0.686
R6024 G.n2026 G.n2025 0.686
R6025 G.n1969 G.n1968 0.686
R6026 G.n1907 G.n1906 0.686
R6027 G.n1839 G.n1838 0.686
R6028 G.n1767 G.n1766 0.686
R6029 G.n1689 G.n1688 0.686
R6030 G.n1606 G.n1605 0.686
R6031 G.n1519 G.n1518 0.686
R6032 G.n1431 G.n1430 0.686
R6033 G.n1343 G.n1342 0.686
R6034 G.n1255 G.n1254 0.686
R6035 G.n1167 G.n1166 0.686
R6036 G.n1079 G.n1078 0.686
R6037 G.n994 G.n993 0.686
R6038 G.n912 G.n911 0.686
R6039 G.n836 G.n835 0.686
R6040 G.n763 G.n762 0.686
R6041 G.n693 G.n692 0.686
R6042 G.n626 G.n625 0.686
R6043 G.n562 G.n561 0.686
R6044 G.n501 G.n500 0.686
R6045 G.n443 G.n442 0.686
R6046 G.n388 G.n387 0.686
R6047 G.n339 G.n338 0.686
R6048 G.n293 G.n292 0.686
R6049 G.n250 G.n249 0.686
R6050 G.n210 G.n209 0.686
R6051 G.n173 G.n172 0.686
R6052 G.n139 G.n138 0.686
R6053 G.n108 G.n107 0.686
R6054 G.n83 G.n82 0.686
R6055 G.n61 G.n60 0.686
R6056 G.n42 G.n41 0.686
R6057 G.n26 G.n25 0.686
R6058 G.n13 G.n12 0.686
R6059 G.n3573 G.n3572 0.686
R6060 G.n3575 G.n3574 0.686
R6061 G.n3584 G.n3583 0.686
R6062 G.n3582 G.n3581 0.686
R6063 G.n2317 G.n2316 0.686
R6064 G.n2319 G.n2318 0.686
R6065 G.n2325 G.n2324 0.686
R6066 G.n2266 G.n2265 0.686
R6067 G.n2246 G.n2245 0.686
R6068 G.n2222 G.n2221 0.686
R6069 G.n2192 G.n2191 0.686
R6070 G.n2157 G.n2156 0.686
R6071 G.n2116 G.n2115 0.686
R6072 G.n2071 G.n2070 0.686
R6073 G.n2020 G.n2019 0.686
R6074 G.n1963 G.n1962 0.686
R6075 G.n1901 G.n1900 0.686
R6076 G.n1833 G.n1832 0.686
R6077 G.n1761 G.n1760 0.686
R6078 G.n1683 G.n1682 0.686
R6079 G.n1600 G.n1599 0.686
R6080 G.n1513 G.n1512 0.686
R6081 G.n1425 G.n1424 0.686
R6082 G.n1337 G.n1336 0.686
R6083 G.n1249 G.n1248 0.686
R6084 G.n1161 G.n1160 0.686
R6085 G.n1073 G.n1072 0.686
R6086 G.n988 G.n987 0.686
R6087 G.n906 G.n905 0.686
R6088 G.n830 G.n829 0.686
R6089 G.n757 G.n756 0.686
R6090 G.n687 G.n686 0.686
R6091 G.n620 G.n619 0.686
R6092 G.n556 G.n555 0.686
R6093 G.n495 G.n494 0.686
R6094 G.n437 G.n436 0.686
R6095 G.n382 G.n381 0.686
R6096 G.n333 G.n332 0.686
R6097 G.n287 G.n286 0.686
R6098 G.n244 G.n243 0.686
R6099 G.n204 G.n203 0.686
R6100 G.n167 G.n166 0.686
R6101 G.n133 G.n132 0.686
R6102 G.n102 G.n101 0.686
R6103 G.n77 G.n76 0.686
R6104 G.n55 G.n54 0.686
R6105 G.n36 G.n35 0.686
R6106 G.n3592 G.n3591 0.686
R6107 G.n3594 G.n3593 0.686
R6108 G.n3596 G.n3595 0.686
R6109 G.n3598 G.n3597 0.686
R6110 G.n3613 G.n3612 0.686
R6111 G.n3611 G.n3610 0.686
R6112 G.n3609 G.n3608 0.686
R6113 G.n3607 G.n3606 0.686
R6114 G.n2332 G.n2331 0.686
R6115 G.n2334 G.n2333 0.686
R6116 G.n2336 G.n2335 0.686
R6117 G.n2345 G.n2344 0.686
R6118 G.n2343 G.n2342 0.686
R6119 G.n2240 G.n2239 0.686
R6120 G.n2216 G.n2215 0.686
R6121 G.n2186 G.n2185 0.686
R6122 G.n2151 G.n2150 0.686
R6123 G.n2110 G.n2109 0.686
R6124 G.n2065 G.n2064 0.686
R6125 G.n2014 G.n2013 0.686
R6126 G.n1957 G.n1956 0.686
R6127 G.n1895 G.n1894 0.686
R6128 G.n1827 G.n1826 0.686
R6129 G.n1755 G.n1754 0.686
R6130 G.n1677 G.n1676 0.686
R6131 G.n1594 G.n1593 0.686
R6132 G.n1507 G.n1506 0.686
R6133 G.n1419 G.n1418 0.686
R6134 G.n1331 G.n1330 0.686
R6135 G.n1243 G.n1242 0.686
R6136 G.n1155 G.n1154 0.686
R6137 G.n1067 G.n1066 0.686
R6138 G.n982 G.n981 0.686
R6139 G.n900 G.n899 0.686
R6140 G.n824 G.n823 0.686
R6141 G.n751 G.n750 0.686
R6142 G.n681 G.n680 0.686
R6143 G.n614 G.n613 0.686
R6144 G.n550 G.n549 0.686
R6145 G.n489 G.n488 0.686
R6146 G.n431 G.n430 0.686
R6147 G.n376 G.n375 0.686
R6148 G.n327 G.n326 0.686
R6149 G.n281 G.n280 0.686
R6150 G.n238 G.n237 0.686
R6151 G.n198 G.n197 0.686
R6152 G.n161 G.n160 0.686
R6153 G.n127 G.n126 0.686
R6154 G.n96 G.n95 0.686
R6155 G.n71 G.n70 0.686
R6156 G.n3623 G.n3622 0.686
R6157 G.n3625 G.n3624 0.686
R6158 G.n3627 G.n3626 0.686
R6159 G.n3629 G.n3628 0.686
R6160 G.n3631 G.n3630 0.686
R6161 G.n3633 G.n3632 0.686
R6162 G.n3654 G.n3653 0.686
R6163 G.n3652 G.n3651 0.686
R6164 G.n3650 G.n3649 0.686
R6165 G.n3648 G.n3647 0.686
R6166 G.n3646 G.n3645 0.686
R6167 G.n3644 G.n3643 0.686
R6168 G.n2353 G.n2352 0.686
R6169 G.n2355 G.n2354 0.686
R6170 G.n2357 G.n2356 0.686
R6171 G.n2359 G.n2358 0.686
R6172 G.n2373 G.n2372 0.686
R6173 G.n2371 G.n2370 0.686
R6174 G.n2369 G.n2368 0.686
R6175 G.n2367 G.n2366 0.686
R6176 G.n2210 G.n2209 0.686
R6177 G.n2180 G.n2179 0.686
R6178 G.n2145 G.n2144 0.686
R6179 G.n2104 G.n2103 0.686
R6180 G.n2059 G.n2058 0.686
R6181 G.n2008 G.n2007 0.686
R6182 G.n1951 G.n1950 0.686
R6183 G.n1889 G.n1888 0.686
R6184 G.n1821 G.n1820 0.686
R6185 G.n1749 G.n1748 0.686
R6186 G.n1671 G.n1670 0.686
R6187 G.n1588 G.n1587 0.686
R6188 G.n1501 G.n1500 0.686
R6189 G.n1413 G.n1412 0.686
R6190 G.n1325 G.n1324 0.686
R6191 G.n1237 G.n1236 0.686
R6192 G.n1149 G.n1148 0.686
R6193 G.n1061 G.n1060 0.686
R6194 G.n976 G.n975 0.686
R6195 G.n894 G.n893 0.686
R6196 G.n818 G.n817 0.686
R6197 G.n745 G.n744 0.686
R6198 G.n675 G.n674 0.686
R6199 G.n608 G.n607 0.686
R6200 G.n544 G.n543 0.686
R6201 G.n483 G.n482 0.686
R6202 G.n425 G.n424 0.686
R6203 G.n370 G.n369 0.686
R6204 G.n321 G.n320 0.686
R6205 G.n275 G.n274 0.686
R6206 G.n232 G.n231 0.686
R6207 G.n192 G.n191 0.686
R6208 G.n155 G.n154 0.686
R6209 G.n121 G.n120 0.686
R6210 G.n3666 G.n3665 0.686
R6211 G.n3668 G.n3667 0.686
R6212 G.n3670 G.n3669 0.686
R6213 G.n3672 G.n3671 0.686
R6214 G.n3674 G.n3673 0.686
R6215 G.n3676 G.n3675 0.686
R6216 G.n3678 G.n3677 0.686
R6217 G.n3680 G.n3679 0.686
R6218 G.n3704 G.n3703 0.686
R6219 G.n3702 G.n3701 0.686
R6220 G.n3700 G.n3699 0.686
R6221 G.n3698 G.n3697 0.686
R6222 G.n3696 G.n3695 0.686
R6223 G.n3694 G.n3693 0.686
R6224 G.n3692 G.n3691 0.686
R6225 G.n2382 G.n2381 0.686
R6226 G.n2384 G.n2383 0.686
R6227 G.n2386 G.n2385 0.686
R6228 G.n2388 G.n2387 0.686
R6229 G.n2390 G.n2389 0.686
R6230 G.n2408 G.n2407 0.686
R6231 G.n2406 G.n2405 0.686
R6232 G.n2404 G.n2403 0.686
R6233 G.n2402 G.n2401 0.686
R6234 G.n2400 G.n2399 0.686
R6235 G.n2139 G.n2138 0.686
R6236 G.n2098 G.n2097 0.686
R6237 G.n2053 G.n2052 0.686
R6238 G.n2002 G.n2001 0.686
R6239 G.n1945 G.n1944 0.686
R6240 G.n1883 G.n1882 0.686
R6241 G.n1815 G.n1814 0.686
R6242 G.n1743 G.n1742 0.686
R6243 G.n1665 G.n1664 0.686
R6244 G.n1582 G.n1581 0.686
R6245 G.n1495 G.n1494 0.686
R6246 G.n1407 G.n1406 0.686
R6247 G.n1319 G.n1318 0.686
R6248 G.n1231 G.n1230 0.686
R6249 G.n1143 G.n1142 0.686
R6250 G.n1055 G.n1054 0.686
R6251 G.n970 G.n969 0.686
R6252 G.n888 G.n887 0.686
R6253 G.n812 G.n811 0.686
R6254 G.n739 G.n738 0.686
R6255 G.n669 G.n668 0.686
R6256 G.n602 G.n601 0.686
R6257 G.n538 G.n537 0.686
R6258 G.n477 G.n476 0.686
R6259 G.n419 G.n418 0.686
R6260 G.n364 G.n363 0.686
R6261 G.n315 G.n314 0.686
R6262 G.n269 G.n268 0.686
R6263 G.n226 G.n225 0.686
R6264 G.n186 G.n185 0.686
R6265 G.n149 G.n148 0.686
R6266 G.n3717 G.n3716 0.686
R6267 G.n3719 G.n3718 0.686
R6268 G.n3721 G.n3720 0.686
R6269 G.n3723 G.n3722 0.686
R6270 G.n3725 G.n3724 0.686
R6271 G.n3727 G.n3726 0.686
R6272 G.n3729 G.n3728 0.686
R6273 G.n3731 G.n3730 0.686
R6274 G.n3733 G.n3732 0.686
R6275 G.n3763 G.n3762 0.686
R6276 G.n3761 G.n3760 0.686
R6277 G.n3759 G.n3758 0.686
R6278 G.n3757 G.n3756 0.686
R6279 G.n3755 G.n3754 0.686
R6280 G.n3753 G.n3752 0.686
R6281 G.n3751 G.n3750 0.686
R6282 G.n3749 G.n3748 0.686
R6283 G.n3747 G.n3746 0.686
R6284 G.n2418 G.n2417 0.686
R6285 G.n2420 G.n2419 0.686
R6286 G.n2422 G.n2421 0.686
R6287 G.n2424 G.n2423 0.686
R6288 G.n2426 G.n2425 0.686
R6289 G.n2428 G.n2427 0.686
R6290 G.n2449 G.n2448 0.686
R6291 G.n2447 G.n2446 0.686
R6292 G.n2445 G.n2444 0.686
R6293 G.n2443 G.n2442 0.686
R6294 G.n2441 G.n2440 0.686
R6295 G.n2439 G.n2438 0.686
R6296 G.n2092 G.n2091 0.686
R6297 G.n2047 G.n2046 0.686
R6298 G.n1996 G.n1995 0.686
R6299 G.n1939 G.n1938 0.686
R6300 G.n1877 G.n1876 0.686
R6301 G.n1809 G.n1808 0.686
R6302 G.n1737 G.n1736 0.686
R6303 G.n1659 G.n1658 0.686
R6304 G.n1576 G.n1575 0.686
R6305 G.n1489 G.n1488 0.686
R6306 G.n1401 G.n1400 0.686
R6307 G.n1313 G.n1312 0.686
R6308 G.n1225 G.n1224 0.686
R6309 G.n1137 G.n1136 0.686
R6310 G.n1049 G.n1048 0.686
R6311 G.n964 G.n963 0.686
R6312 G.n882 G.n881 0.686
R6313 G.n806 G.n805 0.686
R6314 G.n733 G.n732 0.686
R6315 G.n663 G.n662 0.686
R6316 G.n596 G.n595 0.686
R6317 G.n532 G.n531 0.686
R6318 G.n471 G.n470 0.686
R6319 G.n413 G.n412 0.686
R6320 G.n358 G.n357 0.686
R6321 G.n309 G.n308 0.686
R6322 G.n263 G.n262 0.686
R6323 G.n220 G.n219 0.686
R6324 G.n3778 G.n3777 0.686
R6325 G.n3780 G.n3779 0.686
R6326 G.n3782 G.n3781 0.686
R6327 G.n3784 G.n3783 0.686
R6328 G.n3786 G.n3785 0.686
R6329 G.n3788 G.n3787 0.686
R6330 G.n3790 G.n3789 0.686
R6331 G.n3792 G.n3791 0.686
R6332 G.n3794 G.n3793 0.686
R6333 G.n3796 G.n3795 0.686
R6334 G.n3798 G.n3797 0.686
R6335 G.n3834 G.n3833 0.686
R6336 G.n3832 G.n3831 0.686
R6337 G.n3830 G.n3829 0.686
R6338 G.n3828 G.n3827 0.686
R6339 G.n3826 G.n3825 0.686
R6340 G.n3824 G.n3823 0.686
R6341 G.n3822 G.n3821 0.686
R6342 G.n3820 G.n3819 0.686
R6343 G.n3818 G.n3817 0.686
R6344 G.n3816 G.n3815 0.686
R6345 G.n3814 G.n3813 0.686
R6346 G.n2460 G.n2459 0.686
R6347 G.n2462 G.n2461 0.686
R6348 G.n2464 G.n2463 0.686
R6349 G.n2466 G.n2465 0.686
R6350 G.n2468 G.n2467 0.686
R6351 G.n2470 G.n2469 0.686
R6352 G.n2472 G.n2471 0.686
R6353 G.n2496 G.n2495 0.686
R6354 G.n2494 G.n2493 0.686
R6355 G.n2492 G.n2491 0.686
R6356 G.n2490 G.n2489 0.686
R6357 G.n2488 G.n2487 0.686
R6358 G.n2486 G.n2485 0.686
R6359 G.n2484 G.n2483 0.686
R6360 G.n2041 G.n2040 0.686
R6361 G.n1990 G.n1989 0.686
R6362 G.n1933 G.n1932 0.686
R6363 G.n1871 G.n1870 0.686
R6364 G.n1803 G.n1802 0.686
R6365 G.n1731 G.n1730 0.686
R6366 G.n1653 G.n1652 0.686
R6367 G.n1570 G.n1569 0.686
R6368 G.n1483 G.n1482 0.686
R6369 G.n1395 G.n1394 0.686
R6370 G.n1307 G.n1306 0.686
R6371 G.n1219 G.n1218 0.686
R6372 G.n1131 G.n1130 0.686
R6373 G.n1043 G.n1042 0.686
R6374 G.n958 G.n957 0.686
R6375 G.n876 G.n875 0.686
R6376 G.n800 G.n799 0.686
R6377 G.n727 G.n726 0.686
R6378 G.n657 G.n656 0.686
R6379 G.n590 G.n589 0.686
R6380 G.n526 G.n525 0.686
R6381 G.n465 G.n464 0.686
R6382 G.n407 G.n406 0.686
R6383 G.n352 G.n351 0.686
R6384 G.n303 G.n302 0.686
R6385 G.n3851 G.n3850 0.686
R6386 G.n3853 G.n3852 0.686
R6387 G.n3855 G.n3854 0.686
R6388 G.n3857 G.n3856 0.686
R6389 G.n3859 G.n3858 0.686
R6390 G.n3861 G.n3860 0.686
R6391 G.n3863 G.n3862 0.686
R6392 G.n3865 G.n3864 0.686
R6393 G.n3867 G.n3866 0.686
R6394 G.n3869 G.n3868 0.686
R6395 G.n3871 G.n3870 0.686
R6396 G.n3873 G.n3872 0.686
R6397 G.n3875 G.n3874 0.686
R6398 G.n3917 G.n3916 0.686
R6399 G.n3915 G.n3914 0.686
R6400 G.n3913 G.n3912 0.686
R6401 G.n3911 G.n3910 0.686
R6402 G.n3909 G.n3908 0.686
R6403 G.n3907 G.n3906 0.686
R6404 G.n3905 G.n3904 0.686
R6405 G.n3903 G.n3902 0.686
R6406 G.n3901 G.n3900 0.686
R6407 G.n3899 G.n3898 0.686
R6408 G.n3897 G.n3896 0.686
R6409 G.n3895 G.n3894 0.686
R6410 G.n3893 G.n3892 0.686
R6411 G.n2510 G.n2509 0.686
R6412 G.n2512 G.n2511 0.686
R6413 G.n2514 G.n2513 0.686
R6414 G.n2516 G.n2515 0.686
R6415 G.n2518 G.n2517 0.686
R6416 G.n2520 G.n2519 0.686
R6417 G.n2522 G.n2521 0.686
R6418 G.n2524 G.n2523 0.686
R6419 G.n2551 G.n2550 0.686
R6420 G.n2549 G.n2548 0.686
R6421 G.n2547 G.n2546 0.686
R6422 G.n2545 G.n2544 0.686
R6423 G.n2543 G.n2542 0.686
R6424 G.n2541 G.n2540 0.686
R6425 G.n2539 G.n2538 0.686
R6426 G.n2537 G.n2536 0.686
R6427 G.n1984 G.n1983 0.686
R6428 G.n1927 G.n1926 0.686
R6429 G.n1865 G.n1864 0.686
R6430 G.n1797 G.n1796 0.686
R6431 G.n1725 G.n1724 0.686
R6432 G.n1647 G.n1646 0.686
R6433 G.n1564 G.n1563 0.686
R6434 G.n1477 G.n1476 0.686
R6435 G.n1389 G.n1388 0.686
R6436 G.n1301 G.n1300 0.686
R6437 G.n1213 G.n1212 0.686
R6438 G.n1125 G.n1124 0.686
R6439 G.n1037 G.n1036 0.686
R6440 G.n952 G.n951 0.686
R6441 G.n870 G.n869 0.686
R6442 G.n794 G.n793 0.686
R6443 G.n721 G.n720 0.686
R6444 G.n651 G.n650 0.686
R6445 G.n584 G.n583 0.686
R6446 G.n520 G.n519 0.686
R6447 G.n459 G.n458 0.686
R6448 G.n401 G.n400 0.686
R6449 G.n3936 G.n3935 0.686
R6450 G.n3938 G.n3937 0.686
R6451 G.n3940 G.n3939 0.686
R6452 G.n3942 G.n3941 0.686
R6453 G.n3944 G.n3943 0.686
R6454 G.n3946 G.n3945 0.686
R6455 G.n3948 G.n3947 0.686
R6456 G.n3950 G.n3949 0.686
R6457 G.n3952 G.n3951 0.686
R6458 G.n3954 G.n3953 0.686
R6459 G.n3956 G.n3955 0.686
R6460 G.n3958 G.n3957 0.686
R6461 G.n3960 G.n3959 0.686
R6462 G.n3962 G.n3961 0.686
R6463 G.n3964 G.n3963 0.686
R6464 G.n4009 G.n4008 0.686
R6465 G.n4007 G.n4006 0.686
R6466 G.n4005 G.n4004 0.686
R6467 G.n4003 G.n4002 0.686
R6468 G.n4001 G.n4000 0.686
R6469 G.n3999 G.n3998 0.686
R6470 G.n3997 G.n3996 0.686
R6471 G.n3995 G.n3994 0.686
R6472 G.n3993 G.n3992 0.686
R6473 G.n3991 G.n3990 0.686
R6474 G.n3989 G.n3988 0.686
R6475 G.n3987 G.n3986 0.686
R6476 G.n3985 G.n3984 0.686
R6477 G.n3983 G.n3982 0.686
R6478 G.n2566 G.n2565 0.686
R6479 G.n2568 G.n2567 0.686
R6480 G.n2570 G.n2569 0.686
R6481 G.n2572 G.n2571 0.686
R6482 G.n2574 G.n2573 0.686
R6483 G.n2576 G.n2575 0.686
R6484 G.n2578 G.n2577 0.686
R6485 G.n2580 G.n2579 0.686
R6486 G.n2582 G.n2581 0.686
R6487 G.n2612 G.n2611 0.686
R6488 G.n2610 G.n2609 0.686
R6489 G.n2608 G.n2607 0.686
R6490 G.n2606 G.n2605 0.686
R6491 G.n2604 G.n2603 0.686
R6492 G.n2602 G.n2601 0.686
R6493 G.n2600 G.n2599 0.686
R6494 G.n2598 G.n2597 0.686
R6495 G.n2596 G.n2595 0.686
R6496 G.n1921 G.n1920 0.686
R6497 G.n1859 G.n1858 0.686
R6498 G.n1791 G.n1790 0.686
R6499 G.n1719 G.n1718 0.686
R6500 G.n1641 G.n1640 0.686
R6501 G.n1558 G.n1557 0.686
R6502 G.n1471 G.n1470 0.686
R6503 G.n1383 G.n1382 0.686
R6504 G.n1295 G.n1294 0.686
R6505 G.n1207 G.n1206 0.686
R6506 G.n1119 G.n1118 0.686
R6507 G.n1031 G.n1030 0.686
R6508 G.n946 G.n945 0.686
R6509 G.n864 G.n863 0.686
R6510 G.n788 G.n787 0.686
R6511 G.n715 G.n714 0.686
R6512 G.n645 G.n644 0.686
R6513 G.n578 G.n577 0.686
R6514 G.n514 G.n513 0.686
R6515 G.n453 G.n452 0.686
R6516 G.n4029 G.n4028 0.686
R6517 G.n4031 G.n4030 0.686
R6518 G.n4033 G.n4032 0.686
R6519 G.n4035 G.n4034 0.686
R6520 G.n4037 G.n4036 0.686
R6521 G.n4039 G.n4038 0.686
R6522 G.n4041 G.n4040 0.686
R6523 G.n4043 G.n4042 0.686
R6524 G.n4045 G.n4044 0.686
R6525 G.n4047 G.n4046 0.686
R6526 G.n4049 G.n4048 0.686
R6527 G.n4051 G.n4050 0.686
R6528 G.n4053 G.n4052 0.686
R6529 G.n4055 G.n4054 0.686
R6530 G.n4057 G.n4056 0.686
R6531 G.n4059 G.n4058 0.686
R6532 G.n4110 G.n4109 0.686
R6533 G.n4108 G.n4107 0.686
R6534 G.n4106 G.n4105 0.686
R6535 G.n4104 G.n4103 0.686
R6536 G.n4102 G.n4101 0.686
R6537 G.n4100 G.n4099 0.686
R6538 G.n4098 G.n4097 0.686
R6539 G.n4096 G.n4095 0.686
R6540 G.n4094 G.n4093 0.686
R6541 G.n4092 G.n4091 0.686
R6542 G.n4090 G.n4089 0.686
R6543 G.n4088 G.n4087 0.686
R6544 G.n4086 G.n4085 0.686
R6545 G.n4084 G.n4083 0.686
R6546 G.n4082 G.n4081 0.686
R6547 G.n4080 G.n4079 0.686
R6548 G.n2627 G.n2626 0.686
R6549 G.n2629 G.n2628 0.686
R6550 G.n2631 G.n2630 0.686
R6551 G.n2633 G.n2632 0.686
R6552 G.n2635 G.n2634 0.686
R6553 G.n2637 G.n2636 0.686
R6554 G.n2639 G.n2638 0.686
R6555 G.n2641 G.n2640 0.686
R6556 G.n2643 G.n2642 0.686
R6557 G.n2645 G.n2644 0.686
R6558 G.n2647 G.n2646 0.686
R6559 G.n2680 G.n2679 0.686
R6560 G.n2678 G.n2677 0.686
R6561 G.n2676 G.n2675 0.686
R6562 G.n2674 G.n2673 0.686
R6563 G.n2672 G.n2671 0.686
R6564 G.n2670 G.n2669 0.686
R6565 G.n2668 G.n2667 0.686
R6566 G.n2666 G.n2665 0.686
R6567 G.n2664 G.n2663 0.686
R6568 G.n2662 G.n2661 0.686
R6569 G.n1853 G.n1852 0.686
R6570 G.n1785 G.n1784 0.686
R6571 G.n1713 G.n1712 0.686
R6572 G.n1635 G.n1634 0.686
R6573 G.n1552 G.n1551 0.686
R6574 G.n1465 G.n1464 0.686
R6575 G.n1377 G.n1376 0.686
R6576 G.n1289 G.n1288 0.686
R6577 G.n1201 G.n1200 0.686
R6578 G.n1113 G.n1112 0.686
R6579 G.n1025 G.n1024 0.686
R6580 G.n940 G.n939 0.686
R6581 G.n858 G.n857 0.686
R6582 G.n782 G.n781 0.686
R6583 G.n709 G.n708 0.686
R6584 G.n639 G.n638 0.686
R6585 G.n572 G.n571 0.686
R6586 G.n4132 G.n4131 0.686
R6587 G.n4134 G.n4133 0.686
R6588 G.n4136 G.n4135 0.686
R6589 G.n4138 G.n4137 0.686
R6590 G.n4140 G.n4139 0.686
R6591 G.n4142 G.n4141 0.686
R6592 G.n4144 G.n4143 0.686
R6593 G.n4146 G.n4145 0.686
R6594 G.n4148 G.n4147 0.686
R6595 G.n4150 G.n4149 0.686
R6596 G.n4152 G.n4151 0.686
R6597 G.n4154 G.n4153 0.686
R6598 G.n4156 G.n4155 0.686
R6599 G.n4158 G.n4157 0.686
R6600 G.n4160 G.n4159 0.686
R6601 G.n4162 G.n4161 0.686
R6602 G.n4164 G.n4163 0.686
R6603 G.n4166 G.n4165 0.686
R6604 G.n4223 G.n4222 0.686
R6605 G.n4221 G.n4220 0.686
R6606 G.n4219 G.n4218 0.686
R6607 G.n4217 G.n4216 0.686
R6608 G.n4215 G.n4214 0.686
R6609 G.n4213 G.n4212 0.686
R6610 G.n4211 G.n4210 0.686
R6611 G.n4209 G.n4208 0.686
R6612 G.n4207 G.n4206 0.686
R6613 G.n4205 G.n4204 0.686
R6614 G.n4203 G.n4202 0.686
R6615 G.n4201 G.n4200 0.686
R6616 G.n4199 G.n4198 0.686
R6617 G.n4197 G.n4196 0.686
R6618 G.n4195 G.n4194 0.686
R6619 G.n4193 G.n4192 0.686
R6620 G.n4191 G.n4190 0.686
R6621 G.n4189 G.n4188 0.686
R6622 G.n2696 G.n2695 0.686
R6623 G.n2698 G.n2697 0.686
R6624 G.n2700 G.n2699 0.686
R6625 G.n2702 G.n2701 0.686
R6626 G.n2704 G.n2703 0.686
R6627 G.n2706 G.n2705 0.686
R6628 G.n2708 G.n2707 0.686
R6629 G.n2710 G.n2709 0.686
R6630 G.n2712 G.n2711 0.686
R6631 G.n2714 G.n2713 0.686
R6632 G.n2716 G.n2715 0.686
R6633 G.n2718 G.n2717 0.686
R6634 G.n2754 G.n2753 0.686
R6635 G.n2752 G.n2751 0.686
R6636 G.n2750 G.n2749 0.686
R6637 G.n2748 G.n2747 0.686
R6638 G.n2746 G.n2745 0.686
R6639 G.n2744 G.n2743 0.686
R6640 G.n2742 G.n2741 0.686
R6641 G.n2740 G.n2739 0.686
R6642 G.n2738 G.n2737 0.686
R6643 G.n2736 G.n2735 0.686
R6644 G.n2734 G.n2733 0.686
R6645 G.n1779 G.n1778 0.686
R6646 G.n1707 G.n1706 0.686
R6647 G.n1629 G.n1628 0.686
R6648 G.n1546 G.n1545 0.686
R6649 G.n1459 G.n1458 0.686
R6650 G.n1371 G.n1370 0.686
R6651 G.n1283 G.n1282 0.686
R6652 G.n1195 G.n1194 0.686
R6653 G.n1107 G.n1106 0.686
R6654 G.n1019 G.n1018 0.686
R6655 G.n934 G.n933 0.686
R6656 G.n852 G.n851 0.686
R6657 G.n776 G.n775 0.686
R6658 G.n703 G.n702 0.686
R6659 G.n4247 G.n4246 0.686
R6660 G.n4249 G.n4248 0.686
R6661 G.n4251 G.n4250 0.686
R6662 G.n4253 G.n4252 0.686
R6663 G.n4255 G.n4254 0.686
R6664 G.n4257 G.n4256 0.686
R6665 G.n4259 G.n4258 0.686
R6666 G.n4261 G.n4260 0.686
R6667 G.n4263 G.n4262 0.686
R6668 G.n4265 G.n4264 0.686
R6669 G.n4267 G.n4266 0.686
R6670 G.n4269 G.n4268 0.686
R6671 G.n4271 G.n4270 0.686
R6672 G.n4273 G.n4272 0.686
R6673 G.n4275 G.n4274 0.686
R6674 G.n4277 G.n4276 0.686
R6675 G.n4279 G.n4278 0.686
R6676 G.n4281 G.n4280 0.686
R6677 G.n4283 G.n4282 0.686
R6678 G.n4285 G.n4284 0.686
R6679 G.n4348 G.n4347 0.686
R6680 G.n4346 G.n4345 0.686
R6681 G.n4344 G.n4343 0.686
R6682 G.n4342 G.n4341 0.686
R6683 G.n4340 G.n4339 0.686
R6684 G.n4338 G.n4337 0.686
R6685 G.n4336 G.n4335 0.686
R6686 G.n4334 G.n4333 0.686
R6687 G.n4332 G.n4331 0.686
R6688 G.n4330 G.n4329 0.686
R6689 G.n4328 G.n4327 0.686
R6690 G.n4326 G.n4325 0.686
R6691 G.n4324 G.n4323 0.686
R6692 G.n4322 G.n4321 0.686
R6693 G.n4320 G.n4319 0.686
R6694 G.n4318 G.n4317 0.686
R6695 G.n4316 G.n4315 0.686
R6696 G.n4314 G.n4313 0.686
R6697 G.n4312 G.n4311 0.686
R6698 G.n4310 G.n4309 0.686
R6699 G.n2771 G.n2770 0.686
R6700 G.n2773 G.n2772 0.686
R6701 G.n2775 G.n2774 0.686
R6702 G.n2777 G.n2776 0.686
R6703 G.n2779 G.n2778 0.686
R6704 G.n2781 G.n2780 0.686
R6705 G.n2783 G.n2782 0.686
R6706 G.n2785 G.n2784 0.686
R6707 G.n2787 G.n2786 0.686
R6708 G.n2789 G.n2788 0.686
R6709 G.n2791 G.n2790 0.686
R6710 G.n2793 G.n2792 0.686
R6711 G.n2795 G.n2794 0.686
R6712 G.n2836 G.n2835 0.686
R6713 G.n2834 G.n2833 0.686
R6714 G.n2832 G.n2831 0.686
R6715 G.n2830 G.n2829 0.686
R6716 G.n2828 G.n2827 0.686
R6717 G.n2826 G.n2825 0.686
R6718 G.n2824 G.n2823 0.686
R6719 G.n2822 G.n2821 0.686
R6720 G.n2820 G.n2819 0.686
R6721 G.n2818 G.n2817 0.686
R6722 G.n2816 G.n2815 0.686
R6723 G.n2814 G.n2813 0.686
R6724 G.n2812 G.n2811 0.686
R6725 G.n1701 G.n1700 0.686
R6726 G.n1623 G.n1622 0.686
R6727 G.n1540 G.n1539 0.686
R6728 G.n1453 G.n1452 0.686
R6729 G.n1365 G.n1364 0.686
R6730 G.n1277 G.n1276 0.686
R6731 G.n1189 G.n1188 0.686
R6732 G.n1101 G.n1100 0.686
R6733 G.n1013 G.n1012 0.686
R6734 G.n928 G.n927 0.686
R6735 G.n846 G.n845 0.686
R6736 G.n4374 G.n4373 0.686
R6737 G.n4376 G.n4375 0.686
R6738 G.n4378 G.n4377 0.686
R6739 G.n4380 G.n4379 0.686
R6740 G.n4382 G.n4381 0.686
R6741 G.n4384 G.n4383 0.686
R6742 G.n4386 G.n4385 0.686
R6743 G.n4388 G.n4387 0.686
R6744 G.n4390 G.n4389 0.686
R6745 G.n4392 G.n4391 0.686
R6746 G.n4394 G.n4393 0.686
R6747 G.n4396 G.n4395 0.686
R6748 G.n4398 G.n4397 0.686
R6749 G.n4400 G.n4399 0.686
R6750 G.n4402 G.n4401 0.686
R6751 G.n4404 G.n4403 0.686
R6752 G.n4406 G.n4405 0.686
R6753 G.n4408 G.n4407 0.686
R6754 G.n4410 G.n4409 0.686
R6755 G.n4412 G.n4411 0.686
R6756 G.n4414 G.n4413 0.686
R6757 G.n4416 G.n4415 0.686
R6758 G.n4485 G.n4484 0.686
R6759 G.n4483 G.n4482 0.686
R6760 G.n4481 G.n4480 0.686
R6761 G.n4479 G.n4478 0.686
R6762 G.n4477 G.n4476 0.686
R6763 G.n4475 G.n4474 0.686
R6764 G.n4473 G.n4472 0.686
R6765 G.n4471 G.n4470 0.686
R6766 G.n4469 G.n4468 0.686
R6767 G.n4467 G.n4466 0.686
R6768 G.n4465 G.n4464 0.686
R6769 G.n4463 G.n4462 0.686
R6770 G.n4461 G.n4460 0.686
R6771 G.n4459 G.n4458 0.686
R6772 G.n4457 G.n4456 0.686
R6773 G.n4455 G.n4454 0.686
R6774 G.n4453 G.n4452 0.686
R6775 G.n4451 G.n4450 0.686
R6776 G.n4449 G.n4448 0.686
R6777 G.n4447 G.n4446 0.686
R6778 G.n4445 G.n4444 0.686
R6779 G.n4443 G.n4442 0.686
R6780 G.n2854 G.n2853 0.686
R6781 G.n2856 G.n2855 0.686
R6782 G.n2858 G.n2857 0.686
R6783 G.n2860 G.n2859 0.686
R6784 G.n2862 G.n2861 0.686
R6785 G.n2864 G.n2863 0.686
R6786 G.n2866 G.n2865 0.686
R6787 G.n2868 G.n2867 0.686
R6788 G.n2870 G.n2869 0.686
R6789 G.n2872 G.n2871 0.686
R6790 G.n2874 G.n2873 0.686
R6791 G.n2876 G.n2875 0.686
R6792 G.n2878 G.n2877 0.686
R6793 G.n2880 G.n2879 0.686
R6794 G.n2925 G.n2924 0.686
R6795 G.n2923 G.n2922 0.686
R6796 G.n2921 G.n2920 0.686
R6797 G.n2919 G.n2918 0.686
R6798 G.n2917 G.n2916 0.686
R6799 G.n2915 G.n2914 0.686
R6800 G.n2913 G.n2912 0.686
R6801 G.n2911 G.n2910 0.686
R6802 G.n2909 G.n2908 0.686
R6803 G.n2907 G.n2906 0.686
R6804 G.n2905 G.n2904 0.686
R6805 G.n2903 G.n2902 0.686
R6806 G.n2901 G.n2900 0.686
R6807 G.n2899 G.n2898 0.686
R6808 G.n1534 G.n1533 0.686
R6809 G.n1447 G.n1446 0.686
R6810 G.n1359 G.n1358 0.686
R6811 G.n1271 G.n1270 0.686
R6812 G.n1183 G.n1182 0.686
R6813 G.n1095 G.n1094 0.686
R6814 G.n1007 G.n1006 0.686
R6815 G.n922 G.n921 0.686
R6816 G.n4512 G.n4511 0.686
R6817 G.n4514 G.n4513 0.686
R6818 G.n4516 G.n4515 0.686
R6819 G.n4518 G.n4517 0.686
R6820 G.n4520 G.n4519 0.686
R6821 G.n4522 G.n4521 0.686
R6822 G.n4524 G.n4523 0.686
R6823 G.n4526 G.n4525 0.686
R6824 G.n4528 G.n4527 0.686
R6825 G.n4530 G.n4529 0.686
R6826 G.n4532 G.n4531 0.686
R6827 G.n4534 G.n4533 0.686
R6828 G.n4536 G.n4535 0.686
R6829 G.n4538 G.n4537 0.686
R6830 G.n4540 G.n4539 0.686
R6831 G.n4542 G.n4541 0.686
R6832 G.n4544 G.n4543 0.686
R6833 G.n4546 G.n4545 0.686
R6834 G.n4548 G.n4547 0.686
R6835 G.n4550 G.n4549 0.686
R6836 G.n4552 G.n4551 0.686
R6837 G.n4554 G.n4553 0.686
R6838 G.n4556 G.n4555 0.686
R6839 G.n4628 G.n4627 0.686
R6840 G.n4626 G.n4625 0.686
R6841 G.n4624 G.n4623 0.686
R6842 G.n4622 G.n4621 0.686
R6843 G.n4620 G.n4619 0.686
R6844 G.n4618 G.n4617 0.686
R6845 G.n4616 G.n4615 0.686
R6846 G.n4614 G.n4613 0.686
R6847 G.n4612 G.n4611 0.686
R6848 G.n4610 G.n4609 0.686
R6849 G.n4608 G.n4607 0.686
R6850 G.n4606 G.n4605 0.686
R6851 G.n4604 G.n4603 0.686
R6852 G.n4602 G.n4601 0.686
R6853 G.n4600 G.n4599 0.686
R6854 G.n4598 G.n4597 0.686
R6855 G.n4596 G.n4595 0.686
R6856 G.n4594 G.n4593 0.686
R6857 G.n4592 G.n4591 0.686
R6858 G.n4590 G.n4589 0.686
R6859 G.n4588 G.n4587 0.686
R6860 G.n4586 G.n4585 0.686
R6861 G.n4584 G.n4583 0.686
R6862 G.n2944 G.n2943 0.686
R6863 G.n2946 G.n2945 0.686
R6864 G.n2948 G.n2947 0.686
R6865 G.n2950 G.n2949 0.686
R6866 G.n2952 G.n2951 0.686
R6867 G.n2954 G.n2953 0.686
R6868 G.n2956 G.n2955 0.686
R6869 G.n2958 G.n2957 0.686
R6870 G.n2960 G.n2959 0.686
R6871 G.n2962 G.n2961 0.686
R6872 G.n2964 G.n2963 0.686
R6873 G.n2966 G.n2965 0.686
R6874 G.n2968 G.n2967 0.686
R6875 G.n2970 G.n2969 0.686
R6876 G.n2972 G.n2971 0.686
R6877 G.n3020 G.n3019 0.686
R6878 G.n3018 G.n3017 0.686
R6879 G.n3016 G.n3015 0.686
R6880 G.n3014 G.n3013 0.686
R6881 G.n3012 G.n3011 0.686
R6882 G.n3010 G.n3009 0.686
R6883 G.n3008 G.n3007 0.686
R6884 G.n3006 G.n3005 0.686
R6885 G.n3004 G.n3003 0.686
R6886 G.n3002 G.n3001 0.686
R6887 G.n3000 G.n2999 0.686
R6888 G.n2998 G.n2997 0.686
R6889 G.n2996 G.n2995 0.686
R6890 G.n2994 G.n2993 0.686
R6891 G.n2992 G.n2991 0.686
R6892 G.n1441 G.n1440 0.686
R6893 G.n1353 G.n1352 0.686
R6894 G.n1265 G.n1264 0.686
R6895 G.n1177 G.n1176 0.686
R6896 G.n1089 G.n1088 0.686
R6897 G.n4657 G.n4656 0.686
R6898 G.n4659 G.n4658 0.686
R6899 G.n4661 G.n4660 0.686
R6900 G.n4663 G.n4662 0.686
R6901 G.n4665 G.n4664 0.686
R6902 G.n4667 G.n4666 0.686
R6903 G.n4669 G.n4668 0.686
R6904 G.n4671 G.n4670 0.686
R6905 G.n4673 G.n4672 0.686
R6906 G.n4675 G.n4674 0.686
R6907 G.n4677 G.n4676 0.686
R6908 G.n4679 G.n4678 0.686
R6909 G.n4681 G.n4680 0.686
R6910 G.n4683 G.n4682 0.686
R6911 G.n4685 G.n4684 0.686
R6912 G.n4687 G.n4686 0.686
R6913 G.n4689 G.n4688 0.686
R6914 G.n4691 G.n4690 0.686
R6915 G.n4693 G.n4692 0.686
R6916 G.n4695 G.n4694 0.686
R6917 G.n4697 G.n4696 0.686
R6918 G.n4699 G.n4698 0.686
R6919 G.n4701 G.n4700 0.686
R6920 G.n4703 G.n4702 0.686
R6921 G.n4705 G.n4704 0.686
R6922 G.n4782 G.n4781 0.686
R6923 G.n4780 G.n4779 0.686
R6924 G.n4778 G.n4777 0.686
R6925 G.n4776 G.n4775 0.686
R6926 G.n4774 G.n4773 0.686
R6927 G.n4772 G.n4771 0.686
R6928 G.n4770 G.n4769 0.686
R6929 G.n4768 G.n4767 0.686
R6930 G.n4766 G.n4765 0.686
R6931 G.n4764 G.n4763 0.686
R6932 G.n4762 G.n4761 0.686
R6933 G.n4760 G.n4759 0.686
R6934 G.n4758 G.n4757 0.686
R6935 G.n4756 G.n4755 0.686
R6936 G.n4754 G.n4753 0.686
R6937 G.n4752 G.n4751 0.686
R6938 G.n4750 G.n4749 0.686
R6939 G.n4748 G.n4747 0.686
R6940 G.n4746 G.n4745 0.686
R6941 G.n4744 G.n4743 0.686
R6942 G.n4742 G.n4741 0.686
R6943 G.n4740 G.n4739 0.686
R6944 G.n4738 G.n4737 0.686
R6945 G.n4736 G.n4735 0.686
R6946 G.n4734 G.n4733 0.686
R6947 G.n3039 G.n3038 0.686
R6948 G.n3041 G.n3040 0.686
R6949 G.n3043 G.n3042 0.686
R6950 G.n3045 G.n3044 0.686
R6951 G.n3047 G.n3046 0.686
R6952 G.n3049 G.n3048 0.686
R6953 G.n3051 G.n3050 0.686
R6954 G.n3053 G.n3052 0.686
R6955 G.n3055 G.n3054 0.686
R6956 G.n3057 G.n3056 0.686
R6957 G.n3059 G.n3058 0.686
R6958 G.n3061 G.n3060 0.686
R6959 G.n3063 G.n3062 0.686
R6960 G.n3065 G.n3064 0.686
R6961 G.n3067 G.n3066 0.686
R6962 G.n3069 G.n3068 0.686
R6963 G.n3113 G.n3112 0.686
R6964 G.n3111 G.n3110 0.686
R6965 G.n3109 G.n3108 0.686
R6966 G.n3107 G.n3106 0.686
R6967 G.n3105 G.n3104 0.686
R6968 G.n3103 G.n3102 0.686
R6969 G.n3101 G.n3100 0.686
R6970 G.n3099 G.n3098 0.686
R6971 G.n3097 G.n3096 0.686
R6972 G.n3095 G.n3094 0.686
R6973 G.n3093 G.n3092 0.686
R6974 G.n3091 G.n3090 0.686
R6975 G.n3089 G.n3088 0.686
R6976 G.n3087 G.n3086 0.686
R6977 G.n6357 G.n6356 0.686
R6978 G.n6304 G.n6303 0.686
R6979 G.n6250 G.n6249 0.686
R6980 G.n6196 G.n6195 0.686
R6981 G.n6142 G.n6141 0.686
R6982 G.n6088 G.n6087 0.686
R6983 G.n6036 G.n6035 0.686
R6984 G.n4809 G.n4808 0.686
R6985 G.n4811 G.n4810 0.686
R6986 G.n4813 G.n4812 0.686
R6987 G.n4815 G.n4814 0.686
R6988 G.n4817 G.n4816 0.686
R6989 G.n4819 G.n4818 0.686
R6990 G.n4821 G.n4820 0.686
R6991 G.n4823 G.n4822 0.686
R6992 G.n4825 G.n4824 0.686
R6993 G.n4827 G.n4826 0.686
R6994 G.n4829 G.n4828 0.686
R6995 G.n4831 G.n4830 0.686
R6996 G.n4833 G.n4832 0.686
R6997 G.n4835 G.n4834 0.686
R6998 G.n4837 G.n4836 0.686
R6999 G.n4839 G.n4838 0.686
R7000 G.n4841 G.n4840 0.686
R7001 G.n4843 G.n4842 0.686
R7002 G.n4845 G.n4844 0.686
R7003 G.n4847 G.n4846 0.686
R7004 G.n4849 G.n4848 0.686
R7005 G.n4851 G.n4850 0.686
R7006 G.n4853 G.n4852 0.686
R7007 G.n4855 G.n4854 0.686
R7008 G.n4923 G.n4922 0.686
R7009 G.n4921 G.n4920 0.686
R7010 G.n4919 G.n4918 0.686
R7011 G.n4917 G.n4916 0.686
R7012 G.n4915 G.n4914 0.686
R7013 G.n4913 G.n4912 0.686
R7014 G.n4911 G.n4910 0.686
R7015 G.n4909 G.n4908 0.686
R7016 G.n4907 G.n4906 0.686
R7017 G.n4905 G.n4904 0.686
R7018 G.n4903 G.n4902 0.686
R7019 G.n4901 G.n4900 0.686
R7020 G.n4899 G.n4898 0.686
R7021 G.n4897 G.n4896 0.686
R7022 G.n4895 G.n4894 0.686
R7023 G.n4893 G.n4892 0.686
R7024 G.n4891 G.n4890 0.686
R7025 G.n4889 G.n4888 0.686
R7026 G.n4887 G.n4886 0.686
R7027 G.n4885 G.n4884 0.686
R7028 G.n4883 G.n4882 0.686
R7029 G.n4881 G.n4880 0.686
R7030 G.n3131 G.n3130 0.686
R7031 G.n3133 G.n3132 0.686
R7032 G.n3135 G.n3134 0.686
R7033 G.n3137 G.n3136 0.686
R7034 G.n3139 G.n3138 0.686
R7035 G.n3141 G.n3140 0.686
R7036 G.n3143 G.n3142 0.686
R7037 G.n3145 G.n3144 0.686
R7038 G.n3147 G.n3146 0.686
R7039 G.n3149 G.n3148 0.686
R7040 G.n3151 G.n3150 0.686
R7041 G.n3153 G.n3152 0.686
R7042 G.n3155 G.n3154 0.686
R7043 G.n3157 G.n3156 0.686
R7044 G.n3196 G.n3195 0.686
R7045 G.n3194 G.n3193 0.686
R7046 G.n3192 G.n3191 0.686
R7047 G.n3190 G.n3189 0.686
R7048 G.n3188 G.n3187 0.686
R7049 G.n3186 G.n3185 0.686
R7050 G.n3184 G.n3183 0.686
R7051 G.n3182 G.n3181 0.686
R7052 G.n3180 G.n3179 0.686
R7053 G.n3178 G.n3177 0.686
R7054 G.n3176 G.n3175 0.686
R7055 G.n3174 G.n3173 0.686
R7056 G.n6461 G.n6460 0.686
R7057 G.n6413 G.n6412 0.686
R7058 G.n6362 G.n6361 0.686
R7059 G.n6309 G.n6308 0.686
R7060 G.n6255 G.n6254 0.686
R7061 G.n6201 G.n6200 0.686
R7062 G.n6147 G.n6146 0.686
R7063 G.n6093 G.n6092 0.686
R7064 G.n6041 G.n6040 0.686
R7065 G.n5990 G.n5989 0.686
R7066 G.n5941 G.n5940 0.686
R7067 G.n5895 G.n5894 0.686
R7068 G.n4947 G.n4946 0.686
R7069 G.n4949 G.n4948 0.686
R7070 G.n4951 G.n4950 0.686
R7071 G.n4953 G.n4952 0.686
R7072 G.n4955 G.n4954 0.686
R7073 G.n4957 G.n4956 0.686
R7074 G.n4959 G.n4958 0.686
R7075 G.n4961 G.n4960 0.686
R7076 G.n4963 G.n4962 0.686
R7077 G.n4965 G.n4964 0.686
R7078 G.n4967 G.n4966 0.686
R7079 G.n4969 G.n4968 0.686
R7080 G.n4971 G.n4970 0.686
R7081 G.n4973 G.n4972 0.686
R7082 G.n4975 G.n4974 0.686
R7083 G.n4977 G.n4976 0.686
R7084 G.n4979 G.n4978 0.686
R7085 G.n4981 G.n4980 0.686
R7086 G.n4983 G.n4982 0.686
R7087 G.n4985 G.n4984 0.686
R7088 G.n4987 G.n4986 0.686
R7089 G.n5046 G.n5045 0.686
R7090 G.n5044 G.n5043 0.686
R7091 G.n5042 G.n5041 0.686
R7092 G.n5040 G.n5039 0.686
R7093 G.n5038 G.n5037 0.686
R7094 G.n5036 G.n5035 0.686
R7095 G.n5034 G.n5033 0.686
R7096 G.n5032 G.n5031 0.686
R7097 G.n5030 G.n5029 0.686
R7098 G.n5028 G.n5027 0.686
R7099 G.n5026 G.n5025 0.686
R7100 G.n5024 G.n5023 0.686
R7101 G.n5022 G.n5021 0.686
R7102 G.n5020 G.n5019 0.686
R7103 G.n5018 G.n5017 0.686
R7104 G.n5016 G.n5015 0.686
R7105 G.n5014 G.n5013 0.686
R7106 G.n5012 G.n5011 0.686
R7107 G.n5010 G.n5009 0.686
R7108 G.n3212 G.n3211 0.686
R7109 G.n3214 G.n3213 0.686
R7110 G.n3216 G.n3215 0.686
R7111 G.n3218 G.n3217 0.686
R7112 G.n3220 G.n3219 0.686
R7113 G.n3222 G.n3221 0.686
R7114 G.n3224 G.n3223 0.686
R7115 G.n3226 G.n3225 0.686
R7116 G.n3228 G.n3227 0.686
R7117 G.n3230 G.n3229 0.686
R7118 G.n3232 G.n3231 0.686
R7119 G.n3234 G.n3233 0.686
R7120 G.n3268 G.n3267 0.686
R7121 G.n3266 G.n3265 0.686
R7122 G.n3264 G.n3263 0.686
R7123 G.n3262 G.n3261 0.686
R7124 G.n3260 G.n3259 0.686
R7125 G.n3258 G.n3257 0.686
R7126 G.n3256 G.n3255 0.686
R7127 G.n3254 G.n3253 0.686
R7128 G.n3252 G.n3251 0.686
R7129 G.n3250 G.n3249 0.686
R7130 G.n3248 G.n3247 0.686
R7131 G.n6551 G.n6550 0.686
R7132 G.n6510 G.n6509 0.686
R7133 G.n6466 G.n6465 0.686
R7134 G.n6418 G.n6417 0.686
R7135 G.n6367 G.n6366 0.686
R7136 G.n6314 G.n6313 0.686
R7137 G.n6260 G.n6259 0.686
R7138 G.n6206 G.n6205 0.686
R7139 G.n6152 G.n6151 0.686
R7140 G.n6098 G.n6097 0.686
R7141 G.n6046 G.n6045 0.686
R7142 G.n5995 G.n5994 0.686
R7143 G.n5946 G.n5945 0.686
R7144 G.n5900 G.n5899 0.686
R7145 G.n5855 G.n5854 0.686
R7146 G.n5812 G.n5811 0.686
R7147 G.n5772 G.n5771 0.686
R7148 G.n5067 G.n5066 0.686
R7149 G.n5069 G.n5068 0.686
R7150 G.n5071 G.n5070 0.686
R7151 G.n5073 G.n5072 0.686
R7152 G.n5075 G.n5074 0.686
R7153 G.n5077 G.n5076 0.686
R7154 G.n5079 G.n5078 0.686
R7155 G.n5081 G.n5080 0.686
R7156 G.n5083 G.n5082 0.686
R7157 G.n5085 G.n5084 0.686
R7158 G.n5087 G.n5086 0.686
R7159 G.n5089 G.n5088 0.686
R7160 G.n5091 G.n5090 0.686
R7161 G.n5093 G.n5092 0.686
R7162 G.n5095 G.n5094 0.686
R7163 G.n5097 G.n5096 0.686
R7164 G.n5099 G.n5098 0.686
R7165 G.n5101 G.n5100 0.686
R7166 G.n5151 G.n5150 0.686
R7167 G.n5149 G.n5148 0.686
R7168 G.n5147 G.n5146 0.686
R7169 G.n5145 G.n5144 0.686
R7170 G.n5143 G.n5142 0.686
R7171 G.n5141 G.n5140 0.686
R7172 G.n5139 G.n5138 0.686
R7173 G.n5137 G.n5136 0.686
R7174 G.n5135 G.n5134 0.686
R7175 G.n5133 G.n5132 0.686
R7176 G.n5131 G.n5130 0.686
R7177 G.n5129 G.n5128 0.686
R7178 G.n5127 G.n5126 0.686
R7179 G.n5125 G.n5124 0.686
R7180 G.n5123 G.n5122 0.686
R7181 G.n5121 G.n5120 0.686
R7182 G.n3283 G.n3282 0.686
R7183 G.n3285 G.n3284 0.686
R7184 G.n3287 G.n3286 0.686
R7185 G.n3289 G.n3288 0.686
R7186 G.n3291 G.n3290 0.686
R7187 G.n3293 G.n3292 0.686
R7188 G.n3295 G.n3294 0.686
R7189 G.n3297 G.n3296 0.686
R7190 G.n3299 G.n3298 0.686
R7191 G.n3301 G.n3300 0.686
R7192 G.n3330 G.n3329 0.686
R7193 G.n3328 G.n3327 0.686
R7194 G.n3326 G.n3325 0.686
R7195 G.n3324 G.n3323 0.686
R7196 G.n3322 G.n3321 0.686
R7197 G.n3320 G.n3319 0.686
R7198 G.n3318 G.n3317 0.686
R7199 G.n3316 G.n3315 0.686
R7200 G.n3314 G.n3313 0.686
R7201 G.n6593 G.n6592 0.686
R7202 G.n6556 G.n6555 0.686
R7203 G.n6515 G.n6514 0.686
R7204 G.n6471 G.n6470 0.686
R7205 G.n6423 G.n6422 0.686
R7206 G.n6372 G.n6371 0.686
R7207 G.n6319 G.n6318 0.686
R7208 G.n6265 G.n6264 0.686
R7209 G.n6211 G.n6210 0.686
R7210 G.n6157 G.n6156 0.686
R7211 G.n6103 G.n6102 0.686
R7212 G.n6051 G.n6050 0.686
R7213 G.n6000 G.n5999 0.686
R7214 G.n5951 G.n5950 0.686
R7215 G.n5905 G.n5904 0.686
R7216 G.n5860 G.n5859 0.686
R7217 G.n5817 G.n5816 0.686
R7218 G.n5777 G.n5776 0.686
R7219 G.n5738 G.n5737 0.686
R7220 G.n5701 G.n5700 0.686
R7221 G.n5169 G.n5168 0.686
R7222 G.n5171 G.n5170 0.686
R7223 G.n5173 G.n5172 0.686
R7224 G.n5175 G.n5174 0.686
R7225 G.n5177 G.n5176 0.686
R7226 G.n5179 G.n5178 0.686
R7227 G.n5181 G.n5180 0.686
R7228 G.n5183 G.n5182 0.686
R7229 G.n5185 G.n5184 0.686
R7230 G.n5187 G.n5186 0.686
R7231 G.n5189 G.n5188 0.686
R7232 G.n5191 G.n5190 0.686
R7233 G.n5193 G.n5192 0.686
R7234 G.n5195 G.n5194 0.686
R7235 G.n5197 G.n5196 0.686
R7236 G.n5199 G.n5198 0.686
R7237 G.n5240 G.n5239 0.686
R7238 G.n5238 G.n5237 0.686
R7239 G.n5236 G.n5235 0.686
R7240 G.n5234 G.n5233 0.686
R7241 G.n5232 G.n5231 0.686
R7242 G.n5230 G.n5229 0.686
R7243 G.n5228 G.n5227 0.686
R7244 G.n5226 G.n5225 0.686
R7245 G.n5224 G.n5223 0.686
R7246 G.n5222 G.n5221 0.686
R7247 G.n5220 G.n5219 0.686
R7248 G.n5218 G.n5217 0.686
R7249 G.n5216 G.n5215 0.686
R7250 G.n3342 G.n3341 0.686
R7251 G.n3344 G.n3343 0.686
R7252 G.n3346 G.n3345 0.686
R7253 G.n3348 G.n3347 0.686
R7254 G.n3350 G.n3349 0.686
R7255 G.n3352 G.n3351 0.686
R7256 G.n3354 G.n3353 0.686
R7257 G.n3356 G.n3355 0.686
R7258 G.n3358 G.n3357 0.686
R7259 G.n3381 G.n3380 0.686
R7260 G.n3379 G.n3378 0.686
R7261 G.n3377 G.n3376 0.686
R7262 G.n3375 G.n3374 0.686
R7263 G.n3373 G.n3372 0.686
R7264 G.n3371 G.n3370 0.686
R7265 G.n3369 G.n3368 0.686
R7266 G.n6661 G.n6660 0.686
R7267 G.n6631 G.n6630 0.686
R7268 G.n6598 G.n6597 0.686
R7269 G.n6561 G.n6560 0.686
R7270 G.n6520 G.n6519 0.686
R7271 G.n6476 G.n6475 0.686
R7272 G.n6428 G.n6427 0.686
R7273 G.n6377 G.n6376 0.686
R7274 G.n6324 G.n6323 0.686
R7275 G.n6270 G.n6269 0.686
R7276 G.n6216 G.n6215 0.686
R7277 G.n6162 G.n6161 0.686
R7278 G.n6108 G.n6107 0.686
R7279 G.n6056 G.n6055 0.686
R7280 G.n6005 G.n6004 0.686
R7281 G.n5956 G.n5955 0.686
R7282 G.n5910 G.n5909 0.686
R7283 G.n5865 G.n5864 0.686
R7284 G.n5822 G.n5821 0.686
R7285 G.n5782 G.n5781 0.686
R7286 G.n5743 G.n5742 0.686
R7287 G.n5706 G.n5705 0.686
R7288 G.n5672 G.n5671 0.686
R7289 G.n5641 G.n5640 0.686
R7290 G.n5610 G.n5609 0.686
R7291 G.n5255 G.n5254 0.686
R7292 G.n5257 G.n5256 0.686
R7293 G.n5259 G.n5258 0.686
R7294 G.n5261 G.n5260 0.686
R7295 G.n5263 G.n5262 0.686
R7296 G.n5265 G.n5264 0.686
R7297 G.n5267 G.n5266 0.686
R7298 G.n5269 G.n5268 0.686
R7299 G.n5271 G.n5270 0.686
R7300 G.n5273 G.n5272 0.686
R7301 G.n5275 G.n5274 0.686
R7302 G.n5277 G.n5276 0.686
R7303 G.n5279 G.n5278 0.686
R7304 G.n5311 G.n5310 0.686
R7305 G.n5309 G.n5308 0.686
R7306 G.n5307 G.n5306 0.686
R7307 G.n5305 G.n5304 0.686
R7308 G.n5303 G.n5302 0.686
R7309 G.n5301 G.n5300 0.686
R7310 G.n5299 G.n5298 0.686
R7311 G.n5297 G.n5296 0.686
R7312 G.n5295 G.n5294 0.686
R7313 G.n5293 G.n5292 0.686
R7314 G.n3391 G.n3390 0.686
R7315 G.n3393 G.n3392 0.686
R7316 G.n3395 G.n3394 0.686
R7317 G.n3397 G.n3396 0.686
R7318 G.n3399 G.n3398 0.686
R7319 G.n3401 G.n3400 0.686
R7320 G.n3403 G.n3402 0.686
R7321 G.n3420 G.n3419 0.686
R7322 G.n3418 G.n3417 0.686
R7323 G.n3416 G.n3415 0.686
R7324 G.n3414 G.n3413 0.686
R7325 G.n3412 G.n3411 0.686
R7326 G.n6717 G.n6716 0.686
R7327 G.n6693 G.n6692 0.686
R7328 G.n6666 G.n6665 0.686
R7329 G.n6636 G.n6635 0.686
R7330 G.n6603 G.n6602 0.686
R7331 G.n6566 G.n6565 0.686
R7332 G.n6525 G.n6524 0.686
R7333 G.n6481 G.n6480 0.686
R7334 G.n6433 G.n6432 0.686
R7335 G.n6382 G.n6381 0.686
R7336 G.n6329 G.n6328 0.686
R7337 G.n6275 G.n6274 0.686
R7338 G.n6221 G.n6220 0.686
R7339 G.n6167 G.n6166 0.686
R7340 G.n6113 G.n6112 0.686
R7341 G.n6061 G.n6060 0.686
R7342 G.n6010 G.n6009 0.686
R7343 G.n5961 G.n5960 0.686
R7344 G.n5915 G.n5914 0.686
R7345 G.n5870 G.n5869 0.686
R7346 G.n5827 G.n5826 0.686
R7347 G.n5787 G.n5786 0.686
R7348 G.n5748 G.n5747 0.686
R7349 G.n5711 G.n5710 0.686
R7350 G.n5677 G.n5676 0.686
R7351 G.n5646 G.n5645 0.686
R7352 G.n5615 G.n5614 0.686
R7353 G.n5587 G.n5586 0.686
R7354 G.n5562 G.n5561 0.686
R7355 G.n5537 G.n5536 0.686
R7356 G.n5324 G.n5323 0.686
R7357 G.n5326 G.n5325 0.686
R7358 G.n5328 G.n5327 0.686
R7359 G.n5330 G.n5329 0.686
R7360 G.n5332 G.n5331 0.686
R7361 G.n5334 G.n5333 0.686
R7362 G.n5336 G.n5335 0.686
R7363 G.n5338 G.n5337 0.686
R7364 G.n5340 G.n5339 0.686
R7365 G.n5342 G.n5341 0.686
R7366 G.n5365 G.n5364 0.686
R7367 G.n5363 G.n5362 0.686
R7368 G.n5361 G.n5360 0.686
R7369 G.n5359 G.n5358 0.686
R7370 G.n5357 G.n5356 0.686
R7371 G.n5355 G.n5354 0.686
R7372 G.n5353 G.n5352 0.686
R7373 G.n3428 G.n3427 0.686
R7374 G.n3430 G.n3429 0.686
R7375 G.n3432 G.n3431 0.686
R7376 G.n3434 G.n3433 0.686
R7377 G.n3436 G.n3435 0.686
R7378 G.n3447 G.n3446 0.686
R7379 G.n3445 G.n3444 0.686
R7380 G.n3443 G.n3442 0.686
R7381 G.n6761 G.n6760 0.686
R7382 G.n6743 G.n6742 0.686
R7383 G.n6722 G.n6721 0.686
R7384 G.n6698 G.n6697 0.686
R7385 G.n6671 G.n6670 0.686
R7386 G.n6641 G.n6640 0.686
R7387 G.n6608 G.n6607 0.686
R7388 G.n6571 G.n6570 0.686
R7389 G.n6530 G.n6529 0.686
R7390 G.n6486 G.n6485 0.686
R7391 G.n6438 G.n6437 0.686
R7392 G.n6387 G.n6386 0.686
R7393 G.n6334 G.n6333 0.686
R7394 G.n6280 G.n6279 0.686
R7395 G.n6226 G.n6225 0.686
R7396 G.n6172 G.n6171 0.686
R7397 G.n6118 G.n6117 0.686
R7398 G.n6066 G.n6065 0.686
R7399 G.n6015 G.n6014 0.686
R7400 G.n5966 G.n5965 0.686
R7401 G.n5920 G.n5919 0.686
R7402 G.n5875 G.n5874 0.686
R7403 G.n5832 G.n5831 0.686
R7404 G.n5792 G.n5791 0.686
R7405 G.n5753 G.n5752 0.686
R7406 G.n5716 G.n5715 0.686
R7407 G.n5682 G.n5681 0.686
R7408 G.n5651 G.n5650 0.686
R7409 G.n5620 G.n5619 0.686
R7410 G.n5592 G.n5591 0.686
R7411 G.n5567 G.n5566 0.686
R7412 G.n5542 G.n5541 0.686
R7413 G.n5520 G.n5519 0.686
R7414 G.n5501 G.n5500 0.686
R7415 G.n5483 G.n5482 0.686
R7416 G.n5375 G.n5374 0.686
R7417 G.n5377 G.n5376 0.686
R7418 G.n5379 G.n5378 0.686
R7419 G.n5381 G.n5380 0.686
R7420 G.n5383 G.n5382 0.686
R7421 G.n5385 G.n5384 0.686
R7422 G.n5387 G.n5386 0.686
R7423 G.n5400 G.n5399 0.686
R7424 G.n5397 G.n5396 0.686
R7425 G.n5394 G.n5393 0.686
R7426 G.n5391 G.n5390 0.686
R7427 G.n3453 G.n3452 0.686
R7428 G.n3455 G.n3454 0.686
R7429 G.n3457 G.n3456 0.686
R7430 G.n3463 G.n3462 0.686
R7431 G.n3462 G.n3460 0.686
R7432 G.n6780 G.n6773 0.686
R7433 G.n6765 G.n6755 0.686
R7434 G.n6747 G.n6734 0.686
R7435 G.n6726 G.n6710 0.686
R7436 G.n6702 G.n6683 0.686
R7437 G.n6675 G.n6653 0.686
R7438 G.n6645 G.n6620 0.686
R7439 G.n6612 G.n6583 0.686
R7440 G.n6575 G.n6542 0.686
R7441 G.n6534 G.n6498 0.686
R7442 G.n6490 G.n6450 0.686
R7443 G.n6442 G.n6399 0.686
R7444 G.n6391 G.n6346 0.686
R7445 G.n6338 G.n6292 0.686
R7446 G.n6284 G.n6238 0.686
R7447 G.n6230 G.n6184 0.686
R7448 G.n6176 G.n6130 0.686
R7449 G.n6122 G.n6078 0.686
R7450 G.n6070 G.n6027 0.686
R7451 G.n6019 G.n5978 0.686
R7452 G.n5970 G.n5932 0.686
R7453 G.n5924 G.n5887 0.686
R7454 G.n5879 G.n5844 0.686
R7455 G.n5836 G.n5804 0.686
R7456 G.n5796 G.n5765 0.686
R7457 G.n5757 G.n5728 0.686
R7458 G.n5720 G.n5694 0.686
R7459 G.n5686 G.n5663 0.686
R7460 G.n5655 G.n5632 0.686
R7461 G.n5624 G.n5604 0.686
R7462 G.n5596 G.n5579 0.686
R7463 G.n5571 G.n5554 0.686
R7464 G.n5546 G.n5532 0.686
R7465 G.n5524 G.n5513 0.686
R7466 G.n5505 G.n5495 0.686
R7467 G.n5487 G.n5479 0.686
R7468 G.n5471 G.n5466 0.686
R7469 G.n5458 G.n5454 0.686
R7470 G.n5446 G.n5444 0.686
R7471 G.n5406 G.n5405 0.686
R7472 G.n5409 G.n5407 0.686
R7473 G.n5410 G.n5409 0.686
R7474 G.n5414 G.n5412 0.686
R7475 G.n3464 G.n3463 0.686
R7476 G.n6792 G.n6791 0.686
R7477 G.n5407 G.n5406 0.686
R7478 G.n5411 G.n5410 0.686
R7479 G.n5412 G.n5411 0.686
R7480 G.n6803 G.n6799 0.686
R7481 G.n6794 G.n6787 0.686
R7482 G.n6782 G.n6772 0.686
R7483 G.n6767 G.n6754 0.686
R7484 G.n6749 G.n6733 0.686
R7485 G.n6728 G.n6709 0.686
R7486 G.n6704 G.n6682 0.686
R7487 G.n6677 G.n6652 0.686
R7488 G.n6647 G.n6619 0.686
R7489 G.n6614 G.n6582 0.686
R7490 G.n6577 G.n6541 0.686
R7491 G.n6536 G.n6497 0.686
R7492 G.n6492 G.n6449 0.686
R7493 G.n6444 G.n6398 0.686
R7494 G.n6393 G.n6345 0.686
R7495 G.n6340 G.n6291 0.686
R7496 G.n6286 G.n6237 0.686
R7497 G.n6232 G.n6183 0.686
R7498 G.n6178 G.n6129 0.686
R7499 G.n6124 G.n6077 0.686
R7500 G.n6072 G.n6026 0.686
R7501 G.n6021 G.n5977 0.686
R7502 G.n5972 G.n5931 0.686
R7503 G.n5926 G.n5886 0.686
R7504 G.n5881 G.n5843 0.686
R7505 G.n5838 G.n5803 0.686
R7506 G.n5798 G.n5764 0.686
R7507 G.n5759 G.n5727 0.686
R7508 G.n5722 G.n5693 0.686
R7509 G.n5688 G.n5662 0.686
R7510 G.n5657 G.n5631 0.686
R7511 G.n5626 G.n5603 0.686
R7512 G.n5598 G.n5578 0.686
R7513 G.n5573 G.n5553 0.686
R7514 G.n5548 G.n5531 0.686
R7515 G.n5526 G.n5512 0.686
R7516 G.n5507 G.n5494 0.686
R7517 G.n5489 G.n5478 0.686
R7518 G.n5473 G.n5465 0.686
R7519 G.n5460 G.n5453 0.686
R7520 G.n5448 G.n5443 0.686
R7521 G.n5438 G.n5436 0.686
R7522 G.n5431 G.n5430 0.686
R7523 G.n5418 G.n5417 0.686
R7524 G.n5420 G.n5419 0.686
R7525 G.n6811 G.n6810 0.686
R7526 G.n6806 G.n6805 0.686
R7527 G.n6797 G.n6796 0.686
R7528 G.n6785 G.n6784 0.686
R7529 G.n6770 G.n6769 0.686
R7530 G.n6752 G.n6751 0.686
R7531 G.n6731 G.n6730 0.686
R7532 G.n6707 G.n6706 0.686
R7533 G.n6680 G.n6679 0.686
R7534 G.n6650 G.n6649 0.686
R7535 G.n6617 G.n6616 0.686
R7536 G.n6580 G.n6579 0.686
R7537 G.n6539 G.n6538 0.686
R7538 G.n6495 G.n6494 0.686
R7539 G.n6447 G.n6446 0.686
R7540 G.n6396 G.n6395 0.686
R7541 G.n6343 G.n6342 0.686
R7542 G.n6289 G.n6288 0.686
R7543 G.n6235 G.n6234 0.686
R7544 G.n6181 G.n6180 0.686
R7545 G.n6127 G.n6126 0.686
R7546 G.n6075 G.n6074 0.686
R7547 G.n6024 G.n6023 0.686
R7548 G.n5975 G.n5974 0.686
R7549 G.n5929 G.n5928 0.686
R7550 G.n5884 G.n5883 0.686
R7551 G.n5841 G.n5840 0.686
R7552 G.n5801 G.n5800 0.686
R7553 G.n5762 G.n5761 0.686
R7554 G.n5725 G.n5724 0.686
R7555 G.n5691 G.n5690 0.686
R7556 G.n5660 G.n5659 0.686
R7557 G.n5629 G.n5628 0.686
R7558 G.n5601 G.n5600 0.686
R7559 G.n5576 G.n5575 0.686
R7560 G.n5551 G.n5550 0.686
R7561 G.n5529 G.n5528 0.686
R7562 G.n5510 G.n5509 0.686
R7563 G.n5492 G.n5491 0.686
R7564 G.n5476 G.n5475 0.686
R7565 G.n5463 G.n5462 0.686
R7566 G.n5451 G.n5450 0.686
R7567 G.n5441 G.n5440 0.686
R7568 G.n5434 G.n5433 0.686
R7569 G.n5428 G.n5427 0.686
R7570 G.n5423 G.n5422 0.686
R7571 G.n5419 G.n5418 0.686
R7572 G.n3468 G.n3467 0.686
R7573 G.n3458 G.n3457 0.655
R7574 G.n5403 G.n5402 0.655
R7575 G.n3475 G.n3449 0.655
R7576 G.n5388 G.n5387 0.655
R7577 G.n3437 G.n3436 0.655
R7578 G.n5367 G.n5366 0.655
R7579 G.n3477 G.n3422 0.655
R7580 G.n5343 G.n5342 0.655
R7581 G.n3404 G.n3403 0.655
R7582 G.n5313 G.n5312 0.655
R7583 G.n3479 G.n3383 0.655
R7584 G.n5280 G.n5279 0.655
R7585 G.n3359 G.n3358 0.655
R7586 G.n5242 G.n5241 0.655
R7587 G.n3481 G.n3332 0.655
R7588 G.n5200 G.n5199 0.655
R7589 G.n3302 G.n3301 0.655
R7590 G.n5153 G.n5152 0.655
R7591 G.n3483 G.n3270 0.655
R7592 G.n5102 G.n5101 0.655
R7593 G.n3235 G.n3234 0.655
R7594 G.n5048 G.n5047 0.655
R7595 G.n3485 G.n3198 0.655
R7596 G.n4988 G.n4987 0.655
R7597 G.n3158 G.n3157 0.655
R7598 G.n4925 G.n4924 0.655
R7599 G.n3487 G.n3115 0.655
R7600 G.n4856 G.n4855 0.655
R7601 G.n3070 G.n3069 0.655
R7602 G.n4784 G.n4783 0.655
R7603 G.n3489 G.n3022 0.655
R7604 G.n4706 G.n4705 0.655
R7605 G.n2973 G.n2972 0.655
R7606 G.n4630 G.n4629 0.655
R7607 G.n3491 G.n2927 0.655
R7608 G.n4557 G.n4556 0.655
R7609 G.n2881 G.n2880 0.655
R7610 G.n4487 G.n4486 0.655
R7611 G.n3493 G.n2838 0.655
R7612 G.n4417 G.n4416 0.655
R7613 G.n2796 G.n2795 0.655
R7614 G.n4350 G.n4349 0.655
R7615 G.n3495 G.n2756 0.655
R7616 G.n4286 G.n4285 0.655
R7617 G.n2719 G.n2718 0.655
R7618 G.n4225 G.n4224 0.655
R7619 G.n3497 G.n2682 0.655
R7620 G.n4167 G.n4166 0.655
R7621 G.n2648 G.n2647 0.655
R7622 G.n4112 G.n4111 0.655
R7623 G.n3499 G.n2614 0.655
R7624 G.n4060 G.n4059 0.655
R7625 G.n2583 G.n2582 0.655
R7626 G.n4011 G.n4010 0.655
R7627 G.n3501 G.n2553 0.655
R7628 G.n3965 G.n3964 0.655
R7629 G.n2525 G.n2524 0.655
R7630 G.n3919 G.n3918 0.655
R7631 G.n3503 G.n2498 0.655
R7632 G.n3876 G.n3875 0.655
R7633 G.n2473 G.n2472 0.655
R7634 G.n3836 G.n3835 0.655
R7635 G.n3505 G.n2451 0.655
R7636 G.n3799 G.n3798 0.655
R7637 G.n2429 G.n2428 0.655
R7638 G.n3765 G.n3764 0.655
R7639 G.n3507 G.n2410 0.655
R7640 G.n3734 G.n3733 0.655
R7641 G.n2391 G.n2390 0.655
R7642 G.n3706 G.n3705 0.655
R7643 G.n3509 G.n2375 0.655
R7644 G.n3681 G.n3680 0.655
R7645 G.n2360 G.n2359 0.655
R7646 G.n3656 G.n3655 0.655
R7647 G.n3511 G.n2347 0.655
R7648 G.n3634 G.n3633 0.655
R7649 G.n2337 G.n2336 0.655
R7650 G.n3615 G.n3614 0.655
R7651 G.n3513 G.n2327 0.655
R7652 G.n3599 G.n3598 0.655
R7653 G.n2320 G.n2319 0.655
R7654 G.n3586 G.n3585 0.655
R7655 G.n3515 G.n2313 0.655
R7656 G.n3576 G.n3575 0.655
R7657 G.n2309 G.n2308 0.655
R7658 G.n3569 G.n3568 0.655
R7659 G.n3517 G.n2306 0.655
R7660 G.n6908 G.n3565 0.655
R7661 G.n6907 G.n3569 0.655
R7662 G.n3516 G.n2309 0.655
R7663 G.n2313 G.n2312 0.655
R7664 G.n6906 G.n3576 0.655
R7665 G.n6905 G.n3586 0.655
R7666 G.n3514 G.n2320 0.655
R7667 G.n2327 G.n2326 0.655
R7668 G.n6904 G.n3599 0.655
R7669 G.n6903 G.n3615 0.655
R7670 G.n3512 G.n2337 0.655
R7671 G.n2347 G.n2346 0.655
R7672 G.n6902 G.n3634 0.655
R7673 G.n6901 G.n3656 0.655
R7674 G.n3510 G.n2360 0.655
R7675 G.n2375 G.n2374 0.655
R7676 G.n6900 G.n3681 0.655
R7677 G.n6899 G.n3706 0.655
R7678 G.n3508 G.n2391 0.655
R7679 G.n2410 G.n2409 0.655
R7680 G.n6898 G.n3734 0.655
R7681 G.n6897 G.n3765 0.655
R7682 G.n3506 G.n2429 0.655
R7683 G.n2451 G.n2450 0.655
R7684 G.n6896 G.n3799 0.655
R7685 G.n6895 G.n3836 0.655
R7686 G.n3504 G.n2473 0.655
R7687 G.n2498 G.n2497 0.655
R7688 G.n6894 G.n3876 0.655
R7689 G.n6893 G.n3919 0.655
R7690 G.n3502 G.n2525 0.655
R7691 G.n2553 G.n2552 0.655
R7692 G.n6892 G.n3965 0.655
R7693 G.n6891 G.n4011 0.655
R7694 G.n3500 G.n2583 0.655
R7695 G.n2614 G.n2613 0.655
R7696 G.n6890 G.n4060 0.655
R7697 G.n6889 G.n4112 0.655
R7698 G.n3498 G.n2648 0.655
R7699 G.n2682 G.n2681 0.655
R7700 G.n6888 G.n4167 0.655
R7701 G.n6887 G.n4225 0.655
R7702 G.n3496 G.n2719 0.655
R7703 G.n2756 G.n2755 0.655
R7704 G.n6886 G.n4286 0.655
R7705 G.n6885 G.n4350 0.655
R7706 G.n3494 G.n2796 0.655
R7707 G.n2838 G.n2837 0.655
R7708 G.n6884 G.n4417 0.655
R7709 G.n6883 G.n4487 0.655
R7710 G.n3492 G.n2881 0.655
R7711 G.n2927 G.n2926 0.655
R7712 G.n6882 G.n4557 0.655
R7713 G.n6881 G.n4630 0.655
R7714 G.n3490 G.n2973 0.655
R7715 G.n3022 G.n3021 0.655
R7716 G.n6880 G.n4706 0.655
R7717 G.n6879 G.n4784 0.655
R7718 G.n3488 G.n3070 0.655
R7719 G.n3115 G.n3114 0.655
R7720 G.n6878 G.n4856 0.655
R7721 G.n6877 G.n4925 0.655
R7722 G.n3486 G.n3158 0.655
R7723 G.n3198 G.n3197 0.655
R7724 G.n6876 G.n4988 0.655
R7725 G.n6875 G.n5048 0.655
R7726 G.n3484 G.n3235 0.655
R7727 G.n3270 G.n3269 0.655
R7728 G.n6874 G.n5102 0.655
R7729 G.n6873 G.n5153 0.655
R7730 G.n3482 G.n3302 0.655
R7731 G.n3332 G.n3331 0.655
R7732 G.n6872 G.n5200 0.655
R7733 G.n6871 G.n5242 0.655
R7734 G.n3480 G.n3359 0.655
R7735 G.n3383 G.n3382 0.655
R7736 G.n6870 G.n5280 0.655
R7737 G.n6869 G.n5313 0.655
R7738 G.n3478 G.n3404 0.655
R7739 G.n3422 G.n3421 0.655
R7740 G.n6868 G.n5343 0.655
R7741 G.n6867 G.n5367 0.655
R7742 G.n3476 G.n3437 0.655
R7743 G.n3449 G.n3448 0.655
R7744 G.n6866 G.n5388 0.655
R7745 G.n5415 G.n5414 0.655
R7746 G.n6865 G.n5403 0.655
R7747 G.n3474 G.n3458 0.655
R7748 G.n3465 G.n3464 0.655
R7749 G.n3473 G.n3465 0.655
R7750 G.n6864 G.n5415 0.655
R7751 G.n3469 G.n3468 0.655
R7752 G.n5421 G.n5420 0.655
R7753 G.n3471 G.n3470 0.655
R7754 G.n5424 G.n5423 0.655
R7755 G.n6862 G.n5424 0.655
R7756 G.n6863 G.n5421 0.655
R7757 G.n3472 G.n3469 0.655
R7758 G.n6862 G.n6861 0.645
R7759 G.n3518 G.n3517 0.644
R7760 G.n3468 G.n3466 0.624
R7761 G.n5420 G.n5416 0.624
R7762 G.n6861 G.n5425 0.624
R7763 G.n6860 G.n5429 0.624
R7764 G.n5432 G.n5431 0.624
R7765 G.n6859 G.n5435 0.624
R7766 G.n5439 G.n5438 0.624
R7767 G.n6858 G.n5442 0.624
R7768 G.n5449 G.n5448 0.624
R7769 G.n6857 G.n5452 0.624
R7770 G.n5461 G.n5460 0.624
R7771 G.n6856 G.n5464 0.624
R7772 G.n5474 G.n5473 0.624
R7773 G.n6855 G.n5477 0.624
R7774 G.n5490 G.n5489 0.624
R7775 G.n6854 G.n5493 0.624
R7776 G.n5508 G.n5507 0.624
R7777 G.n6853 G.n5511 0.624
R7778 G.n5527 G.n5526 0.624
R7779 G.n6852 G.n5530 0.624
R7780 G.n5549 G.n5548 0.624
R7781 G.n6851 G.n5552 0.624
R7782 G.n5574 G.n5573 0.624
R7783 G.n6850 G.n5577 0.624
R7784 G.n5599 G.n5598 0.624
R7785 G.n6849 G.n5602 0.624
R7786 G.n5627 G.n5626 0.624
R7787 G.n6848 G.n5630 0.624
R7788 G.n5658 G.n5657 0.624
R7789 G.n6847 G.n5661 0.624
R7790 G.n5689 G.n5688 0.624
R7791 G.n6846 G.n5692 0.624
R7792 G.n5723 G.n5722 0.624
R7793 G.n6845 G.n5726 0.624
R7794 G.n5760 G.n5759 0.624
R7795 G.n6844 G.n5763 0.624
R7796 G.n5799 G.n5798 0.624
R7797 G.n6843 G.n5802 0.624
R7798 G.n5839 G.n5838 0.624
R7799 G.n6842 G.n5842 0.624
R7800 G.n5882 G.n5881 0.624
R7801 G.n6841 G.n5885 0.624
R7802 G.n5927 G.n5926 0.624
R7803 G.n6840 G.n5930 0.624
R7804 G.n5973 G.n5972 0.624
R7805 G.n6839 G.n5976 0.624
R7806 G.n6022 G.n6021 0.624
R7807 G.n6838 G.n6025 0.624
R7808 G.n6073 G.n6072 0.624
R7809 G.n6837 G.n6076 0.624
R7810 G.n6125 G.n6124 0.624
R7811 G.n6836 G.n6128 0.624
R7812 G.n6179 G.n6178 0.624
R7813 G.n6835 G.n6182 0.624
R7814 G.n6233 G.n6232 0.624
R7815 G.n6834 G.n6236 0.624
R7816 G.n6287 G.n6286 0.624
R7817 G.n6833 G.n6290 0.624
R7818 G.n6341 G.n6340 0.624
R7819 G.n6832 G.n6344 0.624
R7820 G.n6394 G.n6393 0.624
R7821 G.n6831 G.n6397 0.624
R7822 G.n6445 G.n6444 0.624
R7823 G.n6830 G.n6448 0.624
R7824 G.n6493 G.n6492 0.624
R7825 G.n6829 G.n6496 0.624
R7826 G.n6537 G.n6536 0.624
R7827 G.n6828 G.n6540 0.624
R7828 G.n6578 G.n6577 0.624
R7829 G.n6827 G.n6581 0.624
R7830 G.n6615 G.n6614 0.624
R7831 G.n6826 G.n6618 0.624
R7832 G.n6648 G.n6647 0.624
R7833 G.n6825 G.n6651 0.624
R7834 G.n6678 G.n6677 0.624
R7835 G.n6824 G.n6681 0.624
R7836 G.n6705 G.n6704 0.624
R7837 G.n6823 G.n6708 0.624
R7838 G.n6729 G.n6728 0.624
R7839 G.n6822 G.n6732 0.624
R7840 G.n6750 G.n6749 0.624
R7841 G.n6821 G.n6753 0.624
R7842 G.n6768 G.n6767 0.624
R7843 G.n6820 G.n6771 0.624
R7844 G.n6783 G.n6782 0.624
R7845 G.n6819 G.n6786 0.624
R7846 G.n6795 G.n6794 0.624
R7847 G.n6818 G.n6798 0.624
R7848 G.n6804 G.n6803 0.624
R7849 G.n6817 G.n6807 0.624
R7850 G.n6809 G.n6808 0.624
R7851 G.n6816 G.n6812 0.624
R7852 G.n6812 G.n6811 0.624
R7853 G.n6814 G.n6813 0.624
R7854 G.n6807 G.n6806 0.624
R7855 G.n6798 G.n6797 0.624
R7856 G.n6786 G.n6785 0.624
R7857 G.n6771 G.n6770 0.624
R7858 G.n6753 G.n6752 0.624
R7859 G.n6732 G.n6731 0.624
R7860 G.n6708 G.n6707 0.624
R7861 G.n6681 G.n6680 0.624
R7862 G.n6651 G.n6650 0.624
R7863 G.n6618 G.n6617 0.624
R7864 G.n6581 G.n6580 0.624
R7865 G.n6540 G.n6539 0.624
R7866 G.n6496 G.n6495 0.624
R7867 G.n6448 G.n6447 0.624
R7868 G.n6397 G.n6396 0.624
R7869 G.n6344 G.n6343 0.624
R7870 G.n6290 G.n6289 0.624
R7871 G.n6236 G.n6235 0.624
R7872 G.n6182 G.n6181 0.624
R7873 G.n6128 G.n6127 0.624
R7874 G.n6076 G.n6075 0.624
R7875 G.n6025 G.n6024 0.624
R7876 G.n5976 G.n5975 0.624
R7877 G.n5930 G.n5929 0.624
R7878 G.n5885 G.n5884 0.624
R7879 G.n5842 G.n5841 0.624
R7880 G.n5802 G.n5801 0.624
R7881 G.n5763 G.n5762 0.624
R7882 G.n5726 G.n5725 0.624
R7883 G.n5692 G.n5691 0.624
R7884 G.n5661 G.n5660 0.624
R7885 G.n5630 G.n5629 0.624
R7886 G.n5602 G.n5601 0.624
R7887 G.n5577 G.n5576 0.624
R7888 G.n5552 G.n5551 0.624
R7889 G.n5530 G.n5529 0.624
R7890 G.n5511 G.n5510 0.624
R7891 G.n5493 G.n5492 0.624
R7892 G.n5477 G.n5476 0.624
R7893 G.n5464 G.n5463 0.624
R7894 G.n5452 G.n5451 0.624
R7895 G.n5442 G.n5441 0.624
R7896 G.n5435 G.n5434 0.624
R7897 G.n5429 G.n5428 0.624
R7898 G.n6811 G.n6809 0.624
R7899 G.n6806 G.n6804 0.624
R7900 G.n6797 G.n6795 0.624
R7901 G.n6785 G.n6783 0.624
R7902 G.n6770 G.n6768 0.624
R7903 G.n6752 G.n6750 0.624
R7904 G.n6731 G.n6729 0.624
R7905 G.n6707 G.n6705 0.624
R7906 G.n6680 G.n6678 0.624
R7907 G.n6650 G.n6648 0.624
R7908 G.n6617 G.n6615 0.624
R7909 G.n6580 G.n6578 0.624
R7910 G.n6539 G.n6537 0.624
R7911 G.n6495 G.n6493 0.624
R7912 G.n6447 G.n6445 0.624
R7913 G.n6396 G.n6394 0.624
R7914 G.n6343 G.n6341 0.624
R7915 G.n6289 G.n6287 0.624
R7916 G.n6235 G.n6233 0.624
R7917 G.n6181 G.n6179 0.624
R7918 G.n6127 G.n6125 0.624
R7919 G.n6075 G.n6073 0.624
R7920 G.n6024 G.n6022 0.624
R7921 G.n5975 G.n5973 0.624
R7922 G.n5929 G.n5927 0.624
R7923 G.n5884 G.n5882 0.624
R7924 G.n5841 G.n5839 0.624
R7925 G.n5801 G.n5799 0.624
R7926 G.n5762 G.n5760 0.624
R7927 G.n5725 G.n5723 0.624
R7928 G.n5691 G.n5689 0.624
R7929 G.n5660 G.n5658 0.624
R7930 G.n5629 G.n5627 0.624
R7931 G.n5601 G.n5599 0.624
R7932 G.n5576 G.n5574 0.624
R7933 G.n5551 G.n5549 0.624
R7934 G.n5529 G.n5527 0.624
R7935 G.n5510 G.n5508 0.624
R7936 G.n5492 G.n5490 0.624
R7937 G.n5476 G.n5474 0.624
R7938 G.n5463 G.n5461 0.624
R7939 G.n5451 G.n5449 0.624
R7940 G.n5441 G.n5439 0.624
R7941 G.n5434 G.n5432 0.624
R7942 G.n6794 G.n6793 0.624
R7943 G.n6782 G.n6781 0.624
R7944 G.n6767 G.n6766 0.624
R7945 G.n6749 G.n6748 0.624
R7946 G.n6728 G.n6727 0.624
R7947 G.n6704 G.n6703 0.624
R7948 G.n6677 G.n6676 0.624
R7949 G.n6647 G.n6646 0.624
R7950 G.n6614 G.n6613 0.624
R7951 G.n6577 G.n6576 0.624
R7952 G.n6536 G.n6535 0.624
R7953 G.n6492 G.n6491 0.624
R7954 G.n6444 G.n6443 0.624
R7955 G.n6393 G.n6392 0.624
R7956 G.n6340 G.n6339 0.624
R7957 G.n6286 G.n6285 0.624
R7958 G.n6232 G.n6231 0.624
R7959 G.n6178 G.n6177 0.624
R7960 G.n6124 G.n6123 0.624
R7961 G.n6072 G.n6071 0.624
R7962 G.n6021 G.n6020 0.624
R7963 G.n5972 G.n5971 0.624
R7964 G.n5926 G.n5925 0.624
R7965 G.n5881 G.n5880 0.624
R7966 G.n5838 G.n5837 0.624
R7967 G.n5798 G.n5797 0.624
R7968 G.n5759 G.n5758 0.624
R7969 G.n5722 G.n5721 0.624
R7970 G.n5688 G.n5687 0.624
R7971 G.n5657 G.n5656 0.624
R7972 G.n5626 G.n5625 0.624
R7973 G.n5598 G.n5597 0.624
R7974 G.n5573 G.n5572 0.624
R7975 G.n5548 G.n5547 0.624
R7976 G.n5526 G.n5525 0.624
R7977 G.n5507 G.n5506 0.624
R7978 G.n5489 G.n5488 0.624
R7979 G.n5473 G.n5472 0.624
R7980 G.n5460 G.n5459 0.624
R7981 G.n5448 G.n5447 0.624
R7982 G.n5438 G.n5437 0.624
R7983 G.n6803 G.n6802 0.624
R7984 G.n5414 G.n5413 0.624
R7985 G.n5411 G.n5404 0.624
R7986 G.n5409 G.n5408 0.624
R7987 G.n5447 G.n5446 0.624
R7988 G.n5459 G.n5458 0.624
R7989 G.n5472 G.n5471 0.624
R7990 G.n5488 G.n5487 0.624
R7991 G.n5506 G.n5505 0.624
R7992 G.n5525 G.n5524 0.624
R7993 G.n5547 G.n5546 0.624
R7994 G.n5572 G.n5571 0.624
R7995 G.n5597 G.n5596 0.624
R7996 G.n5625 G.n5624 0.624
R7997 G.n5656 G.n5655 0.624
R7998 G.n5687 G.n5686 0.624
R7999 G.n5721 G.n5720 0.624
R8000 G.n5758 G.n5757 0.624
R8001 G.n5797 G.n5796 0.624
R8002 G.n5837 G.n5836 0.624
R8003 G.n5880 G.n5879 0.624
R8004 G.n5925 G.n5924 0.624
R8005 G.n5971 G.n5970 0.624
R8006 G.n6020 G.n6019 0.624
R8007 G.n6071 G.n6070 0.624
R8008 G.n6123 G.n6122 0.624
R8009 G.n6177 G.n6176 0.624
R8010 G.n6231 G.n6230 0.624
R8011 G.n6285 G.n6284 0.624
R8012 G.n6339 G.n6338 0.624
R8013 G.n6392 G.n6391 0.624
R8014 G.n6443 G.n6442 0.624
R8015 G.n6491 G.n6490 0.624
R8016 G.n6535 G.n6534 0.624
R8017 G.n6576 G.n6575 0.624
R8018 G.n6613 G.n6612 0.624
R8019 G.n6646 G.n6645 0.624
R8020 G.n6676 G.n6675 0.624
R8021 G.n6703 G.n6702 0.624
R8022 G.n6727 G.n6726 0.624
R8023 G.n6748 G.n6747 0.624
R8024 G.n6766 G.n6765 0.624
R8025 G.n6781 G.n6780 0.624
R8026 G.n6793 G.n6792 0.624
R8027 G.n6802 G.n6801 0.624
R8028 G.n3462 G.n3461 0.624
R8029 G.n3464 G.n3459 0.624
R8030 G.n6801 G.n6800 0.624
R8031 G.n6792 G.n6790 0.624
R8032 G.n6780 G.n6779 0.624
R8033 G.n6765 G.n6764 0.624
R8034 G.n6747 G.n6746 0.624
R8035 G.n6726 G.n6725 0.624
R8036 G.n6702 G.n6701 0.624
R8037 G.n6675 G.n6674 0.624
R8038 G.n6645 G.n6644 0.624
R8039 G.n6612 G.n6611 0.624
R8040 G.n6575 G.n6574 0.624
R8041 G.n6534 G.n6533 0.624
R8042 G.n6490 G.n6489 0.624
R8043 G.n6442 G.n6441 0.624
R8044 G.n6391 G.n6390 0.624
R8045 G.n6338 G.n6337 0.624
R8046 G.n6284 G.n6283 0.624
R8047 G.n6230 G.n6229 0.624
R8048 G.n6176 G.n6175 0.624
R8049 G.n6122 G.n6121 0.624
R8050 G.n6070 G.n6069 0.624
R8051 G.n6019 G.n6018 0.624
R8052 G.n5970 G.n5969 0.624
R8053 G.n5924 G.n5923 0.624
R8054 G.n5879 G.n5878 0.624
R8055 G.n5836 G.n5835 0.624
R8056 G.n5796 G.n5795 0.624
R8057 G.n5757 G.n5756 0.624
R8058 G.n5720 G.n5719 0.624
R8059 G.n5686 G.n5685 0.624
R8060 G.n5655 G.n5654 0.624
R8061 G.n5624 G.n5623 0.624
R8062 G.n5596 G.n5595 0.624
R8063 G.n5571 G.n5570 0.624
R8064 G.n5546 G.n5545 0.624
R8065 G.n5524 G.n5523 0.624
R8066 G.n5505 G.n5504 0.624
R8067 G.n5487 G.n5486 0.624
R8068 G.n5471 G.n5470 0.624
R8069 G.n5458 G.n5457 0.624
R8070 G.n5446 G.n5445 0.624
R8071 G.n5387 G.n5368 0.624
R8072 G.n5385 G.n5369 0.624
R8073 G.n5383 G.n5370 0.624
R8074 G.n5381 G.n5371 0.624
R8075 G.n5379 G.n5372 0.624
R8076 G.n5377 G.n5373 0.624
R8077 G.n5484 G.n5483 0.624
R8078 G.n5502 G.n5501 0.624
R8079 G.n5521 G.n5520 0.624
R8080 G.n5543 G.n5542 0.624
R8081 G.n5568 G.n5567 0.624
R8082 G.n5593 G.n5592 0.624
R8083 G.n5621 G.n5620 0.624
R8084 G.n5652 G.n5651 0.624
R8085 G.n5683 G.n5682 0.624
R8086 G.n5717 G.n5716 0.624
R8087 G.n5754 G.n5753 0.624
R8088 G.n5793 G.n5792 0.624
R8089 G.n5833 G.n5832 0.624
R8090 G.n5876 G.n5875 0.624
R8091 G.n5921 G.n5920 0.624
R8092 G.n5967 G.n5966 0.624
R8093 G.n6016 G.n6015 0.624
R8094 G.n6067 G.n6066 0.624
R8095 G.n6119 G.n6118 0.624
R8096 G.n6173 G.n6172 0.624
R8097 G.n6227 G.n6226 0.624
R8098 G.n6281 G.n6280 0.624
R8099 G.n6335 G.n6334 0.624
R8100 G.n6388 G.n6387 0.624
R8101 G.n6439 G.n6438 0.624
R8102 G.n6487 G.n6486 0.624
R8103 G.n6531 G.n6530 0.624
R8104 G.n6572 G.n6571 0.624
R8105 G.n6609 G.n6608 0.624
R8106 G.n6642 G.n6641 0.624
R8107 G.n6672 G.n6671 0.624
R8108 G.n6699 G.n6698 0.624
R8109 G.n6723 G.n6722 0.624
R8110 G.n6744 G.n6743 0.624
R8111 G.n6762 G.n6761 0.624
R8112 G.n6777 G.n6776 0.624
R8113 G.n3444 G.n3440 0.624
R8114 G.n3446 G.n3439 0.624
R8115 G.n3448 G.n3438 0.624
R8116 G.n3436 G.n3423 0.624
R8117 G.n3434 G.n3424 0.624
R8118 G.n3432 G.n3425 0.624
R8119 G.n3430 G.n3426 0.624
R8120 G.n6759 G.n6758 0.624
R8121 G.n6741 G.n6740 0.624
R8122 G.n6720 G.n6719 0.624
R8123 G.n6696 G.n6695 0.624
R8124 G.n6669 G.n6668 0.624
R8125 G.n6639 G.n6638 0.624
R8126 G.n6606 G.n6605 0.624
R8127 G.n6569 G.n6568 0.624
R8128 G.n6528 G.n6527 0.624
R8129 G.n6484 G.n6483 0.624
R8130 G.n6436 G.n6435 0.624
R8131 G.n6385 G.n6384 0.624
R8132 G.n6332 G.n6331 0.624
R8133 G.n6278 G.n6277 0.624
R8134 G.n6224 G.n6223 0.624
R8135 G.n6170 G.n6169 0.624
R8136 G.n6116 G.n6115 0.624
R8137 G.n6064 G.n6063 0.624
R8138 G.n6013 G.n6012 0.624
R8139 G.n5964 G.n5963 0.624
R8140 G.n5918 G.n5917 0.624
R8141 G.n5873 G.n5872 0.624
R8142 G.n5830 G.n5829 0.624
R8143 G.n5790 G.n5789 0.624
R8144 G.n5751 G.n5750 0.624
R8145 G.n5714 G.n5713 0.624
R8146 G.n5680 G.n5679 0.624
R8147 G.n5649 G.n5648 0.624
R8148 G.n5618 G.n5617 0.624
R8149 G.n5590 G.n5589 0.624
R8150 G.n5565 G.n5564 0.624
R8151 G.n5540 G.n5539 0.624
R8152 G.n5518 G.n5517 0.624
R8153 G.n5499 G.n5498 0.624
R8154 G.n5354 G.n5350 0.624
R8155 G.n5356 G.n5349 0.624
R8156 G.n5358 G.n5348 0.624
R8157 G.n5360 G.n5347 0.624
R8158 G.n5362 G.n5346 0.624
R8159 G.n5364 G.n5345 0.624
R8160 G.n5366 G.n5344 0.624
R8161 G.n5342 G.n5314 0.624
R8162 G.n5340 G.n5315 0.624
R8163 G.n5338 G.n5316 0.624
R8164 G.n5336 G.n5317 0.624
R8165 G.n5334 G.n5318 0.624
R8166 G.n5332 G.n5319 0.624
R8167 G.n5330 G.n5320 0.624
R8168 G.n5328 G.n5321 0.624
R8169 G.n5326 G.n5322 0.624
R8170 G.n5538 G.n5537 0.624
R8171 G.n5563 G.n5562 0.624
R8172 G.n5588 G.n5587 0.624
R8173 G.n5616 G.n5615 0.624
R8174 G.n5647 G.n5646 0.624
R8175 G.n5678 G.n5677 0.624
R8176 G.n5712 G.n5711 0.624
R8177 G.n5749 G.n5748 0.624
R8178 G.n5788 G.n5787 0.624
R8179 G.n5828 G.n5827 0.624
R8180 G.n5871 G.n5870 0.624
R8181 G.n5916 G.n5915 0.624
R8182 G.n5962 G.n5961 0.624
R8183 G.n6011 G.n6010 0.624
R8184 G.n6062 G.n6061 0.624
R8185 G.n6114 G.n6113 0.624
R8186 G.n6168 G.n6167 0.624
R8187 G.n6222 G.n6221 0.624
R8188 G.n6276 G.n6275 0.624
R8189 G.n6330 G.n6329 0.624
R8190 G.n6383 G.n6382 0.624
R8191 G.n6434 G.n6433 0.624
R8192 G.n6482 G.n6481 0.624
R8193 G.n6526 G.n6525 0.624
R8194 G.n6567 G.n6566 0.624
R8195 G.n6604 G.n6603 0.624
R8196 G.n6637 G.n6636 0.624
R8197 G.n6667 G.n6666 0.624
R8198 G.n6694 G.n6693 0.624
R8199 G.n6718 G.n6717 0.624
R8200 G.n6739 G.n6738 0.624
R8201 G.n3413 G.n3409 0.624
R8202 G.n3415 G.n3408 0.624
R8203 G.n3417 G.n3407 0.624
R8204 G.n3419 G.n3406 0.624
R8205 G.n3421 G.n3405 0.624
R8206 G.n3403 G.n3384 0.624
R8207 G.n3401 G.n3385 0.624
R8208 G.n3399 G.n3386 0.624
R8209 G.n3397 G.n3387 0.624
R8210 G.n3395 G.n3388 0.624
R8211 G.n3393 G.n3389 0.624
R8212 G.n6715 G.n6714 0.624
R8213 G.n6691 G.n6690 0.624
R8214 G.n6664 G.n6663 0.624
R8215 G.n6634 G.n6633 0.624
R8216 G.n6601 G.n6600 0.624
R8217 G.n6564 G.n6563 0.624
R8218 G.n6523 G.n6522 0.624
R8219 G.n6479 G.n6478 0.624
R8220 G.n6431 G.n6430 0.624
R8221 G.n6380 G.n6379 0.624
R8222 G.n6327 G.n6326 0.624
R8223 G.n6273 G.n6272 0.624
R8224 G.n6219 G.n6218 0.624
R8225 G.n6165 G.n6164 0.624
R8226 G.n6111 G.n6110 0.624
R8227 G.n6059 G.n6058 0.624
R8228 G.n6008 G.n6007 0.624
R8229 G.n5959 G.n5958 0.624
R8230 G.n5913 G.n5912 0.624
R8231 G.n5868 G.n5867 0.624
R8232 G.n5825 G.n5824 0.624
R8233 G.n5785 G.n5784 0.624
R8234 G.n5746 G.n5745 0.624
R8235 G.n5709 G.n5708 0.624
R8236 G.n5675 G.n5674 0.624
R8237 G.n5644 G.n5643 0.624
R8238 G.n5613 G.n5612 0.624
R8239 G.n5585 G.n5584 0.624
R8240 G.n5560 G.n5559 0.624
R8241 G.n5294 G.n5290 0.624
R8242 G.n5296 G.n5289 0.624
R8243 G.n5298 G.n5288 0.624
R8244 G.n5300 G.n5287 0.624
R8245 G.n5302 G.n5286 0.624
R8246 G.n5304 G.n5285 0.624
R8247 G.n5306 G.n5284 0.624
R8248 G.n5308 G.n5283 0.624
R8249 G.n5310 G.n5282 0.624
R8250 G.n5312 G.n5281 0.624
R8251 G.n5279 G.n5243 0.624
R8252 G.n5277 G.n5244 0.624
R8253 G.n5275 G.n5245 0.624
R8254 G.n5273 G.n5246 0.624
R8255 G.n5271 G.n5247 0.624
R8256 G.n5269 G.n5248 0.624
R8257 G.n5267 G.n5249 0.624
R8258 G.n5265 G.n5250 0.624
R8259 G.n5263 G.n5251 0.624
R8260 G.n5261 G.n5252 0.624
R8261 G.n5259 G.n5253 0.624
R8262 G.n5611 G.n5610 0.624
R8263 G.n5642 G.n5641 0.624
R8264 G.n5673 G.n5672 0.624
R8265 G.n5707 G.n5706 0.624
R8266 G.n5744 G.n5743 0.624
R8267 G.n5783 G.n5782 0.624
R8268 G.n5823 G.n5822 0.624
R8269 G.n5866 G.n5865 0.624
R8270 G.n5911 G.n5910 0.624
R8271 G.n5957 G.n5956 0.624
R8272 G.n6006 G.n6005 0.624
R8273 G.n6057 G.n6056 0.624
R8274 G.n6109 G.n6108 0.624
R8275 G.n6163 G.n6162 0.624
R8276 G.n6217 G.n6216 0.624
R8277 G.n6271 G.n6270 0.624
R8278 G.n6325 G.n6324 0.624
R8279 G.n6378 G.n6377 0.624
R8280 G.n6429 G.n6428 0.624
R8281 G.n6477 G.n6476 0.624
R8282 G.n6521 G.n6520 0.624
R8283 G.n6562 G.n6561 0.624
R8284 G.n6599 G.n6598 0.624
R8285 G.n6632 G.n6631 0.624
R8286 G.n6662 G.n6661 0.624
R8287 G.n6689 G.n6688 0.624
R8288 G.n3370 G.n3366 0.624
R8289 G.n3372 G.n3365 0.624
R8290 G.n3374 G.n3364 0.624
R8291 G.n3376 G.n3363 0.624
R8292 G.n3378 G.n3362 0.624
R8293 G.n3380 G.n3361 0.624
R8294 G.n3382 G.n3360 0.624
R8295 G.n3358 G.n3333 0.624
R8296 G.n3356 G.n3334 0.624
R8297 G.n3354 G.n3335 0.624
R8298 G.n3352 G.n3336 0.624
R8299 G.n3350 G.n3337 0.624
R8300 G.n3348 G.n3338 0.624
R8301 G.n3346 G.n3339 0.624
R8302 G.n3344 G.n3340 0.624
R8303 G.n6659 G.n6658 0.624
R8304 G.n6629 G.n6628 0.624
R8305 G.n6596 G.n6595 0.624
R8306 G.n6559 G.n6558 0.624
R8307 G.n6518 G.n6517 0.624
R8308 G.n6474 G.n6473 0.624
R8309 G.n6426 G.n6425 0.624
R8310 G.n6375 G.n6374 0.624
R8311 G.n6322 G.n6321 0.624
R8312 G.n6268 G.n6267 0.624
R8313 G.n6214 G.n6213 0.624
R8314 G.n6160 G.n6159 0.624
R8315 G.n6106 G.n6105 0.624
R8316 G.n6054 G.n6053 0.624
R8317 G.n6003 G.n6002 0.624
R8318 G.n5954 G.n5953 0.624
R8319 G.n5908 G.n5907 0.624
R8320 G.n5863 G.n5862 0.624
R8321 G.n5820 G.n5819 0.624
R8322 G.n5780 G.n5779 0.624
R8323 G.n5741 G.n5740 0.624
R8324 G.n5704 G.n5703 0.624
R8325 G.n5670 G.n5669 0.624
R8326 G.n5639 G.n5638 0.624
R8327 G.n5217 G.n5213 0.624
R8328 G.n5219 G.n5212 0.624
R8329 G.n5221 G.n5211 0.624
R8330 G.n5223 G.n5210 0.624
R8331 G.n5225 G.n5209 0.624
R8332 G.n5227 G.n5208 0.624
R8333 G.n5229 G.n5207 0.624
R8334 G.n5231 G.n5206 0.624
R8335 G.n5233 G.n5205 0.624
R8336 G.n5235 G.n5204 0.624
R8337 G.n5237 G.n5203 0.624
R8338 G.n5239 G.n5202 0.624
R8339 G.n5241 G.n5201 0.624
R8340 G.n5199 G.n5154 0.624
R8341 G.n5197 G.n5155 0.624
R8342 G.n5195 G.n5156 0.624
R8343 G.n5193 G.n5157 0.624
R8344 G.n5191 G.n5158 0.624
R8345 G.n5189 G.n5159 0.624
R8346 G.n5187 G.n5160 0.624
R8347 G.n5185 G.n5161 0.624
R8348 G.n5183 G.n5162 0.624
R8349 G.n5181 G.n5163 0.624
R8350 G.n5179 G.n5164 0.624
R8351 G.n5177 G.n5165 0.624
R8352 G.n5175 G.n5166 0.624
R8353 G.n5173 G.n5167 0.624
R8354 G.n5702 G.n5701 0.624
R8355 G.n5739 G.n5738 0.624
R8356 G.n5778 G.n5777 0.624
R8357 G.n5818 G.n5817 0.624
R8358 G.n5861 G.n5860 0.624
R8359 G.n5906 G.n5905 0.624
R8360 G.n5952 G.n5951 0.624
R8361 G.n6001 G.n6000 0.624
R8362 G.n6052 G.n6051 0.624
R8363 G.n6104 G.n6103 0.624
R8364 G.n6158 G.n6157 0.624
R8365 G.n6212 G.n6211 0.624
R8366 G.n6266 G.n6265 0.624
R8367 G.n6320 G.n6319 0.624
R8368 G.n6373 G.n6372 0.624
R8369 G.n6424 G.n6423 0.624
R8370 G.n6472 G.n6471 0.624
R8371 G.n6516 G.n6515 0.624
R8372 G.n6557 G.n6556 0.624
R8373 G.n6594 G.n6593 0.624
R8374 G.n6627 G.n6626 0.624
R8375 G.n3315 G.n3311 0.624
R8376 G.n3317 G.n3310 0.624
R8377 G.n3319 G.n3309 0.624
R8378 G.n3321 G.n3308 0.624
R8379 G.n3323 G.n3307 0.624
R8380 G.n3325 G.n3306 0.624
R8381 G.n3327 G.n3305 0.624
R8382 G.n3329 G.n3304 0.624
R8383 G.n3331 G.n3303 0.624
R8384 G.n3301 G.n3271 0.624
R8385 G.n3299 G.n3272 0.624
R8386 G.n3297 G.n3273 0.624
R8387 G.n3295 G.n3274 0.624
R8388 G.n3293 G.n3275 0.624
R8389 G.n3291 G.n3276 0.624
R8390 G.n3289 G.n3277 0.624
R8391 G.n3287 G.n3278 0.624
R8392 G.n3285 G.n3279 0.624
R8393 G.n3283 G.n3280 0.624
R8394 G.n6591 G.n6590 0.624
R8395 G.n6554 G.n6553 0.624
R8396 G.n6513 G.n6512 0.624
R8397 G.n6469 G.n6468 0.624
R8398 G.n6421 G.n6420 0.624
R8399 G.n6370 G.n6369 0.624
R8400 G.n6317 G.n6316 0.624
R8401 G.n6263 G.n6262 0.624
R8402 G.n6209 G.n6208 0.624
R8403 G.n6155 G.n6154 0.624
R8404 G.n6101 G.n6100 0.624
R8405 G.n6049 G.n6048 0.624
R8406 G.n5998 G.n5997 0.624
R8407 G.n5949 G.n5948 0.624
R8408 G.n5903 G.n5902 0.624
R8409 G.n5858 G.n5857 0.624
R8410 G.n5815 G.n5814 0.624
R8411 G.n5775 G.n5774 0.624
R8412 G.n5736 G.n5735 0.624
R8413 G.n5122 G.n5118 0.624
R8414 G.n5124 G.n5117 0.624
R8415 G.n5126 G.n5116 0.624
R8416 G.n5128 G.n5115 0.624
R8417 G.n5130 G.n5114 0.624
R8418 G.n5132 G.n5113 0.624
R8419 G.n5134 G.n5112 0.624
R8420 G.n5136 G.n5111 0.624
R8421 G.n5138 G.n5110 0.624
R8422 G.n5140 G.n5109 0.624
R8423 G.n5142 G.n5108 0.624
R8424 G.n5144 G.n5107 0.624
R8425 G.n5146 G.n5106 0.624
R8426 G.n5148 G.n5105 0.624
R8427 G.n5150 G.n5104 0.624
R8428 G.n5152 G.n5103 0.624
R8429 G.n5101 G.n5049 0.624
R8430 G.n5099 G.n5050 0.624
R8431 G.n5097 G.n5051 0.624
R8432 G.n5095 G.n5052 0.624
R8433 G.n5093 G.n5053 0.624
R8434 G.n5091 G.n5054 0.624
R8435 G.n5089 G.n5055 0.624
R8436 G.n5087 G.n5056 0.624
R8437 G.n5085 G.n5057 0.624
R8438 G.n5083 G.n5058 0.624
R8439 G.n5081 G.n5059 0.624
R8440 G.n5079 G.n5060 0.624
R8441 G.n5077 G.n5061 0.624
R8442 G.n5075 G.n5062 0.624
R8443 G.n5073 G.n5063 0.624
R8444 G.n5071 G.n5064 0.624
R8445 G.n5069 G.n5065 0.624
R8446 G.n5773 G.n5772 0.624
R8447 G.n5813 G.n5812 0.624
R8448 G.n5856 G.n5855 0.624
R8449 G.n5901 G.n5900 0.624
R8450 G.n5947 G.n5946 0.624
R8451 G.n5996 G.n5995 0.624
R8452 G.n6047 G.n6046 0.624
R8453 G.n6099 G.n6098 0.624
R8454 G.n6153 G.n6152 0.624
R8455 G.n6207 G.n6206 0.624
R8456 G.n6261 G.n6260 0.624
R8457 G.n6315 G.n6314 0.624
R8458 G.n6368 G.n6367 0.624
R8459 G.n6419 G.n6418 0.624
R8460 G.n6467 G.n6466 0.624
R8461 G.n6511 G.n6510 0.624
R8462 G.n6552 G.n6551 0.624
R8463 G.n3249 G.n3246 0.624
R8464 G.n3251 G.n3245 0.624
R8465 G.n3253 G.n3244 0.624
R8466 G.n3255 G.n3243 0.624
R8467 G.n3257 G.n3242 0.624
R8468 G.n3259 G.n3241 0.624
R8469 G.n3261 G.n3240 0.624
R8470 G.n3263 G.n3239 0.624
R8471 G.n3265 G.n3238 0.624
R8472 G.n3267 G.n3237 0.624
R8473 G.n3269 G.n3236 0.624
R8474 G.n3234 G.n3199 0.624
R8475 G.n3232 G.n3200 0.624
R8476 G.n3230 G.n3201 0.624
R8477 G.n3228 G.n3202 0.624
R8478 G.n3226 G.n3203 0.624
R8479 G.n3224 G.n3204 0.624
R8480 G.n3222 G.n3205 0.624
R8481 G.n3220 G.n3206 0.624
R8482 G.n3218 G.n3207 0.624
R8483 G.n3216 G.n3208 0.624
R8484 G.n3214 G.n3209 0.624
R8485 G.n3212 G.n3210 0.624
R8486 G.n6549 G.n6548 0.624
R8487 G.n6508 G.n6507 0.624
R8488 G.n6464 G.n6463 0.624
R8489 G.n6416 G.n6415 0.624
R8490 G.n6365 G.n6364 0.624
R8491 G.n6312 G.n6311 0.624
R8492 G.n6258 G.n6257 0.624
R8493 G.n6204 G.n6203 0.624
R8494 G.n6150 G.n6149 0.624
R8495 G.n6096 G.n6095 0.624
R8496 G.n6044 G.n6043 0.624
R8497 G.n5993 G.n5992 0.624
R8498 G.n5944 G.n5943 0.624
R8499 G.n5898 G.n5897 0.624
R8500 G.n5853 G.n5852 0.624
R8501 G.n5011 G.n5007 0.624
R8502 G.n5013 G.n5006 0.624
R8503 G.n5015 G.n5005 0.624
R8504 G.n5017 G.n5004 0.624
R8505 G.n5019 G.n5003 0.624
R8506 G.n5021 G.n5002 0.624
R8507 G.n5023 G.n5001 0.624
R8508 G.n5025 G.n5000 0.624
R8509 G.n5027 G.n4999 0.624
R8510 G.n5029 G.n4998 0.624
R8511 G.n5031 G.n4997 0.624
R8512 G.n5033 G.n4996 0.624
R8513 G.n5035 G.n4995 0.624
R8514 G.n5037 G.n4994 0.624
R8515 G.n5039 G.n4993 0.624
R8516 G.n5041 G.n4992 0.624
R8517 G.n5043 G.n4991 0.624
R8518 G.n5045 G.n4990 0.624
R8519 G.n5047 G.n4989 0.624
R8520 G.n4987 G.n4926 0.624
R8521 G.n4985 G.n4927 0.624
R8522 G.n4983 G.n4928 0.624
R8523 G.n4981 G.n4929 0.624
R8524 G.n4979 G.n4930 0.624
R8525 G.n4977 G.n4931 0.624
R8526 G.n4975 G.n4932 0.624
R8527 G.n4973 G.n4933 0.624
R8528 G.n4971 G.n4934 0.624
R8529 G.n4969 G.n4935 0.624
R8530 G.n4967 G.n4936 0.624
R8531 G.n4965 G.n4937 0.624
R8532 G.n4963 G.n4938 0.624
R8533 G.n4961 G.n4939 0.624
R8534 G.n4959 G.n4940 0.624
R8535 G.n4957 G.n4941 0.624
R8536 G.n4955 G.n4942 0.624
R8537 G.n4953 G.n4943 0.624
R8538 G.n4951 G.n4944 0.624
R8539 G.n4949 G.n4945 0.624
R8540 G.n5896 G.n5895 0.624
R8541 G.n5942 G.n5941 0.624
R8542 G.n5991 G.n5990 0.624
R8543 G.n6042 G.n6041 0.624
R8544 G.n6094 G.n6093 0.624
R8545 G.n6148 G.n6147 0.624
R8546 G.n6202 G.n6201 0.624
R8547 G.n6256 G.n6255 0.624
R8548 G.n6310 G.n6309 0.624
R8549 G.n6363 G.n6362 0.624
R8550 G.n6414 G.n6413 0.624
R8551 G.n6462 G.n6461 0.624
R8552 G.n6506 G.n6505 0.624
R8553 G.n3173 G.n3171 0.624
R8554 G.n3175 G.n3170 0.624
R8555 G.n3177 G.n3169 0.624
R8556 G.n3179 G.n3168 0.624
R8557 G.n3181 G.n3167 0.624
R8558 G.n3183 G.n3166 0.624
R8559 G.n3185 G.n3165 0.624
R8560 G.n3187 G.n3164 0.624
R8561 G.n3189 G.n3163 0.624
R8562 G.n3191 G.n3162 0.624
R8563 G.n3193 G.n3161 0.624
R8564 G.n3195 G.n3160 0.624
R8565 G.n3197 G.n3159 0.624
R8566 G.n3157 G.n3116 0.624
R8567 G.n3155 G.n3117 0.624
R8568 G.n3153 G.n3118 0.624
R8569 G.n3151 G.n3119 0.624
R8570 G.n3149 G.n3120 0.624
R8571 G.n3147 G.n3121 0.624
R8572 G.n3145 G.n3122 0.624
R8573 G.n3143 G.n3123 0.624
R8574 G.n3141 G.n3124 0.624
R8575 G.n3139 G.n3125 0.624
R8576 G.n3137 G.n3126 0.624
R8577 G.n3135 G.n3127 0.624
R8578 G.n3133 G.n3128 0.624
R8579 G.n3131 G.n3129 0.624
R8580 G.n6459 G.n6458 0.624
R8581 G.n6411 G.n6410 0.624
R8582 G.n6360 G.n6359 0.624
R8583 G.n6307 G.n6306 0.624
R8584 G.n6253 G.n6252 0.624
R8585 G.n6199 G.n6198 0.624
R8586 G.n6145 G.n6144 0.624
R8587 G.n6091 G.n6090 0.624
R8588 G.n6039 G.n6038 0.624
R8589 G.n5988 G.n5987 0.624
R8590 G.n4882 G.n4878 0.624
R8591 G.n4884 G.n4877 0.624
R8592 G.n4886 G.n4876 0.624
R8593 G.n4888 G.n4875 0.624
R8594 G.n4890 G.n4874 0.624
R8595 G.n4892 G.n4873 0.624
R8596 G.n4894 G.n4872 0.624
R8597 G.n4896 G.n4871 0.624
R8598 G.n4898 G.n4870 0.624
R8599 G.n4900 G.n4869 0.624
R8600 G.n4902 G.n4868 0.624
R8601 G.n4904 G.n4867 0.624
R8602 G.n4906 G.n4866 0.624
R8603 G.n4908 G.n4865 0.624
R8604 G.n4910 G.n4864 0.624
R8605 G.n4912 G.n4863 0.624
R8606 G.n4914 G.n4862 0.624
R8607 G.n4916 G.n4861 0.624
R8608 G.n4918 G.n4860 0.624
R8609 G.n4920 G.n4859 0.624
R8610 G.n4922 G.n4858 0.624
R8611 G.n4924 G.n4857 0.624
R8612 G.n4855 G.n4785 0.624
R8613 G.n4853 G.n4786 0.624
R8614 G.n4851 G.n4787 0.624
R8615 G.n4849 G.n4788 0.624
R8616 G.n4847 G.n4789 0.624
R8617 G.n4845 G.n4790 0.624
R8618 G.n4843 G.n4791 0.624
R8619 G.n4841 G.n4792 0.624
R8620 G.n4839 G.n4793 0.624
R8621 G.n4837 G.n4794 0.624
R8622 G.n4835 G.n4795 0.624
R8623 G.n4833 G.n4796 0.624
R8624 G.n4831 G.n4797 0.624
R8625 G.n4829 G.n4798 0.624
R8626 G.n4827 G.n4799 0.624
R8627 G.n4825 G.n4800 0.624
R8628 G.n4823 G.n4801 0.624
R8629 G.n4821 G.n4802 0.624
R8630 G.n4819 G.n4803 0.624
R8631 G.n4817 G.n4804 0.624
R8632 G.n4815 G.n4805 0.624
R8633 G.n4813 G.n4806 0.624
R8634 G.n4811 G.n4807 0.624
R8635 G.n6037 G.n6036 0.624
R8636 G.n6089 G.n6088 0.624
R8637 G.n6143 G.n6142 0.624
R8638 G.n6197 G.n6196 0.624
R8639 G.n6251 G.n6250 0.624
R8640 G.n6305 G.n6304 0.624
R8641 G.n6358 G.n6357 0.624
R8642 G.n6409 G.n6408 0.624
R8643 G.n3088 G.n3084 0.624
R8644 G.n3090 G.n3083 0.624
R8645 G.n3092 G.n3082 0.624
R8646 G.n3094 G.n3081 0.624
R8647 G.n3096 G.n3080 0.624
R8648 G.n3098 G.n3079 0.624
R8649 G.n3100 G.n3078 0.624
R8650 G.n3102 G.n3077 0.624
R8651 G.n3104 G.n3076 0.624
R8652 G.n3106 G.n3075 0.624
R8653 G.n3108 G.n3074 0.624
R8654 G.n3110 G.n3073 0.624
R8655 G.n3112 G.n3072 0.624
R8656 G.n3114 G.n3071 0.624
R8657 G.n3069 G.n3023 0.624
R8658 G.n3067 G.n3024 0.624
R8659 G.n3065 G.n3025 0.624
R8660 G.n3063 G.n3026 0.624
R8661 G.n3061 G.n3027 0.624
R8662 G.n3059 G.n3028 0.624
R8663 G.n3057 G.n3029 0.624
R8664 G.n3055 G.n3030 0.624
R8665 G.n3053 G.n3031 0.624
R8666 G.n3051 G.n3032 0.624
R8667 G.n3049 G.n3033 0.624
R8668 G.n3047 G.n3034 0.624
R8669 G.n3045 G.n3035 0.624
R8670 G.n3043 G.n3036 0.624
R8671 G.n3041 G.n3037 0.624
R8672 G.n6355 G.n6354 0.624
R8673 G.n6302 G.n6301 0.624
R8674 G.n6248 G.n6247 0.624
R8675 G.n6194 G.n6193 0.624
R8676 G.n6140 G.n6139 0.624
R8677 G.n4735 G.n4731 0.624
R8678 G.n4737 G.n4730 0.624
R8679 G.n4739 G.n4729 0.624
R8680 G.n4741 G.n4728 0.624
R8681 G.n4743 G.n4727 0.624
R8682 G.n4745 G.n4726 0.624
R8683 G.n4747 G.n4725 0.624
R8684 G.n4749 G.n4724 0.624
R8685 G.n4751 G.n4723 0.624
R8686 G.n4753 G.n4722 0.624
R8687 G.n4755 G.n4721 0.624
R8688 G.n4757 G.n4720 0.624
R8689 G.n4759 G.n4719 0.624
R8690 G.n4761 G.n4718 0.624
R8691 G.n4763 G.n4717 0.624
R8692 G.n4765 G.n4716 0.624
R8693 G.n4767 G.n4715 0.624
R8694 G.n4769 G.n4714 0.624
R8695 G.n4771 G.n4713 0.624
R8696 G.n4773 G.n4712 0.624
R8697 G.n4775 G.n4711 0.624
R8698 G.n4777 G.n4710 0.624
R8699 G.n4779 G.n4709 0.624
R8700 G.n4781 G.n4708 0.624
R8701 G.n4783 G.n4707 0.624
R8702 G.n4705 G.n4631 0.624
R8703 G.n4703 G.n4632 0.624
R8704 G.n4701 G.n4633 0.624
R8705 G.n4699 G.n4634 0.624
R8706 G.n4697 G.n4635 0.624
R8707 G.n4695 G.n4636 0.624
R8708 G.n4693 G.n4637 0.624
R8709 G.n4691 G.n4638 0.624
R8710 G.n4689 G.n4639 0.624
R8711 G.n4687 G.n4640 0.624
R8712 G.n4685 G.n4641 0.624
R8713 G.n4683 G.n4642 0.624
R8714 G.n4681 G.n4643 0.624
R8715 G.n4679 G.n4644 0.624
R8716 G.n4677 G.n4645 0.624
R8717 G.n4675 G.n4646 0.624
R8718 G.n4673 G.n4647 0.624
R8719 G.n4671 G.n4648 0.624
R8720 G.n4669 G.n4649 0.624
R8721 G.n4667 G.n4650 0.624
R8722 G.n4665 G.n4651 0.624
R8723 G.n4663 G.n4652 0.624
R8724 G.n4661 G.n4653 0.624
R8725 G.n4659 G.n4654 0.624
R8726 G.n4657 G.n4655 0.624
R8727 G.n1089 G.n1087 0.624
R8728 G.n1177 G.n1175 0.624
R8729 G.n1265 G.n1263 0.624
R8730 G.n1353 G.n1351 0.624
R8731 G.n1441 G.n1439 0.624
R8732 G.n1528 G.n1527 0.624
R8733 G.n2991 G.n2989 0.624
R8734 G.n2993 G.n2988 0.624
R8735 G.n2995 G.n2987 0.624
R8736 G.n2997 G.n2986 0.624
R8737 G.n2999 G.n2985 0.624
R8738 G.n3001 G.n2984 0.624
R8739 G.n3003 G.n2983 0.624
R8740 G.n3005 G.n2982 0.624
R8741 G.n3007 G.n2981 0.624
R8742 G.n3009 G.n2980 0.624
R8743 G.n3011 G.n2979 0.624
R8744 G.n3013 G.n2978 0.624
R8745 G.n3015 G.n2977 0.624
R8746 G.n3017 G.n2976 0.624
R8747 G.n3019 G.n2975 0.624
R8748 G.n3021 G.n2974 0.624
R8749 G.n2972 G.n2928 0.624
R8750 G.n2970 G.n2929 0.624
R8751 G.n2968 G.n2930 0.624
R8752 G.n2966 G.n2931 0.624
R8753 G.n2964 G.n2932 0.624
R8754 G.n2962 G.n2933 0.624
R8755 G.n2960 G.n2934 0.624
R8756 G.n2958 G.n2935 0.624
R8757 G.n2956 G.n2936 0.624
R8758 G.n2954 G.n2937 0.624
R8759 G.n2952 G.n2938 0.624
R8760 G.n2950 G.n2939 0.624
R8761 G.n2948 G.n2940 0.624
R8762 G.n2946 G.n2941 0.624
R8763 G.n2944 G.n2942 0.624
R8764 G.n1615 G.n1614 0.624
R8765 G.n1531 G.n1529 0.624
R8766 G.n1444 G.n1442 0.624
R8767 G.n1356 G.n1354 0.624
R8768 G.n1268 G.n1266 0.624
R8769 G.n1180 G.n1178 0.624
R8770 G.n1092 G.n1090 0.624
R8771 G.n1004 G.n1002 0.624
R8772 G.n4583 G.n4581 0.624
R8773 G.n4585 G.n4580 0.624
R8774 G.n4587 G.n4579 0.624
R8775 G.n4589 G.n4578 0.624
R8776 G.n4591 G.n4577 0.624
R8777 G.n4593 G.n4576 0.624
R8778 G.n4595 G.n4575 0.624
R8779 G.n4597 G.n4574 0.624
R8780 G.n4599 G.n4573 0.624
R8781 G.n4601 G.n4572 0.624
R8782 G.n4603 G.n4571 0.624
R8783 G.n4605 G.n4570 0.624
R8784 G.n4607 G.n4569 0.624
R8785 G.n4609 G.n4568 0.624
R8786 G.n4611 G.n4567 0.624
R8787 G.n4613 G.n4566 0.624
R8788 G.n4615 G.n4565 0.624
R8789 G.n4617 G.n4564 0.624
R8790 G.n4619 G.n4563 0.624
R8791 G.n4621 G.n4562 0.624
R8792 G.n4623 G.n4561 0.624
R8793 G.n4625 G.n4560 0.624
R8794 G.n4627 G.n4559 0.624
R8795 G.n4629 G.n4558 0.624
R8796 G.n4556 G.n4488 0.624
R8797 G.n4554 G.n4489 0.624
R8798 G.n4552 G.n4490 0.624
R8799 G.n4550 G.n4491 0.624
R8800 G.n4548 G.n4492 0.624
R8801 G.n4546 G.n4493 0.624
R8802 G.n4544 G.n4494 0.624
R8803 G.n4542 G.n4495 0.624
R8804 G.n4540 G.n4496 0.624
R8805 G.n4538 G.n4497 0.624
R8806 G.n4536 G.n4498 0.624
R8807 G.n4534 G.n4499 0.624
R8808 G.n4532 G.n4500 0.624
R8809 G.n4530 G.n4501 0.624
R8810 G.n4528 G.n4502 0.624
R8811 G.n4526 G.n4503 0.624
R8812 G.n4524 G.n4504 0.624
R8813 G.n4522 G.n4505 0.624
R8814 G.n4520 G.n4506 0.624
R8815 G.n4518 G.n4507 0.624
R8816 G.n4516 G.n4508 0.624
R8817 G.n4514 G.n4509 0.624
R8818 G.n4512 G.n4510 0.624
R8819 G.n922 G.n920 0.624
R8820 G.n1007 G.n1005 0.624
R8821 G.n1095 G.n1093 0.624
R8822 G.n1183 G.n1181 0.624
R8823 G.n1271 G.n1269 0.624
R8824 G.n1359 G.n1357 0.624
R8825 G.n1447 G.n1445 0.624
R8826 G.n1534 G.n1532 0.624
R8827 G.n1617 G.n1616 0.624
R8828 G.n2898 G.n2896 0.624
R8829 G.n2900 G.n2895 0.624
R8830 G.n2902 G.n2894 0.624
R8831 G.n2904 G.n2893 0.624
R8832 G.n2906 G.n2892 0.624
R8833 G.n2908 G.n2891 0.624
R8834 G.n2910 G.n2890 0.624
R8835 G.n2912 G.n2889 0.624
R8836 G.n2914 G.n2888 0.624
R8837 G.n2916 G.n2887 0.624
R8838 G.n2918 G.n2886 0.624
R8839 G.n2920 G.n2885 0.624
R8840 G.n2922 G.n2884 0.624
R8841 G.n2924 G.n2883 0.624
R8842 G.n2926 G.n2882 0.624
R8843 G.n2880 G.n2839 0.624
R8844 G.n2878 G.n2840 0.624
R8845 G.n2876 G.n2841 0.624
R8846 G.n2874 G.n2842 0.624
R8847 G.n2872 G.n2843 0.624
R8848 G.n2870 G.n2844 0.624
R8849 G.n2868 G.n2845 0.624
R8850 G.n2866 G.n2846 0.624
R8851 G.n2864 G.n2847 0.624
R8852 G.n2862 G.n2848 0.624
R8853 G.n2860 G.n2849 0.624
R8854 G.n2858 G.n2850 0.624
R8855 G.n2856 G.n2851 0.624
R8856 G.n2854 G.n2852 0.624
R8857 G.n1698 G.n1697 0.624
R8858 G.n1620 G.n1618 0.624
R8859 G.n1537 G.n1535 0.624
R8860 G.n1450 G.n1448 0.624
R8861 G.n1362 G.n1360 0.624
R8862 G.n1274 G.n1272 0.624
R8863 G.n1186 G.n1184 0.624
R8864 G.n1098 G.n1096 0.624
R8865 G.n1010 G.n1008 0.624
R8866 G.n925 G.n923 0.624
R8867 G.n4442 G.n4440 0.624
R8868 G.n4444 G.n4439 0.624
R8869 G.n4446 G.n4438 0.624
R8870 G.n4448 G.n4437 0.624
R8871 G.n4450 G.n4436 0.624
R8872 G.n4452 G.n4435 0.624
R8873 G.n4454 G.n4434 0.624
R8874 G.n4456 G.n4433 0.624
R8875 G.n4458 G.n4432 0.624
R8876 G.n4460 G.n4431 0.624
R8877 G.n4462 G.n4430 0.624
R8878 G.n4464 G.n4429 0.624
R8879 G.n4466 G.n4428 0.624
R8880 G.n4468 G.n4427 0.624
R8881 G.n4470 G.n4426 0.624
R8882 G.n4472 G.n4425 0.624
R8883 G.n4474 G.n4424 0.624
R8884 G.n4476 G.n4423 0.624
R8885 G.n4478 G.n4422 0.624
R8886 G.n4480 G.n4421 0.624
R8887 G.n4482 G.n4420 0.624
R8888 G.n4484 G.n4419 0.624
R8889 G.n4486 G.n4418 0.624
R8890 G.n4416 G.n4351 0.624
R8891 G.n4414 G.n4352 0.624
R8892 G.n4412 G.n4353 0.624
R8893 G.n4410 G.n4354 0.624
R8894 G.n4408 G.n4355 0.624
R8895 G.n4406 G.n4356 0.624
R8896 G.n4404 G.n4357 0.624
R8897 G.n4402 G.n4358 0.624
R8898 G.n4400 G.n4359 0.624
R8899 G.n4398 G.n4360 0.624
R8900 G.n4396 G.n4361 0.624
R8901 G.n4394 G.n4362 0.624
R8902 G.n4392 G.n4363 0.624
R8903 G.n4390 G.n4364 0.624
R8904 G.n4388 G.n4365 0.624
R8905 G.n4386 G.n4366 0.624
R8906 G.n4384 G.n4367 0.624
R8907 G.n4382 G.n4368 0.624
R8908 G.n4380 G.n4369 0.624
R8909 G.n4378 G.n4370 0.624
R8910 G.n4376 G.n4371 0.624
R8911 G.n4374 G.n4372 0.624
R8912 G.n846 G.n844 0.624
R8913 G.n928 G.n926 0.624
R8914 G.n1013 G.n1011 0.624
R8915 G.n1101 G.n1099 0.624
R8916 G.n1189 G.n1187 0.624
R8917 G.n1277 G.n1275 0.624
R8918 G.n1365 G.n1363 0.624
R8919 G.n1453 G.n1451 0.624
R8920 G.n1540 G.n1538 0.624
R8921 G.n1623 G.n1621 0.624
R8922 G.n1701 G.n1699 0.624
R8923 G.n2811 G.n2810 0.624
R8924 G.n2813 G.n2809 0.624
R8925 G.n2815 G.n2808 0.624
R8926 G.n2817 G.n2807 0.624
R8927 G.n2819 G.n2806 0.624
R8928 G.n2821 G.n2805 0.624
R8929 G.n2823 G.n2804 0.624
R8930 G.n2825 G.n2803 0.624
R8931 G.n2827 G.n2802 0.624
R8932 G.n2829 G.n2801 0.624
R8933 G.n2831 G.n2800 0.624
R8934 G.n2833 G.n2799 0.624
R8935 G.n2835 G.n2798 0.624
R8936 G.n2837 G.n2797 0.624
R8937 G.n2795 G.n2757 0.624
R8938 G.n2793 G.n2758 0.624
R8939 G.n2791 G.n2759 0.624
R8940 G.n2789 G.n2760 0.624
R8941 G.n2787 G.n2761 0.624
R8942 G.n2785 G.n2762 0.624
R8943 G.n2783 G.n2763 0.624
R8944 G.n2781 G.n2764 0.624
R8945 G.n2779 G.n2765 0.624
R8946 G.n2777 G.n2766 0.624
R8947 G.n2775 G.n2767 0.624
R8948 G.n2773 G.n2768 0.624
R8949 G.n2771 G.n2769 0.624
R8950 G.n1776 G.n1775 0.624
R8951 G.n1704 G.n1702 0.624
R8952 G.n1626 G.n1624 0.624
R8953 G.n1543 G.n1541 0.624
R8954 G.n1456 G.n1454 0.624
R8955 G.n1368 G.n1366 0.624
R8956 G.n1280 G.n1278 0.624
R8957 G.n1192 G.n1190 0.624
R8958 G.n1104 G.n1102 0.624
R8959 G.n1016 G.n1014 0.624
R8960 G.n931 G.n929 0.624
R8961 G.n849 G.n847 0.624
R8962 G.n773 G.n771 0.624
R8963 G.n4309 G.n4307 0.624
R8964 G.n4311 G.n4306 0.624
R8965 G.n4313 G.n4305 0.624
R8966 G.n4315 G.n4304 0.624
R8967 G.n4317 G.n4303 0.624
R8968 G.n4319 G.n4302 0.624
R8969 G.n4321 G.n4301 0.624
R8970 G.n4323 G.n4300 0.624
R8971 G.n4325 G.n4299 0.624
R8972 G.n4327 G.n4298 0.624
R8973 G.n4329 G.n4297 0.624
R8974 G.n4331 G.n4296 0.624
R8975 G.n4333 G.n4295 0.624
R8976 G.n4335 G.n4294 0.624
R8977 G.n4337 G.n4293 0.624
R8978 G.n4339 G.n4292 0.624
R8979 G.n4341 G.n4291 0.624
R8980 G.n4343 G.n4290 0.624
R8981 G.n4345 G.n4289 0.624
R8982 G.n4347 G.n4288 0.624
R8983 G.n4349 G.n4287 0.624
R8984 G.n4285 G.n4226 0.624
R8985 G.n4283 G.n4227 0.624
R8986 G.n4281 G.n4228 0.624
R8987 G.n4279 G.n4229 0.624
R8988 G.n4277 G.n4230 0.624
R8989 G.n4275 G.n4231 0.624
R8990 G.n4273 G.n4232 0.624
R8991 G.n4271 G.n4233 0.624
R8992 G.n4269 G.n4234 0.624
R8993 G.n4267 G.n4235 0.624
R8994 G.n4265 G.n4236 0.624
R8995 G.n4263 G.n4237 0.624
R8996 G.n4261 G.n4238 0.624
R8997 G.n4259 G.n4239 0.624
R8998 G.n4257 G.n4240 0.624
R8999 G.n4255 G.n4241 0.624
R9000 G.n4253 G.n4242 0.624
R9001 G.n4251 G.n4243 0.624
R9002 G.n4249 G.n4244 0.624
R9003 G.n4247 G.n4245 0.624
R9004 G.n703 G.n701 0.624
R9005 G.n776 G.n774 0.624
R9006 G.n852 G.n850 0.624
R9007 G.n934 G.n932 0.624
R9008 G.n1019 G.n1017 0.624
R9009 G.n1107 G.n1105 0.624
R9010 G.n1195 G.n1193 0.624
R9011 G.n1283 G.n1281 0.624
R9012 G.n1371 G.n1369 0.624
R9013 G.n1459 G.n1457 0.624
R9014 G.n1546 G.n1544 0.624
R9015 G.n1629 G.n1627 0.624
R9016 G.n1707 G.n1705 0.624
R9017 G.n1779 G.n1777 0.624
R9018 G.n1848 G.n1847 0.624
R9019 G.n2733 G.n2731 0.624
R9020 G.n2735 G.n2730 0.624
R9021 G.n2737 G.n2729 0.624
R9022 G.n2739 G.n2728 0.624
R9023 G.n2741 G.n2727 0.624
R9024 G.n2743 G.n2726 0.624
R9025 G.n2745 G.n2725 0.624
R9026 G.n2747 G.n2724 0.624
R9027 G.n2749 G.n2723 0.624
R9028 G.n2751 G.n2722 0.624
R9029 G.n2753 G.n2721 0.624
R9030 G.n2755 G.n2720 0.624
R9031 G.n2718 G.n2683 0.624
R9032 G.n2716 G.n2684 0.624
R9033 G.n2714 G.n2685 0.624
R9034 G.n2712 G.n2686 0.624
R9035 G.n2710 G.n2687 0.624
R9036 G.n2708 G.n2688 0.624
R9037 G.n2706 G.n2689 0.624
R9038 G.n2704 G.n2690 0.624
R9039 G.n2702 G.n2691 0.624
R9040 G.n2700 G.n2692 0.624
R9041 G.n2698 G.n2693 0.624
R9042 G.n2696 G.n2694 0.624
R9043 G.n1850 G.n1849 0.624
R9044 G.n1782 G.n1780 0.624
R9045 G.n1710 G.n1708 0.624
R9046 G.n1632 G.n1630 0.624
R9047 G.n1549 G.n1547 0.624
R9048 G.n1462 G.n1460 0.624
R9049 G.n1374 G.n1372 0.624
R9050 G.n1286 G.n1284 0.624
R9051 G.n1198 G.n1196 0.624
R9052 G.n1110 G.n1108 0.624
R9053 G.n1022 G.n1020 0.624
R9054 G.n937 G.n935 0.624
R9055 G.n855 G.n853 0.624
R9056 G.n779 G.n777 0.624
R9057 G.n706 G.n704 0.624
R9058 G.n636 G.n634 0.624
R9059 G.n4188 G.n4186 0.624
R9060 G.n4190 G.n4185 0.624
R9061 G.n4192 G.n4184 0.624
R9062 G.n4194 G.n4183 0.624
R9063 G.n4196 G.n4182 0.624
R9064 G.n4198 G.n4181 0.624
R9065 G.n4200 G.n4180 0.624
R9066 G.n4202 G.n4179 0.624
R9067 G.n4204 G.n4178 0.624
R9068 G.n4206 G.n4177 0.624
R9069 G.n4208 G.n4176 0.624
R9070 G.n4210 G.n4175 0.624
R9071 G.n4212 G.n4174 0.624
R9072 G.n4214 G.n4173 0.624
R9073 G.n4216 G.n4172 0.624
R9074 G.n4218 G.n4171 0.624
R9075 G.n4220 G.n4170 0.624
R9076 G.n4222 G.n4169 0.624
R9077 G.n4224 G.n4168 0.624
R9078 G.n4166 G.n4113 0.624
R9079 G.n4164 G.n4114 0.624
R9080 G.n4162 G.n4115 0.624
R9081 G.n4160 G.n4116 0.624
R9082 G.n4158 G.n4117 0.624
R9083 G.n4156 G.n4118 0.624
R9084 G.n4154 G.n4119 0.624
R9085 G.n4152 G.n4120 0.624
R9086 G.n4150 G.n4121 0.624
R9087 G.n4148 G.n4122 0.624
R9088 G.n4146 G.n4123 0.624
R9089 G.n4144 G.n4124 0.624
R9090 G.n4142 G.n4125 0.624
R9091 G.n4140 G.n4126 0.624
R9092 G.n4138 G.n4127 0.624
R9093 G.n4136 G.n4128 0.624
R9094 G.n4134 G.n4129 0.624
R9095 G.n4132 G.n4130 0.624
R9096 G.n572 G.n570 0.624
R9097 G.n639 G.n637 0.624
R9098 G.n709 G.n707 0.624
R9099 G.n782 G.n780 0.624
R9100 G.n858 G.n856 0.624
R9101 G.n940 G.n938 0.624
R9102 G.n1025 G.n1023 0.624
R9103 G.n1113 G.n1111 0.624
R9104 G.n1201 G.n1199 0.624
R9105 G.n1289 G.n1287 0.624
R9106 G.n1377 G.n1375 0.624
R9107 G.n1465 G.n1463 0.624
R9108 G.n1552 G.n1550 0.624
R9109 G.n1635 G.n1633 0.624
R9110 G.n1713 G.n1711 0.624
R9111 G.n1785 G.n1783 0.624
R9112 G.n1853 G.n1851 0.624
R9113 G.n1916 G.n1915 0.624
R9114 G.n2661 G.n2659 0.624
R9115 G.n2663 G.n2658 0.624
R9116 G.n2665 G.n2657 0.624
R9117 G.n2667 G.n2656 0.624
R9118 G.n2669 G.n2655 0.624
R9119 G.n2671 G.n2654 0.624
R9120 G.n2673 G.n2653 0.624
R9121 G.n2675 G.n2652 0.624
R9122 G.n2677 G.n2651 0.624
R9123 G.n2679 G.n2650 0.624
R9124 G.n2681 G.n2649 0.624
R9125 G.n2647 G.n2615 0.624
R9126 G.n2645 G.n2616 0.624
R9127 G.n2643 G.n2617 0.624
R9128 G.n2641 G.n2618 0.624
R9129 G.n2639 G.n2619 0.624
R9130 G.n2637 G.n2620 0.624
R9131 G.n2635 G.n2621 0.624
R9132 G.n2633 G.n2622 0.624
R9133 G.n2631 G.n2623 0.624
R9134 G.n2629 G.n2624 0.624
R9135 G.n2627 G.n2625 0.624
R9136 G.n1918 G.n1917 0.624
R9137 G.n1856 G.n1854 0.624
R9138 G.n1788 G.n1786 0.624
R9139 G.n1716 G.n1714 0.624
R9140 G.n1638 G.n1636 0.624
R9141 G.n1555 G.n1553 0.624
R9142 G.n1468 G.n1466 0.624
R9143 G.n1380 G.n1378 0.624
R9144 G.n1292 G.n1290 0.624
R9145 G.n1204 G.n1202 0.624
R9146 G.n1116 G.n1114 0.624
R9147 G.n1028 G.n1026 0.624
R9148 G.n943 G.n941 0.624
R9149 G.n861 G.n859 0.624
R9150 G.n785 G.n783 0.624
R9151 G.n712 G.n710 0.624
R9152 G.n642 G.n640 0.624
R9153 G.n575 G.n573 0.624
R9154 G.n511 G.n509 0.624
R9155 G.n4079 G.n4077 0.624
R9156 G.n4081 G.n4076 0.624
R9157 G.n4083 G.n4075 0.624
R9158 G.n4085 G.n4074 0.624
R9159 G.n4087 G.n4073 0.624
R9160 G.n4089 G.n4072 0.624
R9161 G.n4091 G.n4071 0.624
R9162 G.n4093 G.n4070 0.624
R9163 G.n4095 G.n4069 0.624
R9164 G.n4097 G.n4068 0.624
R9165 G.n4099 G.n4067 0.624
R9166 G.n4101 G.n4066 0.624
R9167 G.n4103 G.n4065 0.624
R9168 G.n4105 G.n4064 0.624
R9169 G.n4107 G.n4063 0.624
R9170 G.n4109 G.n4062 0.624
R9171 G.n4111 G.n4061 0.624
R9172 G.n4059 G.n4012 0.624
R9173 G.n4057 G.n4013 0.624
R9174 G.n4055 G.n4014 0.624
R9175 G.n4053 G.n4015 0.624
R9176 G.n4051 G.n4016 0.624
R9177 G.n4049 G.n4017 0.624
R9178 G.n4047 G.n4018 0.624
R9179 G.n4045 G.n4019 0.624
R9180 G.n4043 G.n4020 0.624
R9181 G.n4041 G.n4021 0.624
R9182 G.n4039 G.n4022 0.624
R9183 G.n4037 G.n4023 0.624
R9184 G.n4035 G.n4024 0.624
R9185 G.n4033 G.n4025 0.624
R9186 G.n4031 G.n4026 0.624
R9187 G.n4029 G.n4027 0.624
R9188 G.n453 G.n451 0.624
R9189 G.n514 G.n512 0.624
R9190 G.n578 G.n576 0.624
R9191 G.n645 G.n643 0.624
R9192 G.n715 G.n713 0.624
R9193 G.n788 G.n786 0.624
R9194 G.n864 G.n862 0.624
R9195 G.n946 G.n944 0.624
R9196 G.n1031 G.n1029 0.624
R9197 G.n1119 G.n1117 0.624
R9198 G.n1207 G.n1205 0.624
R9199 G.n1295 G.n1293 0.624
R9200 G.n1383 G.n1381 0.624
R9201 G.n1471 G.n1469 0.624
R9202 G.n1558 G.n1556 0.624
R9203 G.n1641 G.n1639 0.624
R9204 G.n1719 G.n1717 0.624
R9205 G.n1791 G.n1789 0.624
R9206 G.n1859 G.n1857 0.624
R9207 G.n1921 G.n1919 0.624
R9208 G.n1978 G.n1977 0.624
R9209 G.n2595 G.n2593 0.624
R9210 G.n2597 G.n2592 0.624
R9211 G.n2599 G.n2591 0.624
R9212 G.n2601 G.n2590 0.624
R9213 G.n2603 G.n2589 0.624
R9214 G.n2605 G.n2588 0.624
R9215 G.n2607 G.n2587 0.624
R9216 G.n2609 G.n2586 0.624
R9217 G.n2611 G.n2585 0.624
R9218 G.n2613 G.n2584 0.624
R9219 G.n2582 G.n2554 0.624
R9220 G.n2580 G.n2555 0.624
R9221 G.n2578 G.n2556 0.624
R9222 G.n2576 G.n2557 0.624
R9223 G.n2574 G.n2558 0.624
R9224 G.n2572 G.n2559 0.624
R9225 G.n2570 G.n2560 0.624
R9226 G.n2568 G.n2561 0.624
R9227 G.n2566 G.n2562 0.624
R9228 G.n2564 G.n2563 0.624
R9229 G.n1981 G.n1979 0.624
R9230 G.n1924 G.n1922 0.624
R9231 G.n1862 G.n1860 0.624
R9232 G.n1794 G.n1792 0.624
R9233 G.n1722 G.n1720 0.624
R9234 G.n1644 G.n1642 0.624
R9235 G.n1561 G.n1559 0.624
R9236 G.n1474 G.n1472 0.624
R9237 G.n1386 G.n1384 0.624
R9238 G.n1298 G.n1296 0.624
R9239 G.n1210 G.n1208 0.624
R9240 G.n1122 G.n1120 0.624
R9241 G.n1034 G.n1032 0.624
R9242 G.n949 G.n947 0.624
R9243 G.n867 G.n865 0.624
R9244 G.n791 G.n789 0.624
R9245 G.n718 G.n716 0.624
R9246 G.n648 G.n646 0.624
R9247 G.n581 G.n579 0.624
R9248 G.n517 G.n515 0.624
R9249 G.n456 G.n454 0.624
R9250 G.n398 G.n396 0.624
R9251 G.n3982 G.n3980 0.624
R9252 G.n3984 G.n3979 0.624
R9253 G.n3986 G.n3978 0.624
R9254 G.n3988 G.n3977 0.624
R9255 G.n3990 G.n3976 0.624
R9256 G.n3992 G.n3975 0.624
R9257 G.n3994 G.n3974 0.624
R9258 G.n3996 G.n3973 0.624
R9259 G.n3998 G.n3972 0.624
R9260 G.n4000 G.n3971 0.624
R9261 G.n4002 G.n3970 0.624
R9262 G.n4004 G.n3969 0.624
R9263 G.n4006 G.n3968 0.624
R9264 G.n4008 G.n3967 0.624
R9265 G.n4010 G.n3966 0.624
R9266 G.n3964 G.n3920 0.624
R9267 G.n3962 G.n3921 0.624
R9268 G.n3960 G.n3922 0.624
R9269 G.n3958 G.n3923 0.624
R9270 G.n3956 G.n3924 0.624
R9271 G.n3954 G.n3925 0.624
R9272 G.n3952 G.n3926 0.624
R9273 G.n3950 G.n3927 0.624
R9274 G.n3948 G.n3928 0.624
R9275 G.n3946 G.n3929 0.624
R9276 G.n3944 G.n3930 0.624
R9277 G.n3942 G.n3931 0.624
R9278 G.n3940 G.n3932 0.624
R9279 G.n3938 G.n3933 0.624
R9280 G.n3936 G.n3934 0.624
R9281 G.n401 G.n399 0.624
R9282 G.n459 G.n457 0.624
R9283 G.n520 G.n518 0.624
R9284 G.n584 G.n582 0.624
R9285 G.n651 G.n649 0.624
R9286 G.n721 G.n719 0.624
R9287 G.n794 G.n792 0.624
R9288 G.n870 G.n868 0.624
R9289 G.n952 G.n950 0.624
R9290 G.n1037 G.n1035 0.624
R9291 G.n1125 G.n1123 0.624
R9292 G.n1213 G.n1211 0.624
R9293 G.n1301 G.n1299 0.624
R9294 G.n1389 G.n1387 0.624
R9295 G.n1477 G.n1475 0.624
R9296 G.n1564 G.n1562 0.624
R9297 G.n1647 G.n1645 0.624
R9298 G.n1725 G.n1723 0.624
R9299 G.n1797 G.n1795 0.624
R9300 G.n1865 G.n1863 0.624
R9301 G.n1927 G.n1925 0.624
R9302 G.n1984 G.n1982 0.624
R9303 G.n2035 G.n2034 0.624
R9304 G.n2536 G.n2534 0.624
R9305 G.n2538 G.n2533 0.624
R9306 G.n2540 G.n2532 0.624
R9307 G.n2542 G.n2531 0.624
R9308 G.n2544 G.n2530 0.624
R9309 G.n2546 G.n2529 0.624
R9310 G.n2548 G.n2528 0.624
R9311 G.n2550 G.n2527 0.624
R9312 G.n2552 G.n2526 0.624
R9313 G.n2524 G.n2499 0.624
R9314 G.n2522 G.n2500 0.624
R9315 G.n2520 G.n2501 0.624
R9316 G.n2518 G.n2502 0.624
R9317 G.n2516 G.n2503 0.624
R9318 G.n2514 G.n2504 0.624
R9319 G.n2512 G.n2505 0.624
R9320 G.n2510 G.n2506 0.624
R9321 G.n2508 G.n2507 0.624
R9322 G.n2038 G.n2036 0.624
R9323 G.n1987 G.n1985 0.624
R9324 G.n1930 G.n1928 0.624
R9325 G.n1868 G.n1866 0.624
R9326 G.n1800 G.n1798 0.624
R9327 G.n1728 G.n1726 0.624
R9328 G.n1650 G.n1648 0.624
R9329 G.n1567 G.n1565 0.624
R9330 G.n1480 G.n1478 0.624
R9331 G.n1392 G.n1390 0.624
R9332 G.n1304 G.n1302 0.624
R9333 G.n1216 G.n1214 0.624
R9334 G.n1128 G.n1126 0.624
R9335 G.n1040 G.n1038 0.624
R9336 G.n955 G.n953 0.624
R9337 G.n873 G.n871 0.624
R9338 G.n797 G.n795 0.624
R9339 G.n724 G.n722 0.624
R9340 G.n654 G.n652 0.624
R9341 G.n587 G.n585 0.624
R9342 G.n523 G.n521 0.624
R9343 G.n462 G.n460 0.624
R9344 G.n404 G.n402 0.624
R9345 G.n349 G.n347 0.624
R9346 G.n3892 G.n3890 0.624
R9347 G.n3894 G.n3889 0.624
R9348 G.n3896 G.n3888 0.624
R9349 G.n3898 G.n3887 0.624
R9350 G.n3900 G.n3886 0.624
R9351 G.n3902 G.n3885 0.624
R9352 G.n3904 G.n3884 0.624
R9353 G.n3906 G.n3883 0.624
R9354 G.n3908 G.n3882 0.624
R9355 G.n3910 G.n3881 0.624
R9356 G.n3912 G.n3880 0.624
R9357 G.n3914 G.n3879 0.624
R9358 G.n3916 G.n3878 0.624
R9359 G.n3918 G.n3877 0.624
R9360 G.n3875 G.n3837 0.624
R9361 G.n3873 G.n3838 0.624
R9362 G.n3871 G.n3839 0.624
R9363 G.n3869 G.n3840 0.624
R9364 G.n3867 G.n3841 0.624
R9365 G.n3865 G.n3842 0.624
R9366 G.n3863 G.n3843 0.624
R9367 G.n3861 G.n3844 0.624
R9368 G.n3859 G.n3845 0.624
R9369 G.n3857 G.n3846 0.624
R9370 G.n3855 G.n3847 0.624
R9371 G.n3853 G.n3848 0.624
R9372 G.n3851 G.n3849 0.624
R9373 G.n303 G.n301 0.624
R9374 G.n352 G.n350 0.624
R9375 G.n407 G.n405 0.624
R9376 G.n465 G.n463 0.624
R9377 G.n526 G.n524 0.624
R9378 G.n590 G.n588 0.624
R9379 G.n657 G.n655 0.624
R9380 G.n727 G.n725 0.624
R9381 G.n800 G.n798 0.624
R9382 G.n876 G.n874 0.624
R9383 G.n958 G.n956 0.624
R9384 G.n1043 G.n1041 0.624
R9385 G.n1131 G.n1129 0.624
R9386 G.n1219 G.n1217 0.624
R9387 G.n1307 G.n1305 0.624
R9388 G.n1395 G.n1393 0.624
R9389 G.n1483 G.n1481 0.624
R9390 G.n1570 G.n1568 0.624
R9391 G.n1653 G.n1651 0.624
R9392 G.n1731 G.n1729 0.624
R9393 G.n1803 G.n1801 0.624
R9394 G.n1871 G.n1869 0.624
R9395 G.n1933 G.n1931 0.624
R9396 G.n1990 G.n1988 0.624
R9397 G.n2041 G.n2039 0.624
R9398 G.n2086 G.n2085 0.624
R9399 G.n2483 G.n2481 0.624
R9400 G.n2485 G.n2480 0.624
R9401 G.n2487 G.n2479 0.624
R9402 G.n2489 G.n2478 0.624
R9403 G.n2491 G.n2477 0.624
R9404 G.n2493 G.n2476 0.624
R9405 G.n2495 G.n2475 0.624
R9406 G.n2497 G.n2474 0.624
R9407 G.n2472 G.n2452 0.624
R9408 G.n2470 G.n2453 0.624
R9409 G.n2468 G.n2454 0.624
R9410 G.n2466 G.n2455 0.624
R9411 G.n2464 G.n2456 0.624
R9412 G.n2462 G.n2457 0.624
R9413 G.n2460 G.n2458 0.624
R9414 G.n2131 G.n2130 0.624
R9415 G.n2089 G.n2087 0.624
R9416 G.n2044 G.n2042 0.624
R9417 G.n1993 G.n1991 0.624
R9418 G.n1936 G.n1934 0.624
R9419 G.n1874 G.n1872 0.624
R9420 G.n1806 G.n1804 0.624
R9421 G.n1734 G.n1732 0.624
R9422 G.n1656 G.n1654 0.624
R9423 G.n1573 G.n1571 0.624
R9424 G.n1486 G.n1484 0.624
R9425 G.n1398 G.n1396 0.624
R9426 G.n1310 G.n1308 0.624
R9427 G.n1222 G.n1220 0.624
R9428 G.n1134 G.n1132 0.624
R9429 G.n1046 G.n1044 0.624
R9430 G.n961 G.n959 0.624
R9431 G.n879 G.n877 0.624
R9432 G.n803 G.n801 0.624
R9433 G.n730 G.n728 0.624
R9434 G.n660 G.n658 0.624
R9435 G.n593 G.n591 0.624
R9436 G.n529 G.n527 0.624
R9437 G.n468 G.n466 0.624
R9438 G.n410 G.n408 0.624
R9439 G.n355 G.n353 0.624
R9440 G.n306 G.n304 0.624
R9441 G.n260 G.n258 0.624
R9442 G.n3813 G.n3811 0.624
R9443 G.n3815 G.n3810 0.624
R9444 G.n3817 G.n3809 0.624
R9445 G.n3819 G.n3808 0.624
R9446 G.n3821 G.n3807 0.624
R9447 G.n3823 G.n3806 0.624
R9448 G.n3825 G.n3805 0.624
R9449 G.n3827 G.n3804 0.624
R9450 G.n3829 G.n3803 0.624
R9451 G.n3831 G.n3802 0.624
R9452 G.n3833 G.n3801 0.624
R9453 G.n3835 G.n3800 0.624
R9454 G.n3798 G.n3766 0.624
R9455 G.n3796 G.n3767 0.624
R9456 G.n3794 G.n3768 0.624
R9457 G.n3792 G.n3769 0.624
R9458 G.n3790 G.n3770 0.624
R9459 G.n3788 G.n3771 0.624
R9460 G.n3786 G.n3772 0.624
R9461 G.n3784 G.n3773 0.624
R9462 G.n3782 G.n3774 0.624
R9463 G.n3780 G.n3775 0.624
R9464 G.n3778 G.n3776 0.624
R9465 G.n220 G.n218 0.624
R9466 G.n263 G.n261 0.624
R9467 G.n309 G.n307 0.624
R9468 G.n358 G.n356 0.624
R9469 G.n413 G.n411 0.624
R9470 G.n471 G.n469 0.624
R9471 G.n532 G.n530 0.624
R9472 G.n596 G.n594 0.624
R9473 G.n663 G.n661 0.624
R9474 G.n733 G.n731 0.624
R9475 G.n806 G.n804 0.624
R9476 G.n882 G.n880 0.624
R9477 G.n964 G.n962 0.624
R9478 G.n1049 G.n1047 0.624
R9479 G.n1137 G.n1135 0.624
R9480 G.n1225 G.n1223 0.624
R9481 G.n1313 G.n1311 0.624
R9482 G.n1401 G.n1399 0.624
R9483 G.n1489 G.n1487 0.624
R9484 G.n1576 G.n1574 0.624
R9485 G.n1659 G.n1657 0.624
R9486 G.n1737 G.n1735 0.624
R9487 G.n1809 G.n1807 0.624
R9488 G.n1877 G.n1875 0.624
R9489 G.n1939 G.n1937 0.624
R9490 G.n1996 G.n1994 0.624
R9491 G.n2047 G.n2045 0.624
R9492 G.n2092 G.n2090 0.624
R9493 G.n2133 G.n2132 0.624
R9494 G.n2438 G.n2436 0.624
R9495 G.n2440 G.n2435 0.624
R9496 G.n2442 G.n2434 0.624
R9497 G.n2444 G.n2433 0.624
R9498 G.n2446 G.n2432 0.624
R9499 G.n2448 G.n2431 0.624
R9500 G.n2450 G.n2430 0.624
R9501 G.n2428 G.n2411 0.624
R9502 G.n2426 G.n2412 0.624
R9503 G.n2424 G.n2413 0.624
R9504 G.n2422 G.n2414 0.624
R9505 G.n2420 G.n2415 0.624
R9506 G.n2418 G.n2416 0.624
R9507 G.n2172 G.n2171 0.624
R9508 G.n2136 G.n2134 0.624
R9509 G.n2095 G.n2093 0.624
R9510 G.n2050 G.n2048 0.624
R9511 G.n1999 G.n1997 0.624
R9512 G.n1942 G.n1940 0.624
R9513 G.n1880 G.n1878 0.624
R9514 G.n1812 G.n1810 0.624
R9515 G.n1740 G.n1738 0.624
R9516 G.n1662 G.n1660 0.624
R9517 G.n1579 G.n1577 0.624
R9518 G.n1492 G.n1490 0.624
R9519 G.n1404 G.n1402 0.624
R9520 G.n1316 G.n1314 0.624
R9521 G.n1228 G.n1226 0.624
R9522 G.n1140 G.n1138 0.624
R9523 G.n1052 G.n1050 0.624
R9524 G.n967 G.n965 0.624
R9525 G.n885 G.n883 0.624
R9526 G.n809 G.n807 0.624
R9527 G.n736 G.n734 0.624
R9528 G.n666 G.n664 0.624
R9529 G.n599 G.n597 0.624
R9530 G.n535 G.n533 0.624
R9531 G.n474 G.n472 0.624
R9532 G.n416 G.n414 0.624
R9533 G.n361 G.n359 0.624
R9534 G.n312 G.n310 0.624
R9535 G.n266 G.n264 0.624
R9536 G.n223 G.n221 0.624
R9537 G.n183 G.n181 0.624
R9538 G.n3746 G.n3744 0.624
R9539 G.n3748 G.n3743 0.624
R9540 G.n3750 G.n3742 0.624
R9541 G.n3752 G.n3741 0.624
R9542 G.n3754 G.n3740 0.624
R9543 G.n3756 G.n3739 0.624
R9544 G.n3758 G.n3738 0.624
R9545 G.n3760 G.n3737 0.624
R9546 G.n3762 G.n3736 0.624
R9547 G.n3764 G.n3735 0.624
R9548 G.n3733 G.n3707 0.624
R9549 G.n3731 G.n3708 0.624
R9550 G.n3729 G.n3709 0.624
R9551 G.n3727 G.n3710 0.624
R9552 G.n3725 G.n3711 0.624
R9553 G.n3723 G.n3712 0.624
R9554 G.n3721 G.n3713 0.624
R9555 G.n3719 G.n3714 0.624
R9556 G.n3717 G.n3715 0.624
R9557 G.n149 G.n147 0.624
R9558 G.n186 G.n184 0.624
R9559 G.n226 G.n224 0.624
R9560 G.n269 G.n267 0.624
R9561 G.n315 G.n313 0.624
R9562 G.n364 G.n362 0.624
R9563 G.n419 G.n417 0.624
R9564 G.n477 G.n475 0.624
R9565 G.n538 G.n536 0.624
R9566 G.n602 G.n600 0.624
R9567 G.n669 G.n667 0.624
R9568 G.n739 G.n737 0.624
R9569 G.n812 G.n810 0.624
R9570 G.n888 G.n886 0.624
R9571 G.n970 G.n968 0.624
R9572 G.n1055 G.n1053 0.624
R9573 G.n1143 G.n1141 0.624
R9574 G.n1231 G.n1229 0.624
R9575 G.n1319 G.n1317 0.624
R9576 G.n1407 G.n1405 0.624
R9577 G.n1495 G.n1493 0.624
R9578 G.n1582 G.n1580 0.624
R9579 G.n1665 G.n1663 0.624
R9580 G.n1743 G.n1741 0.624
R9581 G.n1815 G.n1813 0.624
R9582 G.n1883 G.n1881 0.624
R9583 G.n1945 G.n1943 0.624
R9584 G.n2002 G.n2000 0.624
R9585 G.n2053 G.n2051 0.624
R9586 G.n2098 G.n2096 0.624
R9587 G.n2139 G.n2137 0.624
R9588 G.n2174 G.n2173 0.624
R9589 G.n2399 G.n2397 0.624
R9590 G.n2401 G.n2396 0.624
R9591 G.n2403 G.n2395 0.624
R9592 G.n2405 G.n2394 0.624
R9593 G.n2407 G.n2393 0.624
R9594 G.n2409 G.n2392 0.624
R9595 G.n2390 G.n2376 0.624
R9596 G.n2388 G.n2377 0.624
R9597 G.n2386 G.n2378 0.624
R9598 G.n2384 G.n2379 0.624
R9599 G.n2382 G.n2380 0.624
R9600 G.n2207 G.n2206 0.624
R9601 G.n2177 G.n2175 0.624
R9602 G.n2142 G.n2140 0.624
R9603 G.n2101 G.n2099 0.624
R9604 G.n2056 G.n2054 0.624
R9605 G.n2005 G.n2003 0.624
R9606 G.n1948 G.n1946 0.624
R9607 G.n1886 G.n1884 0.624
R9608 G.n1818 G.n1816 0.624
R9609 G.n1746 G.n1744 0.624
R9610 G.n1668 G.n1666 0.624
R9611 G.n1585 G.n1583 0.624
R9612 G.n1498 G.n1496 0.624
R9613 G.n1410 G.n1408 0.624
R9614 G.n1322 G.n1320 0.624
R9615 G.n1234 G.n1232 0.624
R9616 G.n1146 G.n1144 0.624
R9617 G.n1058 G.n1056 0.624
R9618 G.n973 G.n971 0.624
R9619 G.n891 G.n889 0.624
R9620 G.n815 G.n813 0.624
R9621 G.n742 G.n740 0.624
R9622 G.n672 G.n670 0.624
R9623 G.n605 G.n603 0.624
R9624 G.n541 G.n539 0.624
R9625 G.n480 G.n478 0.624
R9626 G.n422 G.n420 0.624
R9627 G.n367 G.n365 0.624
R9628 G.n318 G.n316 0.624
R9629 G.n272 G.n270 0.624
R9630 G.n229 G.n227 0.624
R9631 G.n189 G.n187 0.624
R9632 G.n152 G.n150 0.624
R9633 G.n118 G.n116 0.624
R9634 G.n3691 G.n3689 0.624
R9635 G.n3693 G.n3688 0.624
R9636 G.n3695 G.n3687 0.624
R9637 G.n3697 G.n3686 0.624
R9638 G.n3699 G.n3685 0.624
R9639 G.n3701 G.n3684 0.624
R9640 G.n3703 G.n3683 0.624
R9641 G.n3705 G.n3682 0.624
R9642 G.n3680 G.n3657 0.624
R9643 G.n3678 G.n3658 0.624
R9644 G.n3676 G.n3659 0.624
R9645 G.n3674 G.n3660 0.624
R9646 G.n3672 G.n3661 0.624
R9647 G.n3670 G.n3662 0.624
R9648 G.n3668 G.n3663 0.624
R9649 G.n3666 G.n3664 0.624
R9650 G.n121 G.n119 0.624
R9651 G.n155 G.n153 0.624
R9652 G.n192 G.n190 0.624
R9653 G.n232 G.n230 0.624
R9654 G.n275 G.n273 0.624
R9655 G.n321 G.n319 0.624
R9656 G.n370 G.n368 0.624
R9657 G.n425 G.n423 0.624
R9658 G.n483 G.n481 0.624
R9659 G.n544 G.n542 0.624
R9660 G.n608 G.n606 0.624
R9661 G.n675 G.n673 0.624
R9662 G.n745 G.n743 0.624
R9663 G.n818 G.n816 0.624
R9664 G.n894 G.n892 0.624
R9665 G.n976 G.n974 0.624
R9666 G.n1061 G.n1059 0.624
R9667 G.n1149 G.n1147 0.624
R9668 G.n1237 G.n1235 0.624
R9669 G.n1325 G.n1323 0.624
R9670 G.n1413 G.n1411 0.624
R9671 G.n1501 G.n1499 0.624
R9672 G.n1588 G.n1586 0.624
R9673 G.n1671 G.n1669 0.624
R9674 G.n1749 G.n1747 0.624
R9675 G.n1821 G.n1819 0.624
R9676 G.n1889 G.n1887 0.624
R9677 G.n1951 G.n1949 0.624
R9678 G.n2008 G.n2006 0.624
R9679 G.n2059 G.n2057 0.624
R9680 G.n2104 G.n2102 0.624
R9681 G.n2145 G.n2143 0.624
R9682 G.n2180 G.n2178 0.624
R9683 G.n2210 G.n2208 0.624
R9684 G.n2366 G.n2365 0.624
R9685 G.n2368 G.n2364 0.624
R9686 G.n2370 G.n2363 0.624
R9687 G.n2372 G.n2362 0.624
R9688 G.n2374 G.n2361 0.624
R9689 G.n2359 G.n2348 0.624
R9690 G.n2357 G.n2349 0.624
R9691 G.n2355 G.n2350 0.624
R9692 G.n2353 G.n2351 0.624
R9693 G.n2237 G.n2236 0.624
R9694 G.n2213 G.n2211 0.624
R9695 G.n2183 G.n2181 0.624
R9696 G.n2148 G.n2146 0.624
R9697 G.n2107 G.n2105 0.624
R9698 G.n2062 G.n2060 0.624
R9699 G.n2011 G.n2009 0.624
R9700 G.n1954 G.n1952 0.624
R9701 G.n1892 G.n1890 0.624
R9702 G.n1824 G.n1822 0.624
R9703 G.n1752 G.n1750 0.624
R9704 G.n1674 G.n1672 0.624
R9705 G.n1591 G.n1589 0.624
R9706 G.n1504 G.n1502 0.624
R9707 G.n1416 G.n1414 0.624
R9708 G.n1328 G.n1326 0.624
R9709 G.n1240 G.n1238 0.624
R9710 G.n1152 G.n1150 0.624
R9711 G.n1064 G.n1062 0.624
R9712 G.n979 G.n977 0.624
R9713 G.n897 G.n895 0.624
R9714 G.n821 G.n819 0.624
R9715 G.n748 G.n746 0.624
R9716 G.n678 G.n676 0.624
R9717 G.n611 G.n609 0.624
R9718 G.n547 G.n545 0.624
R9719 G.n486 G.n484 0.624
R9720 G.n428 G.n426 0.624
R9721 G.n373 G.n371 0.624
R9722 G.n324 G.n322 0.624
R9723 G.n278 G.n276 0.624
R9724 G.n235 G.n233 0.624
R9725 G.n195 G.n193 0.624
R9726 G.n158 G.n156 0.624
R9727 G.n124 G.n122 0.624
R9728 G.n93 G.n91 0.624
R9729 G.n3643 G.n3641 0.624
R9730 G.n3645 G.n3640 0.624
R9731 G.n3647 G.n3639 0.624
R9732 G.n3649 G.n3638 0.624
R9733 G.n3651 G.n3637 0.624
R9734 G.n3653 G.n3636 0.624
R9735 G.n3655 G.n3635 0.624
R9736 G.n3633 G.n3616 0.624
R9737 G.n3631 G.n3617 0.624
R9738 G.n3629 G.n3618 0.624
R9739 G.n3627 G.n3619 0.624
R9740 G.n3625 G.n3620 0.624
R9741 G.n3623 G.n3621 0.624
R9742 G.n71 G.n69 0.624
R9743 G.n96 G.n94 0.624
R9744 G.n127 G.n125 0.624
R9745 G.n161 G.n159 0.624
R9746 G.n198 G.n196 0.624
R9747 G.n238 G.n236 0.624
R9748 G.n281 G.n279 0.624
R9749 G.n327 G.n325 0.624
R9750 G.n376 G.n374 0.624
R9751 G.n431 G.n429 0.624
R9752 G.n489 G.n487 0.624
R9753 G.n550 G.n548 0.624
R9754 G.n614 G.n612 0.624
R9755 G.n681 G.n679 0.624
R9756 G.n751 G.n749 0.624
R9757 G.n824 G.n822 0.624
R9758 G.n900 G.n898 0.624
R9759 G.n982 G.n980 0.624
R9760 G.n1067 G.n1065 0.624
R9761 G.n1155 G.n1153 0.624
R9762 G.n1243 G.n1241 0.624
R9763 G.n1331 G.n1329 0.624
R9764 G.n1419 G.n1417 0.624
R9765 G.n1507 G.n1505 0.624
R9766 G.n1594 G.n1592 0.624
R9767 G.n1677 G.n1675 0.624
R9768 G.n1755 G.n1753 0.624
R9769 G.n1827 G.n1825 0.624
R9770 G.n1895 G.n1893 0.624
R9771 G.n1957 G.n1955 0.624
R9772 G.n2014 G.n2012 0.624
R9773 G.n2065 G.n2063 0.624
R9774 G.n2110 G.n2108 0.624
R9775 G.n2151 G.n2149 0.624
R9776 G.n2186 G.n2184 0.624
R9777 G.n2216 G.n2214 0.624
R9778 G.n2240 G.n2238 0.624
R9779 G.n2261 G.n2260 0.624
R9780 G.n2342 G.n2340 0.624
R9781 G.n2344 G.n2339 0.624
R9782 G.n2346 G.n2338 0.624
R9783 G.n2336 G.n2328 0.624
R9784 G.n2334 G.n2329 0.624
R9785 G.n2332 G.n2330 0.624
R9786 G.n2263 G.n2262 0.624
R9787 G.n2243 G.n2241 0.624
R9788 G.n2219 G.n2217 0.624
R9789 G.n2189 G.n2187 0.624
R9790 G.n2154 G.n2152 0.624
R9791 G.n2113 G.n2111 0.624
R9792 G.n2068 G.n2066 0.624
R9793 G.n2017 G.n2015 0.624
R9794 G.n1960 G.n1958 0.624
R9795 G.n1898 G.n1896 0.624
R9796 G.n1830 G.n1828 0.624
R9797 G.n1758 G.n1756 0.624
R9798 G.n1680 G.n1678 0.624
R9799 G.n1597 G.n1595 0.624
R9800 G.n1510 G.n1508 0.624
R9801 G.n1422 G.n1420 0.624
R9802 G.n1334 G.n1332 0.624
R9803 G.n1246 G.n1244 0.624
R9804 G.n1158 G.n1156 0.624
R9805 G.n1070 G.n1068 0.624
R9806 G.n985 G.n983 0.624
R9807 G.n903 G.n901 0.624
R9808 G.n827 G.n825 0.624
R9809 G.n754 G.n752 0.624
R9810 G.n684 G.n682 0.624
R9811 G.n617 G.n615 0.624
R9812 G.n553 G.n551 0.624
R9813 G.n492 G.n490 0.624
R9814 G.n434 G.n432 0.624
R9815 G.n379 G.n377 0.624
R9816 G.n330 G.n328 0.624
R9817 G.n284 G.n282 0.624
R9818 G.n241 G.n239 0.624
R9819 G.n201 G.n199 0.624
R9820 G.n164 G.n162 0.624
R9821 G.n130 G.n128 0.624
R9822 G.n99 G.n97 0.624
R9823 G.n74 G.n72 0.624
R9824 G.n52 G.n50 0.624
R9825 G.n3606 G.n3604 0.624
R9826 G.n3608 G.n3603 0.624
R9827 G.n3610 G.n3602 0.624
R9828 G.n3612 G.n3601 0.624
R9829 G.n3614 G.n3600 0.624
R9830 G.n3598 G.n3587 0.624
R9831 G.n3596 G.n3588 0.624
R9832 G.n3594 G.n3589 0.624
R9833 G.n3592 G.n3590 0.624
R9834 G.n36 G.n34 0.624
R9835 G.n55 G.n53 0.624
R9836 G.n77 G.n75 0.624
R9837 G.n102 G.n100 0.624
R9838 G.n133 G.n131 0.624
R9839 G.n167 G.n165 0.624
R9840 G.n204 G.n202 0.624
R9841 G.n244 G.n242 0.624
R9842 G.n287 G.n285 0.624
R9843 G.n333 G.n331 0.624
R9844 G.n382 G.n380 0.624
R9845 G.n437 G.n435 0.624
R9846 G.n495 G.n493 0.624
R9847 G.n556 G.n554 0.624
R9848 G.n620 G.n618 0.624
R9849 G.n687 G.n685 0.624
R9850 G.n757 G.n755 0.624
R9851 G.n830 G.n828 0.624
R9852 G.n906 G.n904 0.624
R9853 G.n988 G.n986 0.624
R9854 G.n1073 G.n1071 0.624
R9855 G.n1161 G.n1159 0.624
R9856 G.n1249 G.n1247 0.624
R9857 G.n1337 G.n1335 0.624
R9858 G.n1425 G.n1423 0.624
R9859 G.n1513 G.n1511 0.624
R9860 G.n1600 G.n1598 0.624
R9861 G.n1683 G.n1681 0.624
R9862 G.n1761 G.n1759 0.624
R9863 G.n1833 G.n1831 0.624
R9864 G.n1901 G.n1899 0.624
R9865 G.n1963 G.n1961 0.624
R9866 G.n2020 G.n2018 0.624
R9867 G.n2071 G.n2069 0.624
R9868 G.n2116 G.n2114 0.624
R9869 G.n2157 G.n2155 0.624
R9870 G.n2192 G.n2190 0.624
R9871 G.n2222 G.n2220 0.624
R9872 G.n2246 G.n2244 0.624
R9873 G.n2266 G.n2264 0.624
R9874 G.n2281 G.n2280 0.624
R9875 G.n2324 G.n2322 0.624
R9876 G.n2326 G.n2321 0.624
R9877 G.n2319 G.n2314 0.624
R9878 G.n2317 G.n2315 0.624
R9879 G.n2283 G.n2282 0.624
R9880 G.n2269 G.n2267 0.624
R9881 G.n2249 G.n2247 0.624
R9882 G.n2225 G.n2223 0.624
R9883 G.n2195 G.n2193 0.624
R9884 G.n2160 G.n2158 0.624
R9885 G.n2119 G.n2117 0.624
R9886 G.n2074 G.n2072 0.624
R9887 G.n2023 G.n2021 0.624
R9888 G.n1966 G.n1964 0.624
R9889 G.n1904 G.n1902 0.624
R9890 G.n1836 G.n1834 0.624
R9891 G.n1764 G.n1762 0.624
R9892 G.n1686 G.n1684 0.624
R9893 G.n1603 G.n1601 0.624
R9894 G.n1516 G.n1514 0.624
R9895 G.n1428 G.n1426 0.624
R9896 G.n1340 G.n1338 0.624
R9897 G.n1252 G.n1250 0.624
R9898 G.n1164 G.n1162 0.624
R9899 G.n1076 G.n1074 0.624
R9900 G.n991 G.n989 0.624
R9901 G.n909 G.n907 0.624
R9902 G.n833 G.n831 0.624
R9903 G.n760 G.n758 0.624
R9904 G.n690 G.n688 0.624
R9905 G.n623 G.n621 0.624
R9906 G.n559 G.n557 0.624
R9907 G.n498 G.n496 0.624
R9908 G.n440 G.n438 0.624
R9909 G.n385 G.n383 0.624
R9910 G.n336 G.n334 0.624
R9911 G.n290 G.n288 0.624
R9912 G.n247 G.n245 0.624
R9913 G.n207 G.n205 0.624
R9914 G.n170 G.n168 0.624
R9915 G.n136 G.n134 0.624
R9916 G.n105 G.n103 0.624
R9917 G.n80 G.n78 0.624
R9918 G.n58 G.n56 0.624
R9919 G.n39 G.n37 0.624
R9920 G.n23 G.n21 0.624
R9921 G.n3581 G.n3579 0.624
R9922 G.n3583 G.n3578 0.624
R9923 G.n3585 G.n3577 0.624
R9924 G.n3575 G.n3570 0.624
R9925 G.n3573 G.n3571 0.624
R9926 G.n13 G.n11 0.624
R9927 G.n26 G.n24 0.624
R9928 G.n42 G.n40 0.624
R9929 G.n61 G.n59 0.624
R9930 G.n83 G.n81 0.624
R9931 G.n108 G.n106 0.624
R9932 G.n139 G.n137 0.624
R9933 G.n173 G.n171 0.624
R9934 G.n210 G.n208 0.624
R9935 G.n250 G.n248 0.624
R9936 G.n293 G.n291 0.624
R9937 G.n339 G.n337 0.624
R9938 G.n388 G.n386 0.624
R9939 G.n443 G.n441 0.624
R9940 G.n501 G.n499 0.624
R9941 G.n562 G.n560 0.624
R9942 G.n626 G.n624 0.624
R9943 G.n693 G.n691 0.624
R9944 G.n763 G.n761 0.624
R9945 G.n836 G.n834 0.624
R9946 G.n912 G.n910 0.624
R9947 G.n994 G.n992 0.624
R9948 G.n1079 G.n1077 0.624
R9949 G.n1167 G.n1165 0.624
R9950 G.n1255 G.n1253 0.624
R9951 G.n1343 G.n1341 0.624
R9952 G.n1431 G.n1429 0.624
R9953 G.n1519 G.n1517 0.624
R9954 G.n1606 G.n1604 0.624
R9955 G.n1689 G.n1687 0.624
R9956 G.n1767 G.n1765 0.624
R9957 G.n1839 G.n1837 0.624
R9958 G.n1907 G.n1905 0.624
R9959 G.n1969 G.n1967 0.624
R9960 G.n2026 G.n2024 0.624
R9961 G.n2077 G.n2075 0.624
R9962 G.n2122 G.n2120 0.624
R9963 G.n2163 G.n2161 0.624
R9964 G.n2198 G.n2196 0.624
R9965 G.n2228 G.n2226 0.624
R9966 G.n2252 G.n2250 0.624
R9967 G.n2272 G.n2270 0.624
R9968 G.n2286 G.n2284 0.624
R9969 G.n2295 G.n2294 0.624
R9970 G.n2312 G.n2310 0.624
R9971 G.n2308 G.n2307 0.624
R9972 G.n2298 G.n2296 0.624
R9973 G.n2289 G.n2287 0.624
R9974 G.n2275 G.n2273 0.624
R9975 G.n2255 G.n2253 0.624
R9976 G.n2231 G.n2229 0.624
R9977 G.n2201 G.n2199 0.624
R9978 G.n2166 G.n2164 0.624
R9979 G.n2125 G.n2123 0.624
R9980 G.n2080 G.n2078 0.624
R9981 G.n2029 G.n2027 0.624
R9982 G.n1972 G.n1970 0.624
R9983 G.n1910 G.n1908 0.624
R9984 G.n1842 G.n1840 0.624
R9985 G.n1770 G.n1768 0.624
R9986 G.n1692 G.n1690 0.624
R9987 G.n1609 G.n1607 0.624
R9988 G.n1522 G.n1520 0.624
R9989 G.n1434 G.n1432 0.624
R9990 G.n1346 G.n1344 0.624
R9991 G.n1258 G.n1256 0.624
R9992 G.n1170 G.n1168 0.624
R9993 G.n1082 G.n1080 0.624
R9994 G.n997 G.n995 0.624
R9995 G.n915 G.n913 0.624
R9996 G.n839 G.n837 0.624
R9997 G.n766 G.n764 0.624
R9998 G.n696 G.n694 0.624
R9999 G.n629 G.n627 0.624
R10000 G.n565 G.n563 0.624
R10001 G.n504 G.n502 0.624
R10002 G.n446 G.n444 0.624
R10003 G.n391 G.n389 0.624
R10004 G.n342 G.n340 0.624
R10005 G.n296 G.n294 0.624
R10006 G.n253 G.n251 0.624
R10007 G.n213 G.n211 0.624
R10008 G.n176 G.n174 0.624
R10009 G.n142 G.n140 0.624
R10010 G.n111 G.n109 0.624
R10011 G.n86 G.n84 0.624
R10012 G.n64 G.n62 0.624
R10013 G.n45 G.n43 0.624
R10014 G.n29 G.n27 0.624
R10015 G.n16 G.n14 0.624
R10016 G.n6 G.n4 0.624
R10017 G.n3568 G.n3566 0.624
R10018 G.n3 G.n2 0.624
R10019 G.n2 G.n0 0.624
R10020 G.n10 G.n9 0.624
R10021 G.n9 G.n7 0.624
R10022 G.n20 G.n19 0.624
R10023 G.n19 G.n17 0.624
R10024 G.n33 G.n32 0.624
R10025 G.n32 G.n30 0.624
R10026 G.n49 G.n48 0.624
R10027 G.n48 G.n46 0.624
R10028 G.n68 G.n67 0.624
R10029 G.n67 G.n65 0.624
R10030 G.n90 G.n89 0.624
R10031 G.n89 G.n87 0.624
R10032 G.n115 G.n114 0.624
R10033 G.n114 G.n112 0.624
R10034 G.n146 G.n145 0.624
R10035 G.n145 G.n143 0.624
R10036 G.n180 G.n179 0.624
R10037 G.n179 G.n177 0.624
R10038 G.n217 G.n216 0.624
R10039 G.n216 G.n214 0.624
R10040 G.n257 G.n256 0.624
R10041 G.n256 G.n254 0.624
R10042 G.n300 G.n299 0.624
R10043 G.n299 G.n297 0.624
R10044 G.n346 G.n345 0.624
R10045 G.n345 G.n343 0.624
R10046 G.n395 G.n394 0.624
R10047 G.n394 G.n392 0.624
R10048 G.n450 G.n449 0.624
R10049 G.n449 G.n447 0.624
R10050 G.n508 G.n507 0.624
R10051 G.n507 G.n505 0.624
R10052 G.n569 G.n568 0.624
R10053 G.n568 G.n566 0.624
R10054 G.n633 G.n632 0.624
R10055 G.n632 G.n630 0.624
R10056 G.n700 G.n699 0.624
R10057 G.n699 G.n697 0.624
R10058 G.n770 G.n769 0.624
R10059 G.n769 G.n767 0.624
R10060 G.n843 G.n842 0.624
R10061 G.n842 G.n840 0.624
R10062 G.n919 G.n918 0.624
R10063 G.n918 G.n916 0.624
R10064 G.n1001 G.n1000 0.624
R10065 G.n1000 G.n998 0.624
R10066 G.n1086 G.n1085 0.624
R10067 G.n1085 G.n1083 0.624
R10068 G.n1174 G.n1173 0.624
R10069 G.n1173 G.n1171 0.624
R10070 G.n1262 G.n1261 0.624
R10071 G.n1261 G.n1259 0.624
R10072 G.n1350 G.n1349 0.624
R10073 G.n1349 G.n1347 0.624
R10074 G.n1438 G.n1437 0.624
R10075 G.n1437 G.n1435 0.624
R10076 G.n1526 G.n1525 0.624
R10077 G.n1525 G.n1523 0.624
R10078 G.n1613 G.n1612 0.624
R10079 G.n1612 G.n1610 0.624
R10080 G.n1696 G.n1695 0.624
R10081 G.n1695 G.n1693 0.624
R10082 G.n1774 G.n1773 0.624
R10083 G.n1773 G.n1771 0.624
R10084 G.n1846 G.n1845 0.624
R10085 G.n1845 G.n1843 0.624
R10086 G.n1914 G.n1913 0.624
R10087 G.n1913 G.n1911 0.624
R10088 G.n1976 G.n1975 0.624
R10089 G.n1975 G.n1973 0.624
R10090 G.n2033 G.n2032 0.624
R10091 G.n2032 G.n2030 0.624
R10092 G.n2084 G.n2083 0.624
R10093 G.n2083 G.n2081 0.624
R10094 G.n2129 G.n2128 0.624
R10095 G.n2128 G.n2126 0.624
R10096 G.n2170 G.n2169 0.624
R10097 G.n2169 G.n2167 0.624
R10098 G.n2205 G.n2204 0.624
R10099 G.n2204 G.n2202 0.624
R10100 G.n2235 G.n2234 0.624
R10101 G.n2234 G.n2232 0.624
R10102 G.n2259 G.n2258 0.624
R10103 G.n2258 G.n2256 0.624
R10104 G.n2279 G.n2278 0.624
R10105 G.n2278 G.n2276 0.624
R10106 G.n2293 G.n2292 0.624
R10107 G.n2292 G.n2290 0.624
R10108 G.n2302 G.n2301 0.624
R10109 G.n2301 G.n2299 0.624
R10110 G.n2305 G.n2304 0.624
R10111 G.n2304 G.n2303 0.624
R10112 G.n3518 G.n2305 0.624
R10113 G.n3519 G.n2302 0.624
R10114 G.n3520 G.n2293 0.624
R10115 G.n3521 G.n2279 0.624
R10116 G.n3522 G.n2259 0.624
R10117 G.n3523 G.n2235 0.624
R10118 G.n3524 G.n2205 0.624
R10119 G.n3525 G.n2170 0.624
R10120 G.n3526 G.n2129 0.624
R10121 G.n3527 G.n2084 0.624
R10122 G.n3528 G.n2033 0.624
R10123 G.n3529 G.n1976 0.624
R10124 G.n3530 G.n1914 0.624
R10125 G.n3531 G.n1846 0.624
R10126 G.n3532 G.n1774 0.624
R10127 G.n3533 G.n1696 0.624
R10128 G.n3534 G.n1613 0.624
R10129 G.n3535 G.n1526 0.624
R10130 G.n3536 G.n1438 0.624
R10131 G.n3537 G.n1350 0.624
R10132 G.n3538 G.n1262 0.624
R10133 G.n3539 G.n1174 0.624
R10134 G.n3540 G.n1086 0.624
R10135 G.n3541 G.n1001 0.624
R10136 G.n3542 G.n919 0.624
R10137 G.n3543 G.n843 0.624
R10138 G.n3544 G.n770 0.624
R10139 G.n3545 G.n700 0.624
R10140 G.n3546 G.n633 0.624
R10141 G.n3547 G.n569 0.624
R10142 G.n3548 G.n508 0.624
R10143 G.n3549 G.n450 0.624
R10144 G.n3550 G.n395 0.624
R10145 G.n3551 G.n346 0.624
R10146 G.n3552 G.n300 0.624
R10147 G.n3553 G.n257 0.624
R10148 G.n3554 G.n217 0.624
R10149 G.n3555 G.n180 0.624
R10150 G.n3556 G.n146 0.624
R10151 G.n3557 G.n115 0.624
R10152 G.n3558 G.n90 0.624
R10153 G.n3559 G.n68 0.624
R10154 G.n3560 G.n49 0.624
R10155 G.n3561 G.n33 0.624
R10156 G.n3562 G.n20 0.624
R10157 G.n3563 G.n10 0.624
R10158 G.n2299 G.n2298 0.624
R10159 G.n2290 G.n2289 0.624
R10160 G.n2276 G.n2275 0.624
R10161 G.n2256 G.n2255 0.624
R10162 G.n2232 G.n2231 0.624
R10163 G.n2202 G.n2201 0.624
R10164 G.n2167 G.n2166 0.624
R10165 G.n2126 G.n2125 0.624
R10166 G.n2081 G.n2080 0.624
R10167 G.n2030 G.n2029 0.624
R10168 G.n1973 G.n1972 0.624
R10169 G.n1911 G.n1910 0.624
R10170 G.n1843 G.n1842 0.624
R10171 G.n1771 G.n1770 0.624
R10172 G.n1693 G.n1692 0.624
R10173 G.n1610 G.n1609 0.624
R10174 G.n1523 G.n1522 0.624
R10175 G.n1435 G.n1434 0.624
R10176 G.n1347 G.n1346 0.624
R10177 G.n1259 G.n1258 0.624
R10178 G.n1171 G.n1170 0.624
R10179 G.n1083 G.n1082 0.624
R10180 G.n998 G.n997 0.624
R10181 G.n916 G.n915 0.624
R10182 G.n840 G.n839 0.624
R10183 G.n767 G.n766 0.624
R10184 G.n697 G.n696 0.624
R10185 G.n630 G.n629 0.624
R10186 G.n566 G.n565 0.624
R10187 G.n505 G.n504 0.624
R10188 G.n447 G.n446 0.624
R10189 G.n392 G.n391 0.624
R10190 G.n343 G.n342 0.624
R10191 G.n297 G.n296 0.624
R10192 G.n254 G.n253 0.624
R10193 G.n214 G.n213 0.624
R10194 G.n177 G.n176 0.624
R10195 G.n143 G.n142 0.624
R10196 G.n112 G.n111 0.624
R10197 G.n87 G.n86 0.624
R10198 G.n65 G.n64 0.624
R10199 G.n46 G.n45 0.624
R10200 G.n30 G.n29 0.624
R10201 G.n17 G.n16 0.624
R10202 G.n2287 G.n2286 0.624
R10203 G.n2273 G.n2272 0.624
R10204 G.n2253 G.n2252 0.624
R10205 G.n2229 G.n2228 0.624
R10206 G.n2199 G.n2198 0.624
R10207 G.n2164 G.n2163 0.624
R10208 G.n2123 G.n2122 0.624
R10209 G.n2078 G.n2077 0.624
R10210 G.n2027 G.n2026 0.624
R10211 G.n1970 G.n1969 0.624
R10212 G.n1908 G.n1907 0.624
R10213 G.n1840 G.n1839 0.624
R10214 G.n1768 G.n1767 0.624
R10215 G.n1690 G.n1689 0.624
R10216 G.n1607 G.n1606 0.624
R10217 G.n1520 G.n1519 0.624
R10218 G.n1432 G.n1431 0.624
R10219 G.n1344 G.n1343 0.624
R10220 G.n1256 G.n1255 0.624
R10221 G.n1168 G.n1167 0.624
R10222 G.n1080 G.n1079 0.624
R10223 G.n995 G.n994 0.624
R10224 G.n913 G.n912 0.624
R10225 G.n837 G.n836 0.624
R10226 G.n764 G.n763 0.624
R10227 G.n694 G.n693 0.624
R10228 G.n627 G.n626 0.624
R10229 G.n563 G.n562 0.624
R10230 G.n502 G.n501 0.624
R10231 G.n444 G.n443 0.624
R10232 G.n389 G.n388 0.624
R10233 G.n340 G.n339 0.624
R10234 G.n294 G.n293 0.624
R10235 G.n251 G.n250 0.624
R10236 G.n211 G.n210 0.624
R10237 G.n174 G.n173 0.624
R10238 G.n140 G.n139 0.624
R10239 G.n109 G.n108 0.624
R10240 G.n84 G.n83 0.624
R10241 G.n62 G.n61 0.624
R10242 G.n43 G.n42 0.624
R10243 G.n27 G.n26 0.624
R10244 G.n14 G.n13 0.624
R10245 G.n2270 G.n2269 0.624
R10246 G.n2250 G.n2249 0.624
R10247 G.n2226 G.n2225 0.624
R10248 G.n2196 G.n2195 0.624
R10249 G.n2161 G.n2160 0.624
R10250 G.n2120 G.n2119 0.624
R10251 G.n2075 G.n2074 0.624
R10252 G.n2024 G.n2023 0.624
R10253 G.n1967 G.n1966 0.624
R10254 G.n1905 G.n1904 0.624
R10255 G.n1837 G.n1836 0.624
R10256 G.n1765 G.n1764 0.624
R10257 G.n1687 G.n1686 0.624
R10258 G.n1604 G.n1603 0.624
R10259 G.n1517 G.n1516 0.624
R10260 G.n1429 G.n1428 0.624
R10261 G.n1341 G.n1340 0.624
R10262 G.n1253 G.n1252 0.624
R10263 G.n1165 G.n1164 0.624
R10264 G.n1077 G.n1076 0.624
R10265 G.n992 G.n991 0.624
R10266 G.n910 G.n909 0.624
R10267 G.n834 G.n833 0.624
R10268 G.n761 G.n760 0.624
R10269 G.n691 G.n690 0.624
R10270 G.n624 G.n623 0.624
R10271 G.n560 G.n559 0.624
R10272 G.n499 G.n498 0.624
R10273 G.n441 G.n440 0.624
R10274 G.n386 G.n385 0.624
R10275 G.n337 G.n336 0.624
R10276 G.n291 G.n290 0.624
R10277 G.n248 G.n247 0.624
R10278 G.n208 G.n207 0.624
R10279 G.n171 G.n170 0.624
R10280 G.n137 G.n136 0.624
R10281 G.n106 G.n105 0.624
R10282 G.n81 G.n80 0.624
R10283 G.n59 G.n58 0.624
R10284 G.n40 G.n39 0.624
R10285 G.n24 G.n23 0.624
R10286 G.n2267 G.n2266 0.624
R10287 G.n2223 G.n2222 0.624
R10288 G.n2193 G.n2192 0.624
R10289 G.n2158 G.n2157 0.624
R10290 G.n2117 G.n2116 0.624
R10291 G.n2072 G.n2071 0.624
R10292 G.n2021 G.n2020 0.624
R10293 G.n1964 G.n1963 0.624
R10294 G.n1902 G.n1901 0.624
R10295 G.n1834 G.n1833 0.624
R10296 G.n1762 G.n1761 0.624
R10297 G.n1684 G.n1683 0.624
R10298 G.n1601 G.n1600 0.624
R10299 G.n1514 G.n1513 0.624
R10300 G.n1426 G.n1425 0.624
R10301 G.n1338 G.n1337 0.624
R10302 G.n1250 G.n1249 0.624
R10303 G.n1162 G.n1161 0.624
R10304 G.n1074 G.n1073 0.624
R10305 G.n989 G.n988 0.624
R10306 G.n907 G.n906 0.624
R10307 G.n831 G.n830 0.624
R10308 G.n758 G.n757 0.624
R10309 G.n688 G.n687 0.624
R10310 G.n621 G.n620 0.624
R10311 G.n557 G.n556 0.624
R10312 G.n496 G.n495 0.624
R10313 G.n438 G.n437 0.624
R10314 G.n383 G.n382 0.624
R10315 G.n334 G.n333 0.624
R10316 G.n288 G.n287 0.624
R10317 G.n245 G.n244 0.624
R10318 G.n205 G.n204 0.624
R10319 G.n168 G.n167 0.624
R10320 G.n134 G.n133 0.624
R10321 G.n103 G.n102 0.624
R10322 G.n78 G.n77 0.624
R10323 G.n56 G.n55 0.624
R10324 G.n37 G.n36 0.624
R10325 G.n2247 G.n2246 0.624
R10326 G.n2264 G.n2263 0.624
R10327 G.n2190 G.n2189 0.624
R10328 G.n2155 G.n2154 0.624
R10329 G.n2114 G.n2113 0.624
R10330 G.n2069 G.n2068 0.624
R10331 G.n2018 G.n2017 0.624
R10332 G.n1961 G.n1960 0.624
R10333 G.n1899 G.n1898 0.624
R10334 G.n1831 G.n1830 0.624
R10335 G.n1759 G.n1758 0.624
R10336 G.n1681 G.n1680 0.624
R10337 G.n1598 G.n1597 0.624
R10338 G.n1511 G.n1510 0.624
R10339 G.n1423 G.n1422 0.624
R10340 G.n1335 G.n1334 0.624
R10341 G.n1247 G.n1246 0.624
R10342 G.n1159 G.n1158 0.624
R10343 G.n1071 G.n1070 0.624
R10344 G.n986 G.n985 0.624
R10345 G.n904 G.n903 0.624
R10346 G.n828 G.n827 0.624
R10347 G.n755 G.n754 0.624
R10348 G.n685 G.n684 0.624
R10349 G.n618 G.n617 0.624
R10350 G.n554 G.n553 0.624
R10351 G.n493 G.n492 0.624
R10352 G.n435 G.n434 0.624
R10353 G.n380 G.n379 0.624
R10354 G.n331 G.n330 0.624
R10355 G.n285 G.n284 0.624
R10356 G.n242 G.n241 0.624
R10357 G.n202 G.n201 0.624
R10358 G.n165 G.n164 0.624
R10359 G.n131 G.n130 0.624
R10360 G.n100 G.n99 0.624
R10361 G.n75 G.n74 0.624
R10362 G.n53 G.n52 0.624
R10363 G.n2220 G.n2219 0.624
R10364 G.n2244 G.n2243 0.624
R10365 G.n2262 G.n2261 0.624
R10366 G.n2187 G.n2186 0.624
R10367 G.n2111 G.n2110 0.624
R10368 G.n2066 G.n2065 0.624
R10369 G.n2015 G.n2014 0.624
R10370 G.n1958 G.n1957 0.624
R10371 G.n1896 G.n1895 0.624
R10372 G.n1828 G.n1827 0.624
R10373 G.n1756 G.n1755 0.624
R10374 G.n1678 G.n1677 0.624
R10375 G.n1595 G.n1594 0.624
R10376 G.n1508 G.n1507 0.624
R10377 G.n1420 G.n1419 0.624
R10378 G.n1332 G.n1331 0.624
R10379 G.n1244 G.n1243 0.624
R10380 G.n1156 G.n1155 0.624
R10381 G.n1068 G.n1067 0.624
R10382 G.n983 G.n982 0.624
R10383 G.n901 G.n900 0.624
R10384 G.n825 G.n824 0.624
R10385 G.n752 G.n751 0.624
R10386 G.n682 G.n681 0.624
R10387 G.n615 G.n614 0.624
R10388 G.n551 G.n550 0.624
R10389 G.n490 G.n489 0.624
R10390 G.n432 G.n431 0.624
R10391 G.n377 G.n376 0.624
R10392 G.n328 G.n327 0.624
R10393 G.n282 G.n281 0.624
R10394 G.n239 G.n238 0.624
R10395 G.n199 G.n198 0.624
R10396 G.n162 G.n161 0.624
R10397 G.n128 G.n127 0.624
R10398 G.n97 G.n96 0.624
R10399 G.n72 G.n71 0.624
R10400 G.n2152 G.n2151 0.624
R10401 G.n2217 G.n2216 0.624
R10402 G.n2241 G.n2240 0.624
R10403 G.n2184 G.n2183 0.624
R10404 G.n2063 G.n2062 0.624
R10405 G.n2012 G.n2011 0.624
R10406 G.n1955 G.n1954 0.624
R10407 G.n1893 G.n1892 0.624
R10408 G.n1825 G.n1824 0.624
R10409 G.n1753 G.n1752 0.624
R10410 G.n1675 G.n1674 0.624
R10411 G.n1592 G.n1591 0.624
R10412 G.n1505 G.n1504 0.624
R10413 G.n1417 G.n1416 0.624
R10414 G.n1329 G.n1328 0.624
R10415 G.n1241 G.n1240 0.624
R10416 G.n1153 G.n1152 0.624
R10417 G.n1065 G.n1064 0.624
R10418 G.n980 G.n979 0.624
R10419 G.n898 G.n897 0.624
R10420 G.n822 G.n821 0.624
R10421 G.n749 G.n748 0.624
R10422 G.n679 G.n678 0.624
R10423 G.n612 G.n611 0.624
R10424 G.n548 G.n547 0.624
R10425 G.n487 G.n486 0.624
R10426 G.n429 G.n428 0.624
R10427 G.n374 G.n373 0.624
R10428 G.n325 G.n324 0.624
R10429 G.n279 G.n278 0.624
R10430 G.n236 G.n235 0.624
R10431 G.n196 G.n195 0.624
R10432 G.n159 G.n158 0.624
R10433 G.n125 G.n124 0.624
R10434 G.n94 G.n93 0.624
R10435 G.n2108 G.n2107 0.624
R10436 G.n2149 G.n2148 0.624
R10437 G.n2214 G.n2213 0.624
R10438 G.n2238 G.n2237 0.624
R10439 G.n2181 G.n2180 0.624
R10440 G.n2060 G.n2059 0.624
R10441 G.n1952 G.n1951 0.624
R10442 G.n1890 G.n1889 0.624
R10443 G.n1822 G.n1821 0.624
R10444 G.n1750 G.n1749 0.624
R10445 G.n1672 G.n1671 0.624
R10446 G.n1589 G.n1588 0.624
R10447 G.n1502 G.n1501 0.624
R10448 G.n1414 G.n1413 0.624
R10449 G.n1326 G.n1325 0.624
R10450 G.n1238 G.n1237 0.624
R10451 G.n1150 G.n1149 0.624
R10452 G.n1062 G.n1061 0.624
R10453 G.n977 G.n976 0.624
R10454 G.n895 G.n894 0.624
R10455 G.n819 G.n818 0.624
R10456 G.n746 G.n745 0.624
R10457 G.n676 G.n675 0.624
R10458 G.n609 G.n608 0.624
R10459 G.n545 G.n544 0.624
R10460 G.n484 G.n483 0.624
R10461 G.n426 G.n425 0.624
R10462 G.n371 G.n370 0.624
R10463 G.n322 G.n321 0.624
R10464 G.n276 G.n275 0.624
R10465 G.n233 G.n232 0.624
R10466 G.n193 G.n192 0.624
R10467 G.n156 G.n155 0.624
R10468 G.n122 G.n121 0.624
R10469 G.n2009 G.n2008 0.624
R10470 G.n2105 G.n2104 0.624
R10471 G.n2146 G.n2145 0.624
R10472 G.n2211 G.n2210 0.624
R10473 G.n2178 G.n2177 0.624
R10474 G.n2057 G.n2056 0.624
R10475 G.n1887 G.n1886 0.624
R10476 G.n1819 G.n1818 0.624
R10477 G.n1747 G.n1746 0.624
R10478 G.n1669 G.n1668 0.624
R10479 G.n1586 G.n1585 0.624
R10480 G.n1499 G.n1498 0.624
R10481 G.n1411 G.n1410 0.624
R10482 G.n1323 G.n1322 0.624
R10483 G.n1235 G.n1234 0.624
R10484 G.n1147 G.n1146 0.624
R10485 G.n1059 G.n1058 0.624
R10486 G.n974 G.n973 0.624
R10487 G.n892 G.n891 0.624
R10488 G.n816 G.n815 0.624
R10489 G.n743 G.n742 0.624
R10490 G.n673 G.n672 0.624
R10491 G.n606 G.n605 0.624
R10492 G.n542 G.n541 0.624
R10493 G.n481 G.n480 0.624
R10494 G.n423 G.n422 0.624
R10495 G.n368 G.n367 0.624
R10496 G.n319 G.n318 0.624
R10497 G.n273 G.n272 0.624
R10498 G.n230 G.n229 0.624
R10499 G.n190 G.n189 0.624
R10500 G.n153 G.n152 0.624
R10501 G.n119 G.n118 0.624
R10502 G.n1949 G.n1948 0.624
R10503 G.n2006 G.n2005 0.624
R10504 G.n2102 G.n2101 0.624
R10505 G.n2143 G.n2142 0.624
R10506 G.n2208 G.n2207 0.624
R10507 G.n2175 G.n2174 0.624
R10508 G.n2054 G.n2053 0.624
R10509 G.n1884 G.n1883 0.624
R10510 G.n1744 G.n1743 0.624
R10511 G.n1666 G.n1665 0.624
R10512 G.n1583 G.n1582 0.624
R10513 G.n1496 G.n1495 0.624
R10514 G.n1408 G.n1407 0.624
R10515 G.n1320 G.n1319 0.624
R10516 G.n1232 G.n1231 0.624
R10517 G.n1144 G.n1143 0.624
R10518 G.n1056 G.n1055 0.624
R10519 G.n971 G.n970 0.624
R10520 G.n889 G.n888 0.624
R10521 G.n813 G.n812 0.624
R10522 G.n740 G.n739 0.624
R10523 G.n670 G.n669 0.624
R10524 G.n603 G.n602 0.624
R10525 G.n539 G.n538 0.624
R10526 G.n478 G.n477 0.624
R10527 G.n420 G.n419 0.624
R10528 G.n365 G.n364 0.624
R10529 G.n316 G.n315 0.624
R10530 G.n270 G.n269 0.624
R10531 G.n227 G.n226 0.624
R10532 G.n187 G.n186 0.624
R10533 G.n150 G.n149 0.624
R10534 G.n1816 G.n1815 0.624
R10535 G.n1946 G.n1945 0.624
R10536 G.n2003 G.n2002 0.624
R10537 G.n2099 G.n2098 0.624
R10538 G.n2140 G.n2139 0.624
R10539 G.n2173 G.n2172 0.624
R10540 G.n2051 G.n2050 0.624
R10541 G.n1881 G.n1880 0.624
R10542 G.n1663 G.n1662 0.624
R10543 G.n1580 G.n1579 0.624
R10544 G.n1493 G.n1492 0.624
R10545 G.n1405 G.n1404 0.624
R10546 G.n1317 G.n1316 0.624
R10547 G.n1229 G.n1228 0.624
R10548 G.n1141 G.n1140 0.624
R10549 G.n1053 G.n1052 0.624
R10550 G.n968 G.n967 0.624
R10551 G.n886 G.n885 0.624
R10552 G.n810 G.n809 0.624
R10553 G.n737 G.n736 0.624
R10554 G.n667 G.n666 0.624
R10555 G.n600 G.n599 0.624
R10556 G.n536 G.n535 0.624
R10557 G.n475 G.n474 0.624
R10558 G.n417 G.n416 0.624
R10559 G.n362 G.n361 0.624
R10560 G.n313 G.n312 0.624
R10561 G.n267 G.n266 0.624
R10562 G.n224 G.n223 0.624
R10563 G.n184 G.n183 0.624
R10564 G.n1741 G.n1740 0.624
R10565 G.n1813 G.n1812 0.624
R10566 G.n1943 G.n1942 0.624
R10567 G.n2000 G.n1999 0.624
R10568 G.n2096 G.n2095 0.624
R10569 G.n2137 G.n2136 0.624
R10570 G.n2048 G.n2047 0.624
R10571 G.n1878 G.n1877 0.624
R10572 G.n1660 G.n1659 0.624
R10573 G.n1490 G.n1489 0.624
R10574 G.n1402 G.n1401 0.624
R10575 G.n1314 G.n1313 0.624
R10576 G.n1226 G.n1225 0.624
R10577 G.n1138 G.n1137 0.624
R10578 G.n1050 G.n1049 0.624
R10579 G.n965 G.n964 0.624
R10580 G.n883 G.n882 0.624
R10581 G.n807 G.n806 0.624
R10582 G.n734 G.n733 0.624
R10583 G.n664 G.n663 0.624
R10584 G.n597 G.n596 0.624
R10585 G.n533 G.n532 0.624
R10586 G.n472 G.n471 0.624
R10587 G.n414 G.n413 0.624
R10588 G.n359 G.n358 0.624
R10589 G.n310 G.n309 0.624
R10590 G.n264 G.n263 0.624
R10591 G.n221 G.n220 0.624
R10592 G.n1577 G.n1576 0.624
R10593 G.n1738 G.n1737 0.624
R10594 G.n1810 G.n1809 0.624
R10595 G.n1940 G.n1939 0.624
R10596 G.n1997 G.n1996 0.624
R10597 G.n2093 G.n2092 0.624
R10598 G.n2134 G.n2133 0.624
R10599 G.n2045 G.n2044 0.624
R10600 G.n1875 G.n1874 0.624
R10601 G.n1657 G.n1656 0.624
R10602 G.n1399 G.n1398 0.624
R10603 G.n1311 G.n1310 0.624
R10604 G.n1223 G.n1222 0.624
R10605 G.n1135 G.n1134 0.624
R10606 G.n1047 G.n1046 0.624
R10607 G.n962 G.n961 0.624
R10608 G.n880 G.n879 0.624
R10609 G.n804 G.n803 0.624
R10610 G.n731 G.n730 0.624
R10611 G.n661 G.n660 0.624
R10612 G.n594 G.n593 0.624
R10613 G.n530 G.n529 0.624
R10614 G.n469 G.n468 0.624
R10615 G.n411 G.n410 0.624
R10616 G.n356 G.n355 0.624
R10617 G.n307 G.n306 0.624
R10618 G.n261 G.n260 0.624
R10619 G.n1487 G.n1486 0.624
R10620 G.n1574 G.n1573 0.624
R10621 G.n1735 G.n1734 0.624
R10622 G.n1807 G.n1806 0.624
R10623 G.n1937 G.n1936 0.624
R10624 G.n1994 G.n1993 0.624
R10625 G.n2090 G.n2089 0.624
R10626 G.n2132 G.n2131 0.624
R10627 G.n2042 G.n2041 0.624
R10628 G.n1872 G.n1871 0.624
R10629 G.n1654 G.n1653 0.624
R10630 G.n1396 G.n1395 0.624
R10631 G.n1220 G.n1219 0.624
R10632 G.n1132 G.n1131 0.624
R10633 G.n1044 G.n1043 0.624
R10634 G.n959 G.n958 0.624
R10635 G.n877 G.n876 0.624
R10636 G.n801 G.n800 0.624
R10637 G.n728 G.n727 0.624
R10638 G.n658 G.n657 0.624
R10639 G.n591 G.n590 0.624
R10640 G.n527 G.n526 0.624
R10641 G.n466 G.n465 0.624
R10642 G.n408 G.n407 0.624
R10643 G.n353 G.n352 0.624
R10644 G.n304 G.n303 0.624
R10645 G.n1308 G.n1307 0.624
R10646 G.n1484 G.n1483 0.624
R10647 G.n1571 G.n1570 0.624
R10648 G.n1732 G.n1731 0.624
R10649 G.n1804 G.n1803 0.624
R10650 G.n1934 G.n1933 0.624
R10651 G.n1991 G.n1990 0.624
R10652 G.n2087 G.n2086 0.624
R10653 G.n2039 G.n2038 0.624
R10654 G.n1869 G.n1868 0.624
R10655 G.n1651 G.n1650 0.624
R10656 G.n1393 G.n1392 0.624
R10657 G.n1129 G.n1128 0.624
R10658 G.n1041 G.n1040 0.624
R10659 G.n956 G.n955 0.624
R10660 G.n874 G.n873 0.624
R10661 G.n798 G.n797 0.624
R10662 G.n725 G.n724 0.624
R10663 G.n655 G.n654 0.624
R10664 G.n588 G.n587 0.624
R10665 G.n524 G.n523 0.624
R10666 G.n463 G.n462 0.624
R10667 G.n405 G.n404 0.624
R10668 G.n350 G.n349 0.624
R10669 G.n1217 G.n1216 0.624
R10670 G.n1305 G.n1304 0.624
R10671 G.n1481 G.n1480 0.624
R10672 G.n1568 G.n1567 0.624
R10673 G.n1729 G.n1728 0.624
R10674 G.n1801 G.n1800 0.624
R10675 G.n1931 G.n1930 0.624
R10676 G.n1988 G.n1987 0.624
R10677 G.n2036 G.n2035 0.624
R10678 G.n1866 G.n1865 0.624
R10679 G.n1648 G.n1647 0.624
R10680 G.n1390 G.n1389 0.624
R10681 G.n1126 G.n1125 0.624
R10682 G.n953 G.n952 0.624
R10683 G.n871 G.n870 0.624
R10684 G.n795 G.n794 0.624
R10685 G.n722 G.n721 0.624
R10686 G.n652 G.n651 0.624
R10687 G.n585 G.n584 0.624
R10688 G.n521 G.n520 0.624
R10689 G.n460 G.n459 0.624
R10690 G.n402 G.n401 0.624
R10691 G.n1038 G.n1037 0.624
R10692 G.n1214 G.n1213 0.624
R10693 G.n1302 G.n1301 0.624
R10694 G.n1478 G.n1477 0.624
R10695 G.n1565 G.n1564 0.624
R10696 G.n1726 G.n1725 0.624
R10697 G.n1798 G.n1797 0.624
R10698 G.n1928 G.n1927 0.624
R10699 G.n1985 G.n1984 0.624
R10700 G.n1863 G.n1862 0.624
R10701 G.n1645 G.n1644 0.624
R10702 G.n1387 G.n1386 0.624
R10703 G.n1123 G.n1122 0.624
R10704 G.n868 G.n867 0.624
R10705 G.n792 G.n791 0.624
R10706 G.n719 G.n718 0.624
R10707 G.n649 G.n648 0.624
R10708 G.n582 G.n581 0.624
R10709 G.n518 G.n517 0.624
R10710 G.n457 G.n456 0.624
R10711 G.n399 G.n398 0.624
R10712 G.n950 G.n949 0.624
R10713 G.n1035 G.n1034 0.624
R10714 G.n1211 G.n1210 0.624
R10715 G.n1299 G.n1298 0.624
R10716 G.n1475 G.n1474 0.624
R10717 G.n1562 G.n1561 0.624
R10718 G.n1723 G.n1722 0.624
R10719 G.n1795 G.n1794 0.624
R10720 G.n1925 G.n1924 0.624
R10721 G.n1982 G.n1981 0.624
R10722 G.n1860 G.n1859 0.624
R10723 G.n1642 G.n1641 0.624
R10724 G.n1384 G.n1383 0.624
R10725 G.n1120 G.n1119 0.624
R10726 G.n865 G.n864 0.624
R10727 G.n716 G.n715 0.624
R10728 G.n646 G.n645 0.624
R10729 G.n579 G.n578 0.624
R10730 G.n515 G.n514 0.624
R10731 G.n454 G.n453 0.624
R10732 G.n789 G.n788 0.624
R10733 G.n947 G.n946 0.624
R10734 G.n1032 G.n1031 0.624
R10735 G.n1208 G.n1207 0.624
R10736 G.n1296 G.n1295 0.624
R10737 G.n1472 G.n1471 0.624
R10738 G.n1559 G.n1558 0.624
R10739 G.n1720 G.n1719 0.624
R10740 G.n1792 G.n1791 0.624
R10741 G.n1922 G.n1921 0.624
R10742 G.n1979 G.n1978 0.624
R10743 G.n1857 G.n1856 0.624
R10744 G.n1639 G.n1638 0.624
R10745 G.n1381 G.n1380 0.624
R10746 G.n1117 G.n1116 0.624
R10747 G.n862 G.n861 0.624
R10748 G.n643 G.n642 0.624
R10749 G.n576 G.n575 0.624
R10750 G.n512 G.n511 0.624
R10751 G.n713 G.n712 0.624
R10752 G.n786 G.n785 0.624
R10753 G.n944 G.n943 0.624
R10754 G.n1029 G.n1028 0.624
R10755 G.n1205 G.n1204 0.624
R10756 G.n1293 G.n1292 0.624
R10757 G.n1469 G.n1468 0.624
R10758 G.n1556 G.n1555 0.624
R10759 G.n1717 G.n1716 0.624
R10760 G.n1789 G.n1788 0.624
R10761 G.n1919 G.n1918 0.624
R10762 G.n1854 G.n1853 0.624
R10763 G.n1636 G.n1635 0.624
R10764 G.n1378 G.n1377 0.624
R10765 G.n1114 G.n1113 0.624
R10766 G.n859 G.n858 0.624
R10767 G.n640 G.n639 0.624
R10768 G.n573 G.n572 0.624
R10769 G.n710 G.n709 0.624
R10770 G.n783 G.n782 0.624
R10771 G.n941 G.n940 0.624
R10772 G.n1026 G.n1025 0.624
R10773 G.n1202 G.n1201 0.624
R10774 G.n1290 G.n1289 0.624
R10775 G.n1466 G.n1465 0.624
R10776 G.n1553 G.n1552 0.624
R10777 G.n1714 G.n1713 0.624
R10778 G.n1786 G.n1785 0.624
R10779 G.n1917 G.n1916 0.624
R10780 G.n1851 G.n1850 0.624
R10781 G.n1633 G.n1632 0.624
R10782 G.n1375 G.n1374 0.624
R10783 G.n1111 G.n1110 0.624
R10784 G.n856 G.n855 0.624
R10785 G.n637 G.n636 0.624
R10786 G.n707 G.n706 0.624
R10787 G.n780 G.n779 0.624
R10788 G.n938 G.n937 0.624
R10789 G.n1023 G.n1022 0.624
R10790 G.n1199 G.n1198 0.624
R10791 G.n1287 G.n1286 0.624
R10792 G.n1463 G.n1462 0.624
R10793 G.n1550 G.n1549 0.624
R10794 G.n1711 G.n1710 0.624
R10795 G.n1783 G.n1782 0.624
R10796 G.n1849 G.n1848 0.624
R10797 G.n1630 G.n1629 0.624
R10798 G.n1372 G.n1371 0.624
R10799 G.n1108 G.n1107 0.624
R10800 G.n853 G.n852 0.624
R10801 G.n704 G.n703 0.624
R10802 G.n777 G.n776 0.624
R10803 G.n935 G.n934 0.624
R10804 G.n1020 G.n1019 0.624
R10805 G.n1196 G.n1195 0.624
R10806 G.n1284 G.n1283 0.624
R10807 G.n1460 G.n1459 0.624
R10808 G.n1547 G.n1546 0.624
R10809 G.n1708 G.n1707 0.624
R10810 G.n1780 G.n1779 0.624
R10811 G.n1627 G.n1626 0.624
R10812 G.n1369 G.n1368 0.624
R10813 G.n1105 G.n1104 0.624
R10814 G.n850 G.n849 0.624
R10815 G.n774 G.n773 0.624
R10816 G.n932 G.n931 0.624
R10817 G.n1017 G.n1016 0.624
R10818 G.n1193 G.n1192 0.624
R10819 G.n1281 G.n1280 0.624
R10820 G.n1457 G.n1456 0.624
R10821 G.n1544 G.n1543 0.624
R10822 G.n1705 G.n1704 0.624
R10823 G.n1777 G.n1776 0.624
R10824 G.n1624 G.n1623 0.624
R10825 G.n1366 G.n1365 0.624
R10826 G.n1102 G.n1101 0.624
R10827 G.n847 G.n846 0.624
R10828 G.n929 G.n928 0.624
R10829 G.n1014 G.n1013 0.624
R10830 G.n1190 G.n1189 0.624
R10831 G.n1278 G.n1277 0.624
R10832 G.n1454 G.n1453 0.624
R10833 G.n1541 G.n1540 0.624
R10834 G.n1702 G.n1701 0.624
R10835 G.n1621 G.n1620 0.624
R10836 G.n1363 G.n1362 0.624
R10837 G.n1099 G.n1098 0.624
R10838 G.n926 G.n925 0.624
R10839 G.n1011 G.n1010 0.624
R10840 G.n1187 G.n1186 0.624
R10841 G.n1275 G.n1274 0.624
R10842 G.n1451 G.n1450 0.624
R10843 G.n1538 G.n1537 0.624
R10844 G.n1699 G.n1698 0.624
R10845 G.n1618 G.n1617 0.624
R10846 G.n1360 G.n1359 0.624
R10847 G.n1096 G.n1095 0.624
R10848 G.n923 G.n922 0.624
R10849 G.n1008 G.n1007 0.624
R10850 G.n1184 G.n1183 0.624
R10851 G.n1272 G.n1271 0.624
R10852 G.n1448 G.n1447 0.624
R10853 G.n1535 G.n1534 0.624
R10854 G.n1616 G.n1615 0.624
R10855 G.n1357 G.n1356 0.624
R10856 G.n1093 G.n1092 0.624
R10857 G.n1005 G.n1004 0.624
R10858 G.n1181 G.n1180 0.624
R10859 G.n1269 G.n1268 0.624
R10860 G.n1445 G.n1444 0.624
R10861 G.n1532 G.n1531 0.624
R10862 G.n1354 G.n1353 0.624
R10863 G.n1090 G.n1089 0.624
R10864 G.n1178 G.n1177 0.624
R10865 G.n1266 G.n1265 0.624
R10866 G.n1442 G.n1441 0.624
R10867 G.n1529 G.n1528 0.624
R10868 G.n6408 G.n6407 0.624
R10869 G.n6250 G.n6248 0.624
R10870 G.n6088 G.n6086 0.624
R10871 G.n6142 G.n6140 0.624
R10872 G.n6196 G.n6194 0.624
R10873 G.n6304 G.n6302 0.624
R10874 G.n6357 G.n6355 0.624
R10875 G.n6410 G.n6409 0.624
R10876 G.n6252 G.n6251 0.624
R10877 G.n6090 G.n6089 0.624
R10878 G.n6038 G.n6037 0.624
R10879 G.n5987 G.n5986 0.624
R10880 G.n6144 G.n6143 0.624
R10881 G.n6198 G.n6197 0.624
R10882 G.n6306 G.n6305 0.624
R10883 G.n6359 G.n6358 0.624
R10884 G.n6458 G.n6457 0.624
R10885 G.n6413 G.n6411 0.624
R10886 G.n6255 G.n6253 0.624
R10887 G.n6093 G.n6091 0.624
R10888 G.n6041 G.n6039 0.624
R10889 G.n5990 G.n5988 0.624
R10890 G.n5941 G.n5939 0.624
R10891 G.n6147 G.n6145 0.624
R10892 G.n6201 G.n6199 0.624
R10893 G.n6309 G.n6307 0.624
R10894 G.n6362 G.n6360 0.624
R10895 G.n6461 G.n6459 0.624
R10896 G.n6415 G.n6414 0.624
R10897 G.n6257 G.n6256 0.624
R10898 G.n6203 G.n6202 0.624
R10899 G.n6149 G.n6148 0.624
R10900 G.n6095 G.n6094 0.624
R10901 G.n6043 G.n6042 0.624
R10902 G.n5992 G.n5991 0.624
R10903 G.n5943 G.n5942 0.624
R10904 G.n5897 G.n5896 0.624
R10905 G.n5852 G.n5851 0.624
R10906 G.n6311 G.n6310 0.624
R10907 G.n6364 G.n6363 0.624
R10908 G.n6463 G.n6462 0.624
R10909 G.n6507 G.n6506 0.624
R10910 G.n6551 G.n6549 0.624
R10911 G.n6418 G.n6416 0.624
R10912 G.n6260 G.n6258 0.624
R10913 G.n6206 G.n6204 0.624
R10914 G.n6152 G.n6150 0.624
R10915 G.n6098 G.n6096 0.624
R10916 G.n6046 G.n6044 0.624
R10917 G.n5995 G.n5993 0.624
R10918 G.n5946 G.n5944 0.624
R10919 G.n5900 G.n5898 0.624
R10920 G.n5855 G.n5853 0.624
R10921 G.n5812 G.n5810 0.624
R10922 G.n6314 G.n6312 0.624
R10923 G.n6367 G.n6365 0.624
R10924 G.n6466 G.n6464 0.624
R10925 G.n6510 G.n6508 0.624
R10926 G.n6553 G.n6552 0.624
R10927 G.n6420 G.n6419 0.624
R10928 G.n6369 G.n6368 0.624
R10929 G.n6316 G.n6315 0.624
R10930 G.n6262 G.n6261 0.624
R10931 G.n6208 G.n6207 0.624
R10932 G.n6154 G.n6153 0.624
R10933 G.n6100 G.n6099 0.624
R10934 G.n6048 G.n6047 0.624
R10935 G.n5997 G.n5996 0.624
R10936 G.n5948 G.n5947 0.624
R10937 G.n5902 G.n5901 0.624
R10938 G.n5857 G.n5856 0.624
R10939 G.n5814 G.n5813 0.624
R10940 G.n5774 G.n5773 0.624
R10941 G.n5735 G.n5734 0.624
R10942 G.n6468 G.n6467 0.624
R10943 G.n6512 G.n6511 0.624
R10944 G.n6590 G.n6589 0.624
R10945 G.n6556 G.n6554 0.624
R10946 G.n6423 G.n6421 0.624
R10947 G.n6372 G.n6370 0.624
R10948 G.n6319 G.n6317 0.624
R10949 G.n6265 G.n6263 0.624
R10950 G.n6211 G.n6209 0.624
R10951 G.n6157 G.n6155 0.624
R10952 G.n6103 G.n6101 0.624
R10953 G.n6051 G.n6049 0.624
R10954 G.n6000 G.n5998 0.624
R10955 G.n5951 G.n5949 0.624
R10956 G.n5905 G.n5903 0.624
R10957 G.n5860 G.n5858 0.624
R10958 G.n5817 G.n5815 0.624
R10959 G.n5777 G.n5775 0.624
R10960 G.n5738 G.n5736 0.624
R10961 G.n5701 G.n5699 0.624
R10962 G.n6471 G.n6469 0.624
R10963 G.n6515 G.n6513 0.624
R10964 G.n6593 G.n6591 0.624
R10965 G.n6626 G.n6625 0.624
R10966 G.n6658 G.n6657 0.624
R10967 G.n6558 G.n6557 0.624
R10968 G.n6517 G.n6516 0.624
R10969 G.n6473 G.n6472 0.624
R10970 G.n6425 G.n6424 0.624
R10971 G.n6374 G.n6373 0.624
R10972 G.n6321 G.n6320 0.624
R10973 G.n6267 G.n6266 0.624
R10974 G.n6213 G.n6212 0.624
R10975 G.n6159 G.n6158 0.624
R10976 G.n6105 G.n6104 0.624
R10977 G.n6053 G.n6052 0.624
R10978 G.n6002 G.n6001 0.624
R10979 G.n5953 G.n5952 0.624
R10980 G.n5907 G.n5906 0.624
R10981 G.n5862 G.n5861 0.624
R10982 G.n5819 G.n5818 0.624
R10983 G.n5779 G.n5778 0.624
R10984 G.n5740 G.n5739 0.624
R10985 G.n5703 G.n5702 0.624
R10986 G.n5669 G.n5668 0.624
R10987 G.n5638 G.n5637 0.624
R10988 G.n6595 G.n6594 0.624
R10989 G.n6628 G.n6627 0.624
R10990 G.n6661 G.n6659 0.624
R10991 G.n6561 G.n6559 0.624
R10992 G.n6520 G.n6518 0.624
R10993 G.n6476 G.n6474 0.624
R10994 G.n6428 G.n6426 0.624
R10995 G.n6377 G.n6375 0.624
R10996 G.n6324 G.n6322 0.624
R10997 G.n6270 G.n6268 0.624
R10998 G.n6216 G.n6214 0.624
R10999 G.n6162 G.n6160 0.624
R11000 G.n6108 G.n6106 0.624
R11001 G.n6056 G.n6054 0.624
R11002 G.n6005 G.n6003 0.624
R11003 G.n5956 G.n5954 0.624
R11004 G.n5910 G.n5908 0.624
R11005 G.n5865 G.n5863 0.624
R11006 G.n5822 G.n5820 0.624
R11007 G.n5782 G.n5780 0.624
R11008 G.n5743 G.n5741 0.624
R11009 G.n5706 G.n5704 0.624
R11010 G.n5672 G.n5670 0.624
R11011 G.n5641 G.n5639 0.624
R11012 G.n5610 G.n5608 0.624
R11013 G.n6598 G.n6596 0.624
R11014 G.n6631 G.n6629 0.624
R11015 G.n6688 G.n6687 0.624
R11016 G.n6663 G.n6662 0.624
R11017 G.n6633 G.n6632 0.624
R11018 G.n6600 G.n6599 0.624
R11019 G.n6563 G.n6562 0.624
R11020 G.n6522 G.n6521 0.624
R11021 G.n6478 G.n6477 0.624
R11022 G.n6430 G.n6429 0.624
R11023 G.n6379 G.n6378 0.624
R11024 G.n6326 G.n6325 0.624
R11025 G.n6272 G.n6271 0.624
R11026 G.n6218 G.n6217 0.624
R11027 G.n6164 G.n6163 0.624
R11028 G.n6110 G.n6109 0.624
R11029 G.n6058 G.n6057 0.624
R11030 G.n6007 G.n6006 0.624
R11031 G.n5958 G.n5957 0.624
R11032 G.n5912 G.n5911 0.624
R11033 G.n5867 G.n5866 0.624
R11034 G.n5824 G.n5823 0.624
R11035 G.n5784 G.n5783 0.624
R11036 G.n5745 G.n5744 0.624
R11037 G.n5708 G.n5707 0.624
R11038 G.n5674 G.n5673 0.624
R11039 G.n5643 G.n5642 0.624
R11040 G.n5612 G.n5611 0.624
R11041 G.n5584 G.n5583 0.624
R11042 G.n5559 G.n5558 0.624
R11043 G.n6690 G.n6689 0.624
R11044 G.n6714 G.n6713 0.624
R11045 G.n6738 G.n6737 0.624
R11046 G.n6666 G.n6664 0.624
R11047 G.n6636 G.n6634 0.624
R11048 G.n6603 G.n6601 0.624
R11049 G.n6566 G.n6564 0.624
R11050 G.n6525 G.n6523 0.624
R11051 G.n6481 G.n6479 0.624
R11052 G.n6433 G.n6431 0.624
R11053 G.n6382 G.n6380 0.624
R11054 G.n6329 G.n6327 0.624
R11055 G.n6275 G.n6273 0.624
R11056 G.n6221 G.n6219 0.624
R11057 G.n6167 G.n6165 0.624
R11058 G.n6113 G.n6111 0.624
R11059 G.n6061 G.n6059 0.624
R11060 G.n6010 G.n6008 0.624
R11061 G.n5961 G.n5959 0.624
R11062 G.n5915 G.n5913 0.624
R11063 G.n5870 G.n5868 0.624
R11064 G.n5827 G.n5825 0.624
R11065 G.n5787 G.n5785 0.624
R11066 G.n5748 G.n5746 0.624
R11067 G.n5711 G.n5709 0.624
R11068 G.n5677 G.n5675 0.624
R11069 G.n5646 G.n5644 0.624
R11070 G.n5615 G.n5613 0.624
R11071 G.n5587 G.n5585 0.624
R11072 G.n5562 G.n5560 0.624
R11073 G.n5537 G.n5535 0.624
R11074 G.n6693 G.n6691 0.624
R11075 G.n6717 G.n6715 0.624
R11076 G.n6740 G.n6739 0.624
R11077 G.n6719 G.n6718 0.624
R11078 G.n6695 G.n6694 0.624
R11079 G.n6668 G.n6667 0.624
R11080 G.n6638 G.n6637 0.624
R11081 G.n6605 G.n6604 0.624
R11082 G.n6568 G.n6567 0.624
R11083 G.n6527 G.n6526 0.624
R11084 G.n6483 G.n6482 0.624
R11085 G.n6435 G.n6434 0.624
R11086 G.n6384 G.n6383 0.624
R11087 G.n6331 G.n6330 0.624
R11088 G.n6277 G.n6276 0.624
R11089 G.n6223 G.n6222 0.624
R11090 G.n6169 G.n6168 0.624
R11091 G.n6115 G.n6114 0.624
R11092 G.n6063 G.n6062 0.624
R11093 G.n6012 G.n6011 0.624
R11094 G.n5963 G.n5962 0.624
R11095 G.n5917 G.n5916 0.624
R11096 G.n5872 G.n5871 0.624
R11097 G.n5829 G.n5828 0.624
R11098 G.n5789 G.n5788 0.624
R11099 G.n5750 G.n5749 0.624
R11100 G.n5713 G.n5712 0.624
R11101 G.n5679 G.n5678 0.624
R11102 G.n5648 G.n5647 0.624
R11103 G.n5617 G.n5616 0.624
R11104 G.n5589 G.n5588 0.624
R11105 G.n5564 G.n5563 0.624
R11106 G.n5539 G.n5538 0.624
R11107 G.n5517 G.n5516 0.624
R11108 G.n6758 G.n6757 0.624
R11109 G.n6743 G.n6741 0.624
R11110 G.n6722 G.n6720 0.624
R11111 G.n6698 G.n6696 0.624
R11112 G.n6671 G.n6669 0.624
R11113 G.n6641 G.n6639 0.624
R11114 G.n6608 G.n6606 0.624
R11115 G.n6571 G.n6569 0.624
R11116 G.n6530 G.n6528 0.624
R11117 G.n6486 G.n6484 0.624
R11118 G.n6438 G.n6436 0.624
R11119 G.n6387 G.n6385 0.624
R11120 G.n6334 G.n6332 0.624
R11121 G.n6280 G.n6278 0.624
R11122 G.n6226 G.n6224 0.624
R11123 G.n6172 G.n6170 0.624
R11124 G.n6118 G.n6116 0.624
R11125 G.n6066 G.n6064 0.624
R11126 G.n6015 G.n6013 0.624
R11127 G.n5966 G.n5964 0.624
R11128 G.n5920 G.n5918 0.624
R11129 G.n5875 G.n5873 0.624
R11130 G.n5832 G.n5830 0.624
R11131 G.n5792 G.n5790 0.624
R11132 G.n5753 G.n5751 0.624
R11133 G.n5716 G.n5714 0.624
R11134 G.n5682 G.n5680 0.624
R11135 G.n5651 G.n5649 0.624
R11136 G.n5620 G.n5618 0.624
R11137 G.n5592 G.n5590 0.624
R11138 G.n5567 G.n5565 0.624
R11139 G.n5542 G.n5540 0.624
R11140 G.n5520 G.n5518 0.624
R11141 G.n5501 G.n5499 0.624
R11142 G.n5483 G.n5481 0.624
R11143 G.n6761 G.n6759 0.624
R11144 G.n6776 G.n6775 0.624
R11145 G.n3455 G.n3451 0.624
R11146 G.n3457 G.n3450 0.624
R11147 G.n6790 G.n6789 0.624
R11148 G.n6789 G.n6788 0.624
R11149 G.n6779 G.n6778 0.624
R11150 G.n6778 G.n6777 0.624
R11151 G.n6764 G.n6763 0.624
R11152 G.n6763 G.n6762 0.624
R11153 G.n6746 G.n6745 0.624
R11154 G.n6745 G.n6744 0.624
R11155 G.n6725 G.n6724 0.624
R11156 G.n6724 G.n6723 0.624
R11157 G.n6701 G.n6700 0.624
R11158 G.n6700 G.n6699 0.624
R11159 G.n6674 G.n6673 0.624
R11160 G.n6673 G.n6672 0.624
R11161 G.n6644 G.n6643 0.624
R11162 G.n6643 G.n6642 0.624
R11163 G.n6611 G.n6610 0.624
R11164 G.n6610 G.n6609 0.624
R11165 G.n6574 G.n6573 0.624
R11166 G.n6573 G.n6572 0.624
R11167 G.n6533 G.n6532 0.624
R11168 G.n6532 G.n6531 0.624
R11169 G.n6489 G.n6488 0.624
R11170 G.n6488 G.n6487 0.624
R11171 G.n6441 G.n6440 0.624
R11172 G.n6440 G.n6439 0.624
R11173 G.n6390 G.n6389 0.624
R11174 G.n6389 G.n6388 0.624
R11175 G.n6337 G.n6336 0.624
R11176 G.n6336 G.n6335 0.624
R11177 G.n6283 G.n6282 0.624
R11178 G.n6282 G.n6281 0.624
R11179 G.n6229 G.n6228 0.624
R11180 G.n6228 G.n6227 0.624
R11181 G.n6175 G.n6174 0.624
R11182 G.n6174 G.n6173 0.624
R11183 G.n6121 G.n6120 0.624
R11184 G.n6120 G.n6119 0.624
R11185 G.n6069 G.n6068 0.624
R11186 G.n6068 G.n6067 0.624
R11187 G.n6018 G.n6017 0.624
R11188 G.n6017 G.n6016 0.624
R11189 G.n5969 G.n5968 0.624
R11190 G.n5968 G.n5967 0.624
R11191 G.n5923 G.n5922 0.624
R11192 G.n5922 G.n5921 0.624
R11193 G.n5878 G.n5877 0.624
R11194 G.n5877 G.n5876 0.624
R11195 G.n5835 G.n5834 0.624
R11196 G.n5834 G.n5833 0.624
R11197 G.n5795 G.n5794 0.624
R11198 G.n5794 G.n5793 0.624
R11199 G.n5756 G.n5755 0.624
R11200 G.n5755 G.n5754 0.624
R11201 G.n5719 G.n5718 0.624
R11202 G.n5718 G.n5717 0.624
R11203 G.n5685 G.n5684 0.624
R11204 G.n5684 G.n5683 0.624
R11205 G.n5654 G.n5653 0.624
R11206 G.n5653 G.n5652 0.624
R11207 G.n5623 G.n5622 0.624
R11208 G.n5622 G.n5621 0.624
R11209 G.n5595 G.n5594 0.624
R11210 G.n5594 G.n5593 0.624
R11211 G.n5570 G.n5569 0.624
R11212 G.n5569 G.n5568 0.624
R11213 G.n5545 G.n5544 0.624
R11214 G.n5544 G.n5543 0.624
R11215 G.n5523 G.n5522 0.624
R11216 G.n5522 G.n5521 0.624
R11217 G.n5504 G.n5503 0.624
R11218 G.n5503 G.n5502 0.624
R11219 G.n5486 G.n5485 0.624
R11220 G.n5485 G.n5484 0.624
R11221 G.n5470 G.n5469 0.624
R11222 G.n5469 G.n5468 0.624
R11223 G.n5457 G.n5456 0.624
R11224 G.n5393 G.n5392 0.624
R11225 G.n5396 G.n5395 0.624
R11226 G.n5399 G.n5398 0.624
R11227 G.n5402 G.n5401 0.624
R11228 G.n2282 G.n2281 0.624
R11229 G.n2284 G.n2283 0.624
R11230 G.n2296 G.n2295 0.624
R11231 G.n7 G.n6 0.624
R11232 G.n3564 G.n3 0.624
R11233 G.n5428 G.n5426 0.624
R11234 G.n6815 G.n6814 0.624
R11235 G G.n3564 0.339
R11236 G.n6816 G.n6815 0.305
R11237 G.n6817 G.n6816 0.305
R11238 G.n6818 G.n6817 0.305
R11239 G.n6819 G.n6818 0.305
R11240 G.n6820 G.n6819 0.305
R11241 G.n6821 G.n6820 0.305
R11242 G.n6822 G.n6821 0.305
R11243 G.n6823 G.n6822 0.305
R11244 G.n6824 G.n6823 0.305
R11245 G.n6825 G.n6824 0.305
R11246 G.n6826 G.n6825 0.305
R11247 G.n6827 G.n6826 0.305
R11248 G.n6828 G.n6827 0.305
R11249 G.n6829 G.n6828 0.305
R11250 G.n6830 G.n6829 0.305
R11251 G.n6831 G.n6830 0.305
R11252 G.n6832 G.n6831 0.305
R11253 G.n6833 G.n6832 0.305
R11254 G.n6834 G.n6833 0.305
R11255 G.n6835 G.n6834 0.305
R11256 G.n6836 G.n6835 0.305
R11257 G.n6837 G.n6836 0.305
R11258 G.n6838 G.n6837 0.305
R11259 G.n6839 G.n6838 0.305
R11260 G.n6840 G.n6839 0.305
R11261 G.n6841 G.n6840 0.305
R11262 G.n6842 G.n6841 0.305
R11263 G.n6843 G.n6842 0.305
R11264 G.n6844 G.n6843 0.305
R11265 G.n6845 G.n6844 0.305
R11266 G.n6846 G.n6845 0.305
R11267 G.n6847 G.n6846 0.305
R11268 G.n6848 G.n6847 0.305
R11269 G.n6849 G.n6848 0.305
R11270 G.n6850 G.n6849 0.305
R11271 G.n6851 G.n6850 0.305
R11272 G.n6852 G.n6851 0.305
R11273 G.n6853 G.n6852 0.305
R11274 G.n6854 G.n6853 0.305
R11275 G.n6855 G.n6854 0.305
R11276 G.n6856 G.n6855 0.305
R11277 G.n6857 G.n6856 0.305
R11278 G.n6858 G.n6857 0.305
R11279 G.n6859 G.n6858 0.305
R11280 G.n6860 G.n6859 0.305
R11281 G.n6861 G.n6860 0.305
R11282 G.n3519 G.n3518 0.305
R11283 G.n3520 G.n3519 0.305
R11284 G.n3521 G.n3520 0.305
R11285 G.n3522 G.n3521 0.305
R11286 G.n3523 G.n3522 0.305
R11287 G.n3524 G.n3523 0.305
R11288 G.n3525 G.n3524 0.305
R11289 G.n3526 G.n3525 0.305
R11290 G.n3527 G.n3526 0.305
R11291 G.n3528 G.n3527 0.305
R11292 G.n3529 G.n3528 0.305
R11293 G.n3530 G.n3529 0.305
R11294 G.n3531 G.n3530 0.305
R11295 G.n3532 G.n3531 0.305
R11296 G.n3533 G.n3532 0.305
R11297 G.n3534 G.n3533 0.305
R11298 G.n3535 G.n3534 0.305
R11299 G.n3536 G.n3535 0.305
R11300 G.n3537 G.n3536 0.305
R11301 G.n3538 G.n3537 0.305
R11302 G.n3539 G.n3538 0.305
R11303 G.n3540 G.n3539 0.305
R11304 G.n3541 G.n3540 0.305
R11305 G.n3542 G.n3541 0.305
R11306 G.n3543 G.n3542 0.305
R11307 G.n3544 G.n3543 0.305
R11308 G.n3545 G.n3544 0.305
R11309 G.n3546 G.n3545 0.305
R11310 G.n3547 G.n3546 0.305
R11311 G.n3548 G.n3547 0.305
R11312 G.n3549 G.n3548 0.305
R11313 G.n3550 G.n3549 0.305
R11314 G.n3551 G.n3550 0.305
R11315 G.n3552 G.n3551 0.305
R11316 G.n3553 G.n3552 0.305
R11317 G.n3554 G.n3553 0.305
R11318 G.n3555 G.n3554 0.305
R11319 G.n3556 G.n3555 0.305
R11320 G.n3557 G.n3556 0.305
R11321 G.n3558 G.n3557 0.305
R11322 G.n3559 G.n3558 0.305
R11323 G.n3560 G.n3559 0.305
R11324 G.n3561 G.n3560 0.305
R11325 G.n3562 G.n3561 0.305
R11326 G.n3563 G.n3562 0.305
R11327 G.n3564 G.n3563 0.305
R11328 G.n3472 G.n3471 0.305
R11329 G.n3473 G.n3472 0.305
R11330 G.n3474 G.n3473 0.305
R11331 G.n3475 G.n3474 0.305
R11332 G.n3476 G.n3475 0.305
R11333 G.n3477 G.n3476 0.305
R11334 G.n3478 G.n3477 0.305
R11335 G.n3479 G.n3478 0.305
R11336 G.n3480 G.n3479 0.305
R11337 G.n3481 G.n3480 0.305
R11338 G.n3482 G.n3481 0.305
R11339 G.n3483 G.n3482 0.305
R11340 G.n3484 G.n3483 0.305
R11341 G.n3485 G.n3484 0.305
R11342 G.n3486 G.n3485 0.305
R11343 G.n3487 G.n3486 0.305
R11344 G.n3488 G.n3487 0.305
R11345 G.n3489 G.n3488 0.305
R11346 G.n3490 G.n3489 0.305
R11347 G.n3491 G.n3490 0.305
R11348 G.n3492 G.n3491 0.305
R11349 G.n3493 G.n3492 0.305
R11350 G.n3494 G.n3493 0.305
R11351 G.n3495 G.n3494 0.305
R11352 G.n3496 G.n3495 0.305
R11353 G.n3497 G.n3496 0.305
R11354 G.n3498 G.n3497 0.305
R11355 G.n3499 G.n3498 0.305
R11356 G.n3500 G.n3499 0.305
R11357 G.n3501 G.n3500 0.305
R11358 G.n3502 G.n3501 0.305
R11359 G.n3503 G.n3502 0.305
R11360 G.n3504 G.n3503 0.305
R11361 G.n3505 G.n3504 0.305
R11362 G.n3506 G.n3505 0.305
R11363 G.n3507 G.n3506 0.305
R11364 G.n3508 G.n3507 0.305
R11365 G.n3509 G.n3508 0.305
R11366 G.n3510 G.n3509 0.305
R11367 G.n3511 G.n3510 0.305
R11368 G.n3512 G.n3511 0.305
R11369 G.n3513 G.n3512 0.305
R11370 G.n3514 G.n3513 0.305
R11371 G.n3515 G.n3514 0.305
R11372 G.n3516 G.n3515 0.305
R11373 G.n3517 G.n3516 0.305
R11374 G.n6863 G.n6862 0.305
R11375 G.n6864 G.n6863 0.305
R11376 G.n6865 G.n6864 0.305
R11377 G.n6866 G.n6865 0.305
R11378 G.n6867 G.n6866 0.305
R11379 G.n6868 G.n6867 0.305
R11380 G.n6869 G.n6868 0.305
R11381 G.n6870 G.n6869 0.305
R11382 G.n6871 G.n6870 0.305
R11383 G.n6872 G.n6871 0.305
R11384 G.n6873 G.n6872 0.305
R11385 G.n6874 G.n6873 0.305
R11386 G.n6875 G.n6874 0.305
R11387 G.n6876 G.n6875 0.305
R11388 G.n6877 G.n6876 0.305
R11389 G.n6878 G.n6877 0.305
R11390 G.n6879 G.n6878 0.305
R11391 G.n6880 G.n6879 0.305
R11392 G.n6881 G.n6880 0.305
R11393 G.n6882 G.n6881 0.305
R11394 G.n6883 G.n6882 0.305
R11395 G.n6884 G.n6883 0.305
R11396 G.n6885 G.n6884 0.305
R11397 G.n6886 G.n6885 0.305
R11398 G.n6887 G.n6886 0.305
R11399 G.n6888 G.n6887 0.305
R11400 G.n6889 G.n6888 0.305
R11401 G.n6890 G.n6889 0.305
R11402 G.n6891 G.n6890 0.305
R11403 G.n6892 G.n6891 0.305
R11404 G.n6893 G.n6892 0.305
R11405 G.n6894 G.n6893 0.305
R11406 G.n6895 G.n6894 0.305
R11407 G.n6896 G.n6895 0.305
R11408 G.n6897 G.n6896 0.305
R11409 G.n6898 G.n6897 0.305
R11410 G.n6899 G.n6898 0.305
R11411 G.n6900 G.n6899 0.305
R11412 G.n6901 G.n6900 0.305
R11413 G.n6902 G.n6901 0.305
R11414 G.n6903 G.n6902 0.305
R11415 G.n6904 G.n6903 0.305
R11416 G.n6905 G.n6904 0.305
R11417 G.n6906 G.n6905 0.305
R11418 G.n6907 G.n6906 0.305
R11419 G.n6908 G.n6907 0.305
R11420 G G.n6908 0.305
R11421 D.n7835 D.t282 7.599
R11422 D.n7825 D.t2794 7.599
R11423 D.n447 D.t3021 7.599
R11424 D.n438 D.t792 7.599
R11425 D.n28 D.t4247 7.599
R11426 D.n7930 D.t440 7.599
R11427 D.n7955 D.t358 7.599
R11428 D.n7940 D.t1940 7.599
R11429 D.n14061 D.t606 7.599
R11430 D.n14043 D.t905 7.599
R11431 D.n14025 D.t2054 7.599
R11432 D.n14007 D.t3812 7.599
R11433 D.n13989 D.t4380 7.599
R11434 D.n13971 D.t3634 7.599
R11435 D.n13953 D.t3584 7.599
R11436 D.n13935 D.t4100 7.599
R11437 D.n13917 D.t4155 7.599
R11438 D.n13899 D.t4169 7.599
R11439 D.n13881 D.t3296 7.599
R11440 D.n13863 D.t475 7.599
R11441 D.n13845 D.t1573 7.599
R11442 D.n13827 D.t2856 7.599
R11443 D.n13809 D.t1039 7.599
R11444 D.n13791 D.t1015 7.599
R11445 D.n13773 D.t1067 7.599
R11446 D.n13755 D.t728 7.599
R11447 D.n13737 D.t2099 7.599
R11448 D.n13719 D.t3558 7.599
R11449 D.n13701 D.t3106 7.599
R11450 D.n13682 D.t380 7.599
R11451 D.n13691 D.t3795 7.599
R11452 D.n13709 D.t130 7.599
R11453 D.n13727 D.t4381 7.599
R11454 D.n13745 D.t3306 7.599
R11455 D.n13763 D.t2190 7.599
R11456 D.n13781 D.t1358 7.599
R11457 D.n13799 D.t1862 7.599
R11458 D.n13817 D.t271 7.599
R11459 D.n13835 D.t1336 7.599
R11460 D.n13853 D.t2829 7.599
R11461 D.n13871 D.t851 7.599
R11462 D.n13889 D.t1135 7.599
R11463 D.n13907 D.t4477 7.599
R11464 D.n13925 D.t4396 7.599
R11465 D.n13943 D.t1893 7.599
R11466 D.n13961 D.t2488 7.599
R11467 D.n13979 D.t1832 7.599
R11468 D.n13997 D.t744 7.599
R11469 D.n14015 D.t3461 7.599
R11470 D.n14033 D.t3721 7.599
R11471 D.n14051 D.t3556 7.599
R11472 D.n14073 D.t428 7.599
R11473 D.n14090 D.t1999 7.599
R11474 D.n13207 D.t118 7.599
R11475 D.n13227 D.t947 7.599
R11476 D.n13247 D.t3630 7.599
R11477 D.n13267 D.t1811 7.599
R11478 D.n13287 D.t1774 7.599
R11479 D.n13307 D.t3426 7.599
R11480 D.n13327 D.t3935 7.599
R11481 D.n13347 D.t3684 7.599
R11482 D.n13367 D.t3378 7.599
R11483 D.n13387 D.t842 7.599
R11484 D.n13407 D.t4442 7.599
R11485 D.n13427 D.t3198 7.599
R11486 D.n13447 D.t529 7.599
R11487 D.n13467 D.t4053 7.599
R11488 D.n13487 D.t4143 7.599
R11489 D.n13507 D.t154 7.599
R11490 D.n13527 D.t303 7.599
R11491 D.n13547 D.t1248 7.599
R11492 D.n13567 D.t1935 7.599
R11493 D.n13587 D.t2486 7.599
R11494 D.n13607 D.t1795 7.599
R11495 D.n13595 D.t2958 7.599
R11496 D.n13575 D.t2847 7.599
R11497 D.n13555 D.t864 7.599
R11498 D.n13535 D.t1094 7.599
R11499 D.n13515 D.t676 7.599
R11500 D.n13495 D.t893 7.599
R11501 D.n13475 D.t1853 7.599
R11502 D.n13455 D.t4507 7.599
R11503 D.n13435 D.t3934 7.599
R11504 D.n13415 D.t2311 7.599
R11505 D.n13395 D.t246 7.599
R11506 D.n13375 D.t3635 7.599
R11507 D.n13355 D.t1220 7.599
R11508 D.n13335 D.t2294 7.599
R11509 D.n13315 D.t2642 7.599
R11510 D.n13295 D.t365 7.599
R11511 D.n13275 D.t3631 7.599
R11512 D.n13255 D.t95 7.599
R11513 D.n13235 D.t494 7.599
R11514 D.n13215 D.t621 7.599
R11515 D.n13190 D.t2698 7.599
R11516 D.n13177 D.t593 7.599
R11517 D.n13098 D.t1607 7.599
R11518 D.n13080 D.t1780 7.599
R11519 D.n13062 D.t102 7.599
R11520 D.n13044 D.t1172 7.599
R11521 D.n13026 D.t1104 7.599
R11522 D.n13008 D.t521 7.599
R11523 D.n12990 D.t523 7.599
R11524 D.n12972 D.t1861 7.599
R11525 D.n12954 D.t115 7.599
R11526 D.n12936 D.t3628 7.599
R11527 D.n12918 D.t4225 7.599
R11528 D.n12900 D.t1966 7.599
R11529 D.n12882 D.t2639 7.599
R11530 D.n12864 D.t3190 7.599
R11531 D.n12846 D.t3109 7.599
R11532 D.n12828 D.t2559 7.599
R11533 D.n12810 D.t1003 7.599
R11534 D.n12792 D.t1083 7.599
R11535 D.n12774 D.t2985 7.599
R11536 D.n12755 D.t3316 7.599
R11537 D.n12764 D.t1997 7.599
R11538 D.n12782 D.t2323 7.599
R11539 D.n12800 D.t1366 7.599
R11540 D.n12818 D.t1333 7.599
R11541 D.n12836 D.t644 7.599
R11542 D.n12854 D.t2764 7.599
R11543 D.n12872 D.t3912 7.599
R11544 D.n12890 D.t557 7.599
R11545 D.n12908 D.t1808 7.599
R11546 D.n12926 D.t4496 7.599
R11547 D.n12944 D.t4068 7.599
R11548 D.n12962 D.t3726 7.599
R11549 D.n12980 D.t2039 7.599
R11550 D.n12998 D.t1742 7.599
R11551 D.n13016 D.t2692 7.599
R11552 D.n13034 D.t4373 7.599
R11553 D.n13052 D.t4286 7.599
R11554 D.n13070 D.t4201 7.599
R11555 D.n13088 D.t3245 7.599
R11556 D.n13109 D.t1678 7.599
R11557 D.n13120 D.t357 7.599
R11558 D.n12324 D.t4161 7.599
R11559 D.n12344 D.t4089 7.599
R11560 D.n12364 D.t3070 7.599
R11561 D.n12384 D.t3582 7.599
R11562 D.n12404 D.t4213 7.599
R11563 D.n12424 D.t3443 7.599
R11564 D.n12444 D.t4394 7.599
R11565 D.n12464 D.t4300 7.599
R11566 D.n12484 D.t4114 7.599
R11567 D.n12504 D.t1445 7.599
R11568 D.n12524 D.t2955 7.599
R11569 D.n12544 D.t3962 7.599
R11570 D.n12564 D.t3522 7.599
R11571 D.n12584 D.t2448 7.599
R11572 D.n12604 D.t3984 7.599
R11573 D.n12624 D.t3317 7.599
R11574 D.n12644 D.t1544 7.599
R11575 D.n12664 D.t733 7.599
R11576 D.n12684 D.t1772 7.599
R11577 D.n12672 D.t1030 7.599
R11578 D.n12652 D.t659 7.599
R11579 D.n12632 D.t12 7.599
R11580 D.n12612 D.t4108 7.599
R11581 D.n12592 D.t854 7.599
R11582 D.n12572 D.t1221 7.599
R11583 D.n12552 D.t3871 7.599
R11584 D.n12532 D.t1838 7.599
R11585 D.n12512 D.t1991 7.599
R11586 D.n12492 D.t582 7.599
R11587 D.n12472 D.t4287 7.599
R11588 D.n12452 D.t4265 7.599
R11589 D.n12432 D.t2223 7.599
R11590 D.n12412 D.t3160 7.599
R11591 D.n12392 D.t341 7.599
R11592 D.n12372 D.t3543 7.599
R11593 D.n12352 D.t1258 7.599
R11594 D.n12332 D.t2474 7.599
R11595 D.n12307 D.t2788 7.599
R11596 D.n12294 D.t1575 7.599
R11597 D.n12213 D.t3280 7.599
R11598 D.n12195 D.t965 7.599
R11599 D.n12177 D.t200 7.599
R11600 D.n12159 D.t1803 7.599
R11601 D.n12141 D.t657 7.599
R11602 D.n12123 D.t3870 7.599
R11603 D.n12105 D.t3419 7.599
R11604 D.n12087 D.t3390 7.599
R11605 D.n12069 D.t2855 7.599
R11606 D.n12051 D.t2391 7.599
R11607 D.n12033 D.t3813 7.599
R11608 D.n12015 D.t4061 7.599
R11609 D.n11997 D.t2814 7.599
R11610 D.n11979 D.t294 7.599
R11611 D.n11961 D.t620 7.599
R11612 D.n11943 D.t2998 7.599
R11613 D.n11925 D.t794 7.599
R11614 D.n11906 D.t2782 7.599
R11615 D.n11915 D.t3209 7.599
R11616 D.n11933 D.t1214 7.599
R11617 D.n11951 D.t773 7.599
R11618 D.n11969 D.t4218 7.599
R11619 D.n11987 D.t1667 7.599
R11620 D.n12005 D.t2467 7.599
R11621 D.n12023 D.t1281 7.599
R11622 D.n12041 D.t2540 7.599
R11623 D.n12059 D.t2845 7.599
R11624 D.n12077 D.t899 7.599
R11625 D.n12095 D.t3181 7.599
R11626 D.n12113 D.t2508 7.599
R11627 D.n12131 D.t2458 7.599
R11628 D.n12149 D.t1876 7.599
R11629 D.n12167 D.t1646 7.599
R11630 D.n12185 D.t337 7.599
R11631 D.n12203 D.t2111 7.599
R11632 D.n12225 D.t1219 7.599
R11633 D.n12242 D.t420 7.599
R11634 D.n11515 D.t1016 7.599
R11635 D.n11535 D.t1743 7.599
R11636 D.n11555 D.t81 7.599
R11637 D.n11575 D.t467 7.599
R11638 D.n11595 D.t1108 7.599
R11639 D.n11615 D.t2279 7.599
R11640 D.n11635 D.t978 7.599
R11641 D.n11655 D.t3184 7.599
R11642 D.n11675 D.t1065 7.599
R11643 D.n11695 D.t858 7.599
R11644 D.n11715 D.t2506 7.599
R11645 D.n11735 D.t3119 7.599
R11646 D.n11755 D.t4101 7.599
R11647 D.n11775 D.t3262 7.599
R11648 D.n11795 D.t1988 7.599
R11649 D.n11815 D.t3313 7.599
R11650 D.n11835 D.t181 7.599
R11651 D.n11823 D.t4504 7.599
R11652 D.n11803 D.t2902 7.599
R11653 D.n11783 D.t2991 7.599
R11654 D.n11763 D.t2485 7.599
R11655 D.n11743 D.t2078 7.599
R11656 D.n11723 D.t2820 7.599
R11657 D.n11703 D.t2773 7.599
R11658 D.n11683 D.t822 7.599
R11659 D.n11663 D.t789 7.599
R11660 D.n11643 D.t1955 7.599
R11661 D.n11623 D.t1056 7.599
R11662 D.n11603 D.t1405 7.599
R11663 D.n11583 D.t259 7.599
R11664 D.n11563 D.t1052 7.599
R11665 D.n11543 D.t2444 7.599
R11666 D.n11523 D.t4086 7.599
R11667 D.n11500 D.t1501 7.599
R11668 D.n11490 D.t1101 7.599
R11669 D.n11414 D.t3654 7.599
R11670 D.n11396 D.t3709 7.599
R11671 D.n11378 D.t3104 7.599
R11672 D.n11360 D.t3163 7.599
R11673 D.n11342 D.t4276 7.599
R11674 D.n11324 D.t3604 7.599
R11675 D.n11306 D.t85 7.599
R11676 D.n11288 D.t3216 7.599
R11677 D.n11270 D.t312 7.599
R11678 D.n11252 D.t1210 7.599
R11679 D.n11234 D.t2246 7.599
R11680 D.n11216 D.t3936 7.599
R11681 D.n11198 D.t4251 7.599
R11682 D.n11180 D.t968 7.599
R11683 D.n11162 D.t3575 7.599
R11684 D.n11143 D.t3171 7.599
R11685 D.n11152 D.t558 7.599
R11686 D.n11170 D.t3814 7.599
R11687 D.n11188 D.t2118 7.599
R11688 D.n11206 D.t176 7.599
R11689 D.n11224 D.t4001 7.599
R11690 D.n11242 D.t1717 7.599
R11691 D.n11260 D.t1288 7.599
R11692 D.n11278 D.t607 7.599
R11693 D.n11296 D.t3923 7.599
R11694 D.n11314 D.t3286 7.599
R11695 D.n11332 D.t3147 7.599
R11696 D.n11350 D.t4056 7.599
R11697 D.n11368 D.t4302 7.599
R11698 D.n11386 D.t4187 7.599
R11699 D.n11404 D.t2470 7.599
R11700 D.n11426 D.t2433 7.599
R11701 D.n11443 D.t2877 7.599
R11702 D.n10792 D.t3277 7.599
R11703 D.n10812 D.t471 7.599
R11704 D.n10832 D.t1290 7.599
R11705 D.n10852 D.t1537 7.599
R11706 D.n10872 D.t554 7.599
R11707 D.n10892 D.t3072 7.599
R11708 D.n10912 D.t3059 7.599
R11709 D.n10932 D.t2865 7.599
R11710 D.n10952 D.t3150 7.599
R11711 D.n10972 D.t143 7.599
R11712 D.n10992 D.t563 7.599
R11713 D.n11012 D.t1234 7.599
R11714 D.n11032 D.t4328 7.599
R11715 D.n11052 D.t3564 7.599
R11716 D.n11072 D.t4395 7.599
R11717 D.n11060 D.t2023 7.599
R11718 D.n11040 D.t108 7.599
R11719 D.n11020 D.t4018 7.599
R11720 D.n11000 D.t4170 7.599
R11721 D.n10980 D.t2518 7.599
R11722 D.n10960 D.t1107 7.599
R11723 D.n10940 D.t119 7.599
R11724 D.n10920 D.t859 7.599
R11725 D.n10900 D.t3903 7.599
R11726 D.n10880 D.t1349 7.599
R11727 D.n10860 D.t1572 7.599
R11728 D.n10840 D.t848 7.599
R11729 D.n10820 D.t1919 7.599
R11730 D.n10800 D.t2492 7.599
R11731 D.n10777 D.t3977 7.599
R11732 D.n10767 D.t1824 7.599
R11733 D.n10695 D.t1025 7.599
R11734 D.n10677 D.t1759 7.599
R11735 D.n10659 D.t68 7.599
R11736 D.n10641 D.t4059 7.599
R11737 D.n10623 D.t185 7.599
R11738 D.n10605 D.t1211 7.599
R11739 D.n10587 D.t2352 7.599
R11740 D.n10569 D.t660 7.599
R11741 D.n10551 D.t2423 7.599
R11742 D.n10533 D.t3643 7.599
R11743 D.n10515 D.t2103 7.599
R11744 D.n10497 D.t1323 7.599
R11745 D.n10479 D.t3780 7.599
R11746 D.n10460 D.t324 7.599
R11747 D.n10469 D.t1216 7.599
R11748 D.n10487 D.t4312 7.599
R11749 D.n10505 D.t1928 7.599
R11750 D.n10523 D.t229 7.599
R11751 D.n10541 D.t1522 7.599
R11752 D.n10559 D.t351 7.599
R11753 D.n10577 D.t3231 7.599
R11754 D.n10595 D.t4112 7.599
R11755 D.n10613 D.t3464 7.599
R11756 D.n10631 D.t3911 7.599
R11757 D.n10649 D.t1794 7.599
R11758 D.n10667 D.t2566 7.599
R11759 D.n10685 D.t2656 7.599
R11760 D.n10707 D.t1954 7.599
R11761 D.n10724 D.t3690 7.599
R11762 D.n10149 D.t3879 7.599
R11763 D.n10169 D.t4426 7.599
R11764 D.n10189 D.t2933 7.599
R11765 D.n10209 D.t574 7.599
R11766 D.n10229 D.t367 7.599
R11767 D.n10249 D.t359 7.599
R11768 D.n10269 D.t3034 7.599
R11769 D.n10289 D.t2679 7.599
R11770 D.n10309 D.t156 7.599
R11771 D.n10329 D.t3765 7.599
R11772 D.n10349 D.t2175 7.599
R11773 D.n10369 D.t2274 7.599
R11774 D.n10389 D.t828 7.599
R11775 D.n10377 D.t3065 7.599
R11776 D.n10357 D.t640 7.599
R11777 D.n10337 D.t1360 7.599
R11778 D.n10317 D.t2 7.599
R11779 D.n10297 D.t1468 7.599
R11780 D.n10277 D.t3401 7.599
R11781 D.n10257 D.t3361 7.599
R11782 D.n10237 D.t3672 7.599
R11783 D.n10217 D.t240 7.599
R11784 D.n10197 D.t4366 7.599
R11785 D.n10177 D.t4238 7.599
R11786 D.n10157 D.t4074 7.599
R11787 D.n10132 D.t1995 7.599
R11788 D.n10119 D.t1149 7.599
R11789 D.n10056 D.t1489 7.599
R11790 D.n10038 D.t1604 7.599
R11791 D.n10020 D.t1729 7.599
R11792 D.n10002 D.t3123 7.599
R11793 D.n9984 D.t2919 7.599
R11794 D.n9966 D.t3060 7.599
R11795 D.n9948 D.t3050 7.599
R11796 D.n9930 D.t3052 7.599
R11797 D.n9912 D.t2888 7.599
R11798 D.n9894 D.t3092 7.599
R11799 D.n9876 D.t4360 7.599
R11800 D.n9857 D.t1663 7.599
R11801 D.n9866 D.t2344 7.599
R11802 D.n9884 D.t7 7.599
R11803 D.n9902 D.t1379 7.599
R11804 D.n9920 D.t537 7.599
R11805 D.n9938 D.t3661 7.599
R11806 D.n9956 D.t2576 7.599
R11807 D.n9974 D.t1981 7.599
R11808 D.n9992 D.t310 7.599
R11809 D.n10010 D.t1844 7.599
R11810 D.n10028 D.t456 7.599
R11811 D.n10046 D.t2482 7.599
R11812 D.n10067 D.t716 7.599
R11813 D.n10078 D.t2960 7.599
R11814 D.n9586 D.t1033 7.599
R11815 D.n9606 D.t2027 7.599
R11816 D.n9626 D.t2237 7.599
R11817 D.n9646 D.t2382 7.599
R11818 D.n9666 D.t273 7.599
R11819 D.n9686 D.t987 7.599
R11820 D.n9706 D.t2257 7.599
R11821 D.n9726 D.t2434 7.599
R11822 D.n9746 D.t1660 7.599
R11823 D.n9766 D.t3679 7.599
R11824 D.n9786 D.t1978 7.599
R11825 D.n9774 D.t2180 7.599
R11826 D.n9754 D.t3725 7.599
R11827 D.n9734 D.t1165 7.599
R11828 D.n9714 D.t1276 7.599
R11829 D.n9694 D.t4135 7.599
R11830 D.n9674 D.t3856 7.599
R11831 D.n9654 D.t3897 7.599
R11832 D.n9634 D.t758 7.599
R11833 D.n9614 D.t3785 7.599
R11834 D.n9594 D.t2612 7.599
R11835 D.n9569 D.t526 7.599
R11836 D.n9556 D.t1226 7.599
R11837 D.n9491 D.t3992 7.599
R11838 D.n9473 D.t2153 7.599
R11839 D.n9455 D.t2205 7.599
R11840 D.n9437 D.t4509 7.599
R11841 D.n9419 D.t1225 7.599
R11842 D.n9401 D.t2626 7.599
R11843 D.n9383 D.t132 7.599
R11844 D.n9365 D.t91 7.599
R11845 D.n9347 D.t2659 7.599
R11846 D.n9328 D.t2682 7.599
R11847 D.n9337 D.t1395 7.599
R11848 D.n9355 D.t795 7.599
R11849 D.n9373 D.t3351 7.599
R11850 D.n9391 D.t3222 7.599
R11851 D.n9409 D.t3460 7.599
R11852 D.n9427 D.t1722 7.599
R11853 D.n9445 D.t1419 7.599
R11854 D.n9463 D.t3478 7.599
R11855 D.n9481 D.t3678 7.599
R11856 D.n9503 D.t4455 7.599
R11857 D.n9520 D.t1484 7.599
R11858 D.n9097 D.t803 7.599
R11859 D.n9117 D.t1363 7.599
R11860 D.n9137 D.t561 7.599
R11861 D.n9157 D.t3102 7.599
R11862 D.n9177 D.t2795 7.599
R11863 D.n9197 D.t2908 7.599
R11864 D.n9217 D.t3073 7.599
R11865 D.n9237 D.t2953 7.599
R11866 D.n9257 D.t2915 7.599
R11867 D.n9245 D.t2008 7.599
R11868 D.n9225 D.t3315 7.599
R11869 D.n9205 D.t4142 7.599
R11870 D.n9185 D.t3384 7.599
R11871 D.n9165 D.t1268 7.599
R11872 D.n9145 D.t1813 7.599
R11873 D.n9125 D.t4105 7.599
R11874 D.n9105 D.t3194 7.599
R11875 D.n9082 D.t496 7.599
R11876 D.n9072 D.t4266 7.599
R11877 D.n9012 D.t1775 7.599
R11878 D.n8994 D.t1951 7.599
R11879 D.n8976 D.t2135 7.599
R11880 D.n8958 D.t2367 7.599
R11881 D.n8940 D.t2317 7.599
R11882 D.n8922 D.t838 7.599
R11883 D.n8904 D.t2250 7.599
R11884 D.n8885 D.t1046 7.599
R11885 D.n8894 D.t3859 7.599
R11886 D.n8912 D.t3416 7.599
R11887 D.n8930 D.t2033 7.599
R11888 D.n8948 D.t2305 7.599
R11889 D.n8966 D.t1045 7.599
R11890 D.n8984 D.t3965 7.599
R11891 D.n9002 D.t3325 7.599
R11892 D.n9024 D.t4430 7.599
R11893 D.n9041 D.t2270 7.599
R11894 D.n8694 D.t2548 7.599
R11895 D.n8714 D.t4031 7.599
R11896 D.n8734 D.t2197 7.599
R11897 D.n8754 D.t4494 7.599
R11898 D.n8774 D.t1655 7.599
R11899 D.n8794 D.t1541 7.599
R11900 D.n8814 D.t4501 7.599
R11901 D.n8802 D.t3819 7.599
R11902 D.n8782 D.t4076 7.599
R11903 D.n8762 D.t1377 7.599
R11904 D.n8742 D.t349 7.599
R11905 D.n8722 D.t3671 7.599
R11906 D.n8702 D.t3405 7.599
R11907 D.n8677 D.t853 7.599
R11908 D.n8664 D.t3055 7.599
R11909 D.n8613 D.t2567 7.599
R11910 D.n8595 D.t737 7.599
R11911 D.n8577 D.t544 7.599
R11912 D.n8559 D.t3027 7.599
R11913 D.n8541 D.t2873 7.599
R11914 D.n8522 D.t548 7.599
R11915 D.n8531 D.t1948 7.599
R11916 D.n8549 D.t363 7.599
R11917 D.n8567 D.t1467 7.599
R11918 D.n8585 D.t3403 7.599
R11919 D.n8603 D.t2647 7.599
R11920 D.n8624 D.t2769 7.599
R11921 D.n8635 D.t1032 7.599
R11922 D.n8371 D.t1533 7.599
R11923 D.n8391 D.t1513 7.599
R11924 D.n8411 D.t2123 7.599
R11925 D.n8431 D.t2364 7.599
R11926 D.n8451 D.t1799 7.599
R11927 D.n8439 D.t3485 7.599
R11928 D.n8419 D.t1858 7.599
R11929 D.n8399 D.t3771 7.599
R11930 D.n8379 D.t3939 7.599
R11931 D.n8354 D.t4109 7.599
R11932 D.n8341 D.t906 7.599
R11933 D.n8288 D.t2531 7.599
R11934 D.n8270 D.t4022 7.599
R11935 D.n8252 D.t2192 7.599
R11936 D.n8233 D.t2537 7.599
R11937 D.n8242 D.t3459 7.599
R11938 D.n8260 D.t3297 7.599
R11939 D.n8278 D.t3466 7.599
R11940 D.n8300 D.t2222 7.599
R11941 D.n8317 D.t3829 7.599
R11942 D.n8122 D.t2326 7.599
R11943 D.n8142 D.t678 7.599
R11944 D.n8162 D.t1330 7.599
R11945 D.n8150 D.t513 7.599
R11946 D.n8130 D.t3301 7.599
R11947 D.n8107 D.t4297 7.599
R11948 D.n8097 D.t1865 7.599
R11949 D.n8049 D.t655 7.599
R11950 D.n8030 D.t674 7.599
R11951 D.n8039 D.t4122 7.599
R11952 D.n8061 D.t446 7.599
R11953 D.n8078 D.t2179 7.599
R11954 D.n7909 D.t3851 7.599
R11955 D.n50 D.t553 7.599
R11956 D.n59 D.t3334 7.599
R11957 D.n68 D.t2435 7.599
R11958 D.n77 D.t2947 7.599
R11959 D.n86 D.t1517 7.599
R11960 D.n95 D.t1495 7.599
R11961 D.n104 D.t3617 7.599
R11962 D.n113 D.t2469 7.599
R11963 D.n122 D.t4377 7.599
R11964 D.n131 D.t3000 7.599
R11965 D.n140 D.t2627 7.599
R11966 D.n149 D.t971 7.599
R11967 D.n158 D.t3800 7.599
R11968 D.n167 D.t1324 7.599
R11969 D.n176 D.t405 7.599
R11970 D.n185 D.t2677 7.599
R11971 D.n194 D.t896 7.599
R11972 D.n203 D.t3603 7.599
R11973 D.n212 D.t219 7.599
R11974 D.n221 D.t336 7.599
R11975 D.n230 D.t4376 7.599
R11976 D.n239 D.t1859 7.599
R11977 D.n248 D.t3675 7.599
R11978 D.n257 D.t83 7.599
R11979 D.n266 D.t2093 7.599
R11980 D.n275 D.t3067 7.599
R11981 D.n284 D.t31 7.599
R11982 D.n293 D.t293 7.599
R11983 D.n302 D.t4323 7.599
R11984 D.n311 D.t1969 7.599
R11985 D.n320 D.t4203 7.599
R11986 D.n329 D.t493 7.599
R11987 D.n338 D.t3754 7.599
R11988 D.n347 D.t612 7.599
R11989 D.n356 D.t2793 7.599
R11990 D.n365 D.t1911 7.599
R11991 D.n374 D.t3712 7.599
R11992 D.n383 D.t2581 7.599
R11993 D.n392 D.t4102 7.599
R11994 D.n401 D.t715 7.599
R11995 D.n410 D.t4080 7.599
R11996 D.n419 D.t1685 7.599
R11997 D.n428 D.t3707 7.599
R11998 D.n523 D.t672 7.599
R11999 D.n539 D.t609 7.599
R12000 D.n1127 D.t1399 7.599
R12001 D.n1113 D.t2831 7.599
R12002 D.n1099 D.t3574 7.599
R12003 D.n1085 D.t3591 7.599
R12004 D.n1071 D.t711 7.599
R12005 D.n1057 D.t1194 7.599
R12006 D.n1043 D.t2378 7.599
R12007 D.n1029 D.t1510 7.599
R12008 D.n1015 D.t3423 7.599
R12009 D.n1001 D.t3486 7.599
R12010 D.n987 D.t3107 7.599
R12011 D.n973 D.t652 7.599
R12012 D.n959 D.t929 7.599
R12013 D.n945 D.t2167 7.599
R12014 D.n931 D.t1890 7.599
R12015 D.n917 D.t3183 7.599
R12016 D.n903 D.t1031 7.599
R12017 D.n889 D.t2430 7.599
R12018 D.n875 D.t2927 7.599
R12019 D.n861 D.t1167 7.599
R12020 D.n847 D.t360 7.599
R12021 D.n833 D.t3615 7.599
R12022 D.n819 D.t3185 7.599
R12023 D.n805 D.t3040 7.599
R12024 D.n791 D.t1609 7.599
R12025 D.n777 D.t3412 7.599
R12026 D.n763 D.t2539 7.599
R12027 D.n749 D.t2381 7.599
R12028 D.n735 D.t3300 7.599
R12029 D.n721 D.t266 7.599
R12030 D.n707 D.t3462 7.599
R12031 D.n693 D.t1311 7.599
R12032 D.n679 D.t3720 7.599
R12033 D.n665 D.t2665 7.599
R12034 D.n651 D.t3950 7.599
R12035 D.n637 D.t1638 7.599
R12036 D.n623 D.t1386 7.599
R12037 D.n609 D.t437 7.599
R12038 D.n595 D.t1705 7.599
R12039 D.n581 D.t1982 7.599
R12040 D.n567 D.t427 7.599
R12041 D.n553 D.t1133 7.599
R12042 D.n1150 D.t3777 7.599
R12043 D.n1166 D.t1347 7.599
R12044 D.n1726 D.t1903 7.599
R12045 D.n1712 D.t4104 7.599
R12046 D.n1698 D.t958 7.599
R12047 D.n1684 D.t570 7.599
R12048 D.n1670 D.t3753 7.599
R12049 D.n1656 D.t1461 7.599
R12050 D.n1642 D.t3322 7.599
R12051 D.n1628 D.t3224 7.599
R12052 D.n1614 D.t1726 7.599
R12053 D.n1600 D.t104 7.599
R12054 D.n1586 D.t2049 7.599
R12055 D.n1572 D.t2280 7.599
R12056 D.n1558 D.t4398 7.599
R12057 D.n1544 D.t2073 7.599
R12058 D.n1530 D.t1307 7.599
R12059 D.n1516 D.t3146 7.599
R12060 D.n1502 D.t244 7.599
R12061 D.n1488 D.t1492 7.599
R12062 D.n1474 D.t707 7.599
R12063 D.n1460 D.t1182 7.599
R12064 D.n1446 D.t2781 7.599
R12065 D.n1432 D.t2297 7.599
R12066 D.n1418 D.t3599 7.599
R12067 D.n1404 D.t3738 7.599
R12068 D.n1390 D.t1085 7.599
R12069 D.n1376 D.t2883 7.599
R12070 D.n1362 D.t1503 7.599
R12071 D.n1348 D.t812 7.599
R12072 D.n1334 D.t3743 7.599
R12073 D.n1320 D.t872 7.599
R12074 D.n1306 D.t4103 7.599
R12075 D.n1292 D.t1922 7.599
R12076 D.n1278 D.t3441 7.599
R12077 D.n1264 D.t3830 7.599
R12078 D.n1250 D.t4472 7.599
R12079 D.n1236 D.t3436 7.599
R12080 D.n1222 D.t736 7.599
R12081 D.n1208 D.t3363 7.599
R12082 D.n1194 D.t205 7.599
R12083 D.n1180 D.t3673 7.599
R12084 D.n1749 D.t3465 7.599
R12085 D.n1765 D.t2543 7.599
R12086 D.n2297 D.t680 7.599
R12087 D.n2283 D.t1694 7.599
R12088 D.n2269 D.t894 7.599
R12089 D.n2255 D.t4129 7.599
R12090 D.n2241 D.t139 7.599
R12091 D.n2227 D.t1451 7.599
R12092 D.n2213 D.t4510 7.599
R12093 D.n2199 D.t2361 7.599
R12094 D.n2185 D.t3714 7.599
R12095 D.n2171 D.t1321 7.599
R12096 D.n2157 D.t3741 7.599
R12097 D.n2143 D.t1188 7.599
R12098 D.n2129 D.t3098 7.599
R12099 D.n2115 D.t100 7.599
R12100 D.n2101 D.t1902 7.599
R12101 D.n2087 D.t4292 7.599
R12102 D.n2073 D.t625 7.599
R12103 D.n2059 D.t646 7.599
R12104 D.n2045 D.t3836 7.599
R12105 D.n2031 D.t2400 7.599
R12106 D.n2017 D.t3427 7.599
R12107 D.n2003 D.t1131 7.599
R12108 D.n1989 D.t1525 7.599
R12109 D.n1975 D.t2693 7.599
R12110 D.n1961 D.t2429 7.599
R12111 D.n1947 D.t4311 7.599
R12112 D.n1933 D.t877 7.599
R12113 D.n1919 D.t3728 7.599
R12114 D.n1905 D.t3957 7.599
R12115 D.n1891 D.t4249 7.599
R12116 D.n1877 D.t1983 7.599
R12117 D.n1863 D.t4306 7.599
R12118 D.n1849 D.t2414 7.599
R12119 D.n1835 D.t3773 7.599
R12120 D.n1821 D.t2195 7.599
R12121 D.n1807 D.t4385 7.599
R12122 D.n1793 D.t4028 7.599
R12123 D.n1779 D.t3534 7.599
R12124 D.n2320 D.t3904 7.599
R12125 D.n2336 D.t1869 7.599
R12126 D.n2840 D.t2712 7.599
R12127 D.n2826 D.t14 7.599
R12128 D.n2812 D.t1863 7.599
R12129 D.n2798 D.t1371 7.599
R12130 D.n2784 D.t487 7.599
R12131 D.n2770 D.t2754 7.599
R12132 D.n2756 D.t1118 7.599
R12133 D.n2742 D.t1425 7.599
R12134 D.n2728 D.t4437 7.599
R12135 D.n2714 D.t3978 7.599
R12136 D.n2700 D.t4060 7.599
R12137 D.n2686 D.t1212 7.599
R12138 D.n2672 D.t4285 7.599
R12139 D.n2658 D.t3487 7.599
R12140 D.n2644 D.t675 7.599
R12141 D.n2630 D.t3766 7.599
R12142 D.n2616 D.t636 7.599
R12143 D.n2602 D.t3153 7.599
R12144 D.n2588 D.t111 7.599
R12145 D.n2574 D.t1458 7.599
R12146 D.n2560 D.t53 7.599
R12147 D.n2546 D.t2348 7.599
R12148 D.n2532 D.t2943 7.599
R12149 D.n2518 D.t483 7.599
R12150 D.n2504 D.t1491 7.599
R12151 D.n2490 D.t3596 7.599
R12152 D.n2476 D.t1113 7.599
R12153 D.n2462 D.t2812 7.599
R12154 D.n2448 D.t3364 7.599
R12155 D.n2434 D.t2022 7.599
R12156 D.n2420 D.t2948 7.599
R12157 D.n2406 D.t1153 7.599
R12158 D.n2392 D.t2366 7.599
R12159 D.n2378 D.t2259 7.599
R12160 D.n2364 D.t2128 7.599
R12161 D.n2350 D.t107 7.599
R12162 D.n2863 D.t3346 7.599
R12163 D.n2879 D.t560 7.599
R12164 D.n3355 D.t3244 7.599
R12165 D.n3341 D.t459 7.599
R12166 D.n3327 D.t1915 7.599
R12167 D.n3313 D.t297 7.599
R12168 D.n3299 D.t433 7.599
R12169 D.n3285 D.t4327 7.599
R12170 D.n3271 D.t1150 7.599
R12171 D.n3257 D.t3396 7.599
R12172 D.n3243 D.t4489 7.599
R12173 D.n3229 D.t1747 7.599
R12174 D.n3215 D.t2254 7.599
R12175 D.n3201 D.t2551 7.599
R12176 D.n3187 D.t2189 7.599
R12177 D.n3173 D.t2289 7.599
R12178 D.n3159 D.t1570 7.599
R12179 D.n3145 D.t1562 7.599
R12180 D.n3131 D.t1857 7.599
R12181 D.n3117 D.t3537 7.599
R12182 D.n3103 D.t145 7.599
R12183 D.n3089 D.t2783 7.599
R12184 D.n3075 D.t172 7.599
R12185 D.n3061 D.t1411 7.599
R12186 D.n3047 D.t3508 7.599
R12187 D.n3033 D.t3637 7.599
R12188 D.n3019 D.t608 7.599
R12189 D.n3005 D.t1670 7.599
R12190 D.n2991 D.t1827 7.599
R12191 D.n2977 D.t1961 7.599
R12192 D.n2963 D.t3206 7.599
R12193 D.n2949 D.t3383 7.599
R12194 D.n2935 D.t2826 7.599
R12195 D.n2921 D.t3311 7.599
R12196 D.n2907 D.t3085 7.599
R12197 D.n2893 D.t3815 7.599
R12198 D.n3379 D.t3843 7.599
R12199 D.n3395 D.t4505 7.599
R12200 D.n3843 D.t2171 7.599
R12201 D.n3829 D.t217 7.599
R12202 D.n3815 D.t117 7.599
R12203 D.n3801 D.t3215 7.599
R12204 D.n3787 D.t1800 7.599
R12205 D.n3773 D.t422 7.599
R12206 D.n3759 D.t384 7.599
R12207 D.n3745 D.t211 7.599
R12208 D.n3731 D.t30 7.599
R12209 D.n3717 D.t746 7.599
R12210 D.n3703 D.t2359 7.599
R12211 D.n3689 D.t3669 7.599
R12212 D.n3675 D.t2614 7.599
R12213 D.n3661 D.t839 7.599
R12214 D.n3647 D.t4248 7.599
R12215 D.n3633 D.t3200 7.599
R12216 D.n3619 D.t404 7.599
R12217 D.n3605 D.t2144 7.599
R12218 D.n3591 D.t3824 7.599
R12219 D.n3577 D.t4358 7.599
R12220 D.n3563 D.t78 7.599
R12221 D.n3549 D.t3242 7.599
R12222 D.n3535 D.t1689 7.599
R12223 D.n3521 D.t2215 7.599
R12224 D.n3507 D.t3039 7.599
R12225 D.n3493 D.t2987 7.599
R12226 D.n3479 D.t300 7.599
R12227 D.n3465 D.t617 7.599
R12228 D.n3451 D.t2683 7.599
R12229 D.n3437 D.t3568 7.599
R12230 D.n3423 D.t901 7.599
R12231 D.n3409 D.t3963 7.599
R12232 D.n3867 D.t1676 7.599
R12233 D.n3883 D.t3210 7.599
R12234 D.n4303 D.t2136 7.599
R12235 D.n4289 D.t3627 7.599
R12236 D.n4275 D.t4270 7.599
R12237 D.n4261 D.t1160 7.599
R12238 D.n4247 D.t2571 7.599
R12239 D.n4233 D.t4110 7.599
R12240 D.n4219 D.t2402 7.599
R12241 D.n4205 D.t889 7.599
R12242 D.n4191 D.t1511 7.599
R12243 D.n4177 D.t1088 7.599
R12244 D.n4163 D.t599 7.599
R12245 D.n4149 D.t2969 7.599
R12246 D.n4135 D.t641 7.599
R12247 D.n4121 D.t1649 7.599
R12248 D.n4107 D.t2166 7.599
R12249 D.n4093 D.t3269 7.599
R12250 D.n4079 D.t1 7.599
R12251 D.n4065 D.t2145 7.599
R12252 D.n4051 D.t1538 7.599
R12253 D.n4037 D.t418 7.599
R12254 D.n4023 D.t2321 7.599
R12255 D.n4009 D.t3008 7.599
R12256 D.n3995 D.t44 7.599
R12257 D.n3981 D.t748 7.599
R12258 D.n3967 D.t225 7.599
R12259 D.n3953 D.t3246 7.599
R12260 D.n3939 D.t2372 7.599
R12261 D.n3925 D.t3480 7.599
R12262 D.n3911 D.t985 7.599
R12263 D.n3897 D.t2631 7.599
R12264 D.n4327 D.t3611 7.599
R12265 D.n4343 D.t3080 7.599
R12266 D.n4735 D.t520 7.599
R12267 D.n4721 D.t919 7.599
R12268 D.n4707 D.t4039 7.599
R12269 D.n4693 D.t1239 7.599
R12270 D.n4679 D.t3007 7.599
R12271 D.n4665 D.t3987 7.599
R12272 D.n4651 D.t1460 7.599
R12273 D.n4637 D.t4347 7.599
R12274 D.n4623 D.t3223 7.599
R12275 D.n4609 D.t1270 7.599
R12276 D.n4595 D.t3732 7.599
R12277 D.n4581 D.t4405 7.599
R12278 D.n4567 D.t2276 7.599
R12279 D.n4553 D.t3047 7.599
R12280 D.n4539 D.t2072 7.599
R12281 D.n4525 D.t342 7.599
R12282 D.n4511 D.t4275 7.599
R12283 D.n4497 D.t518 7.599
R12284 D.n4483 D.t2568 7.599
R12285 D.n4469 D.t2662 7.599
R12286 D.n4455 D.t3840 7.599
R12287 D.n4441 D.t1078 7.599
R12288 D.n4427 D.t4173 7.599
R12289 D.n4413 D.t1002 7.599
R12290 D.n4399 D.t843 7.599
R12291 D.n4385 D.t2554 7.599
R12292 D.n4371 D.t1921 7.599
R12293 D.n4357 D.t2996 7.599
R12294 D.n4759 D.t4424 7.599
R12295 D.n4775 D.t3715 7.599
R12296 D.n5139 D.t2225 7.599
R12297 D.n5125 D.t3425 7.599
R12298 D.n5111 D.t501 7.599
R12299 D.n5097 D.t2014 7.599
R12300 D.n5083 D.t4239 7.599
R12301 D.n5069 D.t2669 7.599
R12302 D.n5055 D.t1436 7.599
R12303 D.n5041 D.t3081 7.599
R12304 D.n5027 D.t2353 7.599
R12305 D.n5013 D.t692 7.599
R12306 D.n4999 D.t3155 7.599
R12307 D.n4985 D.t1357 7.599
R12308 D.n4971 D.t1187 7.599
R12309 D.n4957 D.t4375 7.599
R12310 D.n4943 D.t2282 7.599
R12311 D.n4929 D.t3676 7.599
R12312 D.n4915 D.t4029 7.599
R12313 D.n4901 D.t1100 7.599
R12314 D.n4887 D.t4354 7.599
R12315 D.n4873 D.t3025 7.599
R12316 D.n4859 D.t194 7.599
R12317 D.n4845 D.t1205 7.599
R12318 D.n4831 D.t3997 7.599
R12319 D.n4817 D.t316 7.599
R12320 D.n4803 D.t2680 7.599
R12321 D.n4789 D.t96 7.599
R12322 D.n5163 D.t1021 7.599
R12323 D.n5179 D.t3017 7.599
R12324 D.n5515 D.t857 7.599
R12325 D.n5501 D.t1728 7.599
R12326 D.n5487 D.t3203 7.599
R12327 D.n5473 D.t2383 7.599
R12328 D.n5459 D.t3169 7.599
R12329 D.n5445 D.t1181 7.599
R12330 D.n5431 D.t2799 7.599
R12331 D.n5417 D.t2524 7.599
R12332 D.n5403 D.t1424 7.599
R12333 D.n5389 D.t2930 7.599
R12334 D.n5375 D.t4231 7.599
R12335 D.n5361 D.t2634 7.599
R12336 D.n5347 D.t3420 7.599
R12337 D.n5333 D.t3762 7.599
R12338 D.n5319 D.t2132 7.599
R12339 D.n5305 D.t2986 7.599
R12340 D.n5291 D.t956 7.599
R12341 D.n5277 D.t1535 7.599
R12342 D.n5263 D.t2483 7.599
R12343 D.n5249 D.t3159 7.599
R12344 D.n5235 D.t2019 7.599
R12345 D.n5221 D.t726 7.599
R12346 D.n5207 D.t2720 7.599
R12347 D.n5193 D.t2332 7.599
R12348 D.n5539 D.t964 7.599
R12349 D.n5555 D.t1264 7.599
R12350 D.n5863 D.t1650 7.599
R12351 D.n5849 D.t3857 7.599
R12352 D.n5835 D.t2006 7.599
R12353 D.n5821 D.t3975 7.599
R12354 D.n5807 D.t2239 7.599
R12355 D.n5793 D.t1506 7.599
R12356 D.n5779 D.t4460 7.599
R12357 D.n5765 D.t1201 7.599
R12358 D.n5751 D.t3395 7.599
R12359 D.n5737 D.t2051 7.599
R12360 D.n5723 D.t3764 7.599
R12361 D.n5709 D.t1829 7.599
R12362 D.n5695 D.t3097 7.599
R12363 D.n5681 D.t4062 7.599
R12364 D.n5667 D.t2493 7.599
R12365 D.n5653 D.t2421 7.599
R12366 D.n5639 D.t4235 7.599
R12367 D.n5625 D.t835 7.599
R12368 D.n5611 D.t1664 7.599
R12369 D.n5597 D.t2062 7.599
R12370 D.n5583 D.t2463 7.599
R12371 D.n5569 D.t2994 7.599
R12372 D.n5887 D.t2858 7.599
R12373 D.n5903 D.t3882 7.599
R12374 D.n6183 D.t4139 7.599
R12375 D.n6169 D.t3333 7.599
R12376 D.n6155 D.t3270 7.599
R12377 D.n6141 D.t579 7.599
R12378 D.n6127 D.t2703 7.599
R12379 D.n6113 D.t3850 7.599
R12380 D.n6099 D.t421 7.599
R12381 D.n6085 D.t2579 7.599
R12382 D.n6071 D.t3058 7.599
R12383 D.n6057 D.t124 7.599
R12384 D.n6043 D.t2760 7.599
R12385 D.n6029 D.t662 7.599
R12386 D.n6015 D.t4192 7.599
R12387 D.n6001 D.t2805 7.599
R12388 D.n5987 D.t3188 7.599
R12389 D.n5973 D.t1493 7.599
R12390 D.n5959 D.t684 7.599
R12391 D.n5945 D.t988 7.599
R12392 D.n5931 D.t2303 7.599
R12393 D.n5917 D.t653 7.599
R12394 D.n6207 D.t1209 7.599
R12395 D.n6223 D.t3069 7.599
R12396 D.n6475 D.t3149 7.599
R12397 D.n6461 D.t4491 7.599
R12398 D.n6447 D.t743 7.599
R12399 D.n6433 D.t4124 7.599
R12400 D.n6419 D.t1964 7.599
R12401 D.n6405 D.t1599 7.599
R12402 D.n6391 D.t2623 7.599
R12403 D.n6377 D.t1446 7.599
R12404 D.n6363 D.t3327 7.599
R12405 D.n6349 D.t397 7.599
R12406 D.n6335 D.t1051 7.599
R12407 D.n6321 D.t169 7.599
R12408 D.n6307 D.t786 7.599
R12409 D.n6293 D.t3567 7.599
R12410 D.n6279 D.t3273 7.599
R12411 D.n6265 D.t647 7.599
R12412 D.n6251 D.t2763 7.599
R12413 D.n6237 D.t1480 7.599
R12414 D.n6499 D.t3665 7.599
R12415 D.n6515 D.t1846 7.599
R12416 D.n6739 D.t4434 7.599
R12417 D.n6725 D.t1128 7.599
R12418 D.n6711 D.t4149 7.599
R12419 D.n6697 D.t4470 7.599
R12420 D.n6683 D.t2586 7.599
R12421 D.n6669 D.t3797 7.599
R12422 D.n6655 D.t1765 7.599
R12423 D.n6641 D.t2590 7.599
R12424 D.n6627 D.t356 7.599
R12425 D.n6613 D.t4440 7.599
R12426 D.n6599 D.t3688 7.599
R12427 D.n6585 D.t69 7.599
R12428 D.n6571 D.t3121 7.599
R12429 D.n6557 D.t1690 7.599
R12430 D.n6543 D.t883 7.599
R12431 D.n6529 D.t2776 7.599
R12432 D.n6763 D.t3531 7.599
R12433 D.n6779 D.t3406 7.599
R12434 D.n6975 D.t3787 7.599
R12435 D.n6961 D.t2410 7.599
R12436 D.n6947 D.t2928 7.599
R12437 D.n6933 D.t27 7.599
R12438 D.n6919 D.t924 7.599
R12439 D.n6905 D.t3706 7.599
R12440 D.n6891 D.t2597 7.599
R12441 D.n6877 D.t2258 7.599
R12442 D.n6863 D.t729 7.599
R12443 D.n6849 D.t2191 7.599
R12444 D.n6835 D.t514 7.599
R12445 D.n6821 D.t2337 7.599
R12446 D.n6807 D.t4178 7.599
R12447 D.n6793 D.t43 7.599
R12448 D.n6999 D.t19 7.599
R12449 D.n7015 D.t3967 7.599
R12450 D.n7183 D.t3253 7.599
R12451 D.n7169 D.t2516 7.599
R12452 D.n7155 D.t4212 7.599
R12453 D.n7141 D.t540 7.599
R12454 D.n7127 D.t3367 7.599
R12455 D.n7113 D.t3310 7.599
R12456 D.n7099 D.t2066 7.599
R12457 D.n7085 D.t2356 7.599
R12458 D.n7071 D.t3043 7.599
R12459 D.n7057 D.t2621 7.599
R12460 D.n7043 D.t2012 7.599
R12461 D.n7029 D.t3841 7.599
R12462 D.n7207 D.t381 7.599
R12463 D.n7223 D.t1822 7.599
R12464 D.n7363 D.t1576 7.599
R12465 D.n7349 D.t3385 7.599
R12466 D.n7335 D.t3448 7.599
R12467 D.n7321 D.t4066 7.599
R12468 D.n7307 D.t1193 7.599
R12469 D.n7293 D.t2785 7.599
R12470 D.n7279 D.t1171 7.599
R12471 D.n7265 D.t600 7.599
R12472 D.n7251 D.t779 7.599
R12473 D.n7237 D.t642 7.599
R12474 D.n7387 D.t2277 7.599
R12475 D.n7403 D.t3724 7.599
R12476 D.n7515 D.t1294 7.599
R12477 D.n7501 D.t3979 7.599
R12478 D.n7487 D.t568 7.599
R12479 D.n7473 D.t1190 7.599
R12480 D.n7459 D.t1455 7.599
R12481 D.n7445 D.t4363 7.599
R12482 D.n7431 D.t3 7.599
R12483 D.n7417 D.t3733 7.599
R12484 D.n7539 D.t3151 7.599
R12485 D.n7555 D.t1414 7.599
R12486 D.n7639 D.t1693 7.599
R12487 D.n7625 D.t2235 7.599
R12488 D.n7611 D.t2838 7.599
R12489 D.n7597 D.t3868 7.599
R12490 D.n7583 D.t1449 7.599
R12491 D.n7569 D.t3291 7.599
R12492 D.n7663 D.t376 7.599
R12493 D.n7679 D.t3015 7.599
R12494 D.n7735 D.t16 7.599
R12495 D.n7721 D.t592 7.599
R12496 D.n7707 D.t3900 7.599
R12497 D.n7693 D.t3749 7.599
R12498 D.n7758 D.t984 7.599
R12499 D.n7774 D.t309 7.599
R12500 D.n7802 D.t2017 7.599
R12501 D.n7788 D.t3545 7.599
R12502 D.n7839 D.t3587 7.493
R12503 D.n7829 D.t747 7.493
R12504 D.n450 D.t3952 7.493
R12505 D.n441 D.t2441 7.493
R12506 D.n32 D.t2632 7.493
R12507 D.n7892 D.t2343 7.493
R12508 D.n7976 D.t268 7.493
R12509 D.n7959 D.t3782 7.493
R12510 D.n7944 D.t3468 7.493
R12511 D.n14064 D.t4253 7.493
R12512 D.n14046 D.t2824 7.493
R12513 D.n14028 D.t3908 7.493
R12514 D.n14010 D.t4208 7.493
R12515 D.n13992 D.t3016 7.493
R12516 D.n13974 D.t1916 7.493
R12517 D.n13956 D.t1388 7.493
R12518 D.n13938 D.t4495 7.493
R12519 D.n13920 D.t2100 7.493
R12520 D.n13902 D.t476 7.493
R12521 D.n13884 D.t2497 7.493
R12522 D.n13866 D.t3089 7.493
R12523 D.n13848 D.t3763 7.493
R12524 D.n13830 D.t2247 7.493
R12525 D.n13812 D.t3781 7.493
R12526 D.n13794 D.t3120 7.493
R12527 D.n13776 D.t2536 7.493
R12528 D.n13758 D.t2730 7.493
R12529 D.n13740 D.t4246 7.493
R12530 D.n13722 D.t2967 7.493
R12531 D.n13704 D.t93 7.493
R12532 D.n13685 D.t1112 7.493
R12533 D.n13659 D.t2526 7.493
R12534 D.n13695 D.t2979 7.493
R12535 D.n13713 D.t361 7.493
R12536 D.n13731 D.t2462 7.493
R12537 D.n13749 D.t2938 7.493
R12538 D.n13767 D.t831 7.493
R12539 D.n13785 D.t1236 7.493
R12540 D.n13803 D.t1605 7.493
R12541 D.n13821 D.t3282 7.493
R12542 D.n13839 D.t4144 7.493
R12543 D.n13857 D.t1837 7.493
R12544 D.n13875 D.t3577 7.493
R12545 D.n13893 D.t4342 7.493
R12546 D.n13911 D.t949 7.493
R12547 D.n13929 D.t508 7.493
R12548 D.n13947 D.t3514 7.493
R12549 D.n13965 D.t3670 7.493
R12550 D.n13983 D.t3613 7.493
R12551 D.n14001 D.t3386 7.493
R12552 D.n14019 D.t3100 7.493
R12553 D.n14037 D.t2104 7.493
R12554 D.n14055 D.t1720 7.493
R12555 D.n14077 D.t2275 7.493
R12556 D.n13210 D.t3336 7.493
R12557 D.n13230 D.t694 7.493
R12558 D.n13250 D.t2504 7.493
R12559 D.n13270 D.t2397 7.493
R12560 D.n13290 D.t2585 7.493
R12561 D.n13310 D.t2580 7.493
R12562 D.n13330 D.t581 7.493
R12563 D.n13350 D.t2920 7.493
R12564 D.n13370 D.t2844 7.493
R12565 D.n13390 D.t474 7.493
R12566 D.n13410 D.t2139 7.493
R12567 D.n13430 D.t3549 7.493
R12568 D.n13450 D.t2152 7.493
R12569 D.n13470 D.t564 7.493
R12570 D.n13490 D.t1259 7.493
R12571 D.n13510 D.t1329 7.493
R12572 D.n13530 D.t2599 7.493
R12573 D.n13550 D.t3998 7.493
R12574 D.n13570 D.t3144 7.493
R12575 D.n13590 D.t3705 7.493
R12576 D.n13610 D.t2625 7.493
R12577 D.n13624 D.t693 7.493
R12578 D.n13599 D.t334 7.493
R12579 D.n13579 D.t2077 7.493
R12580 D.n13559 D.t394 7.493
R12581 D.n13539 D.t2452 7.493
R12582 D.n13519 D.t1018 7.493
R12583 D.n13499 D.t3509 7.493
R12584 D.n13479 D.t2918 7.493
R12585 D.n13459 D.t782 7.493
R12586 D.n13439 D.t1972 7.493
R12587 D.n13419 D.t3761 7.493
R12588 D.n13399 D.t2966 7.493
R12589 D.n13379 D.t517 7.493
R12590 D.n13359 D.t1058 7.493
R12591 D.n13339 D.t1089 7.493
R12592 D.n13319 D.t3861 7.493
R12593 D.n13299 D.t2646 7.493
R12594 D.n13279 D.t1845 7.493
R12595 D.n13259 D.t980 7.493
R12596 D.n13239 D.t2131 7.493
R12597 D.n13219 D.t4008 7.493
R12598 D.n13194 D.t1494 7.493
R12599 D.n13101 D.t3057 7.493
R12600 D.n13083 D.t1882 7.493
R12601 D.n13065 D.t4461 7.493
R12602 D.n13047 D.t4511 7.493
R12603 D.n13029 D.t3074 7.493
R12604 D.n13011 D.t1512 7.493
R12605 D.n12993 D.t2117 7.493
R12606 D.n12975 D.t2357 7.493
R12607 D.n12957 D.t2607 7.493
R12608 D.n12939 D.t4036 7.493
R12609 D.n12921 D.t510 7.493
R12610 D.n12903 D.t804 7.493
R12611 D.n12885 D.t4290 7.493
R12612 D.n12867 D.t2106 7.493
R12613 D.n12849 D.t1334 7.493
R12614 D.n12831 D.t1110 7.493
R12615 D.n12813 D.t844 7.493
R12616 D.n12795 D.t3755 7.493
R12617 D.n12777 D.t3551 7.493
R12618 D.n12758 D.t2766 7.493
R12619 D.n12736 D.t3498 7.493
R12620 D.n12768 D.t1657 7.493
R12621 D.n12786 D.t1206 7.493
R12622 D.n12804 D.t302 7.493
R12623 D.n12822 D.t90 7.493
R12624 D.n12840 D.t3451 7.493
R12625 D.n12858 D.t3681 7.493
R12626 D.n12876 D.t3758 7.493
R12627 D.n12894 D.t1782 7.493
R12628 D.n12912 D.t4057 7.493
R12629 D.n12930 D.t4148 7.493
R12630 D.n12948 D.t1697 7.493
R12631 D.n12966 D.t415 7.493
R12632 D.n12984 D.t3510 7.493
R12633 D.n13002 D.t3642 7.493
R12634 D.n13020 D.t3569 7.493
R12635 D.n13038 D.t4210 7.493
R12636 D.n13056 D.t4409 7.493
R12637 D.n13074 D.t4450 7.493
R12638 D.n13092 D.t4033 7.493
R12639 D.n13113 D.t1763 7.493
R12640 D.n12327 D.t1777 7.493
R12641 D.n12347 D.t1364 7.493
R12642 D.n12367 D.t1727 7.493
R12643 D.n12387 D.t3091 7.493
R12644 D.n12407 D.t907 7.493
R12645 D.n12427 D.t4021 7.493
R12646 D.n12447 D.t2187 7.493
R12647 D.n12467 D.t4486 7.493
R12648 D.n12487 D.t1589 7.493
R12649 D.n12507 D.t4339 7.493
R12650 D.n12527 D.t2309 7.493
R12651 D.n12547 D.t1809 7.493
R12652 D.n12567 D.t3523 7.493
R12653 D.n12587 D.t2177 7.493
R12654 D.n12607 D.t2644 7.493
R12655 D.n12627 D.t1520 7.493
R12656 D.n12647 D.t3629 7.493
R12657 D.n12667 D.t4165 7.493
R12658 D.n12687 D.t2256 7.493
R12659 D.n12701 D.t2168 7.493
R12660 D.n12676 D.t1075 7.493
R12661 D.n12656 D.t1005 7.493
R12662 D.n12636 D.t757 7.493
R12663 D.n12616 D.t2988 7.493
R12664 D.n12596 D.t1735 7.493
R12665 D.n12576 D.t2032 7.493
R12666 D.n12556 D.t1184 7.493
R12667 D.n12536 D.t4190 7.493
R12668 D.n12516 D.t3948 7.493
R12669 D.n12496 D.t936 7.493
R12670 D.n12476 D.t572 7.493
R12671 D.n12456 D.t3400 7.493
R12672 D.n12436 D.t3682 7.493
R12673 D.n12416 D.t3365 7.493
R12674 D.n12396 D.t3370 7.493
R12675 D.n12376 D.t3417 7.493
R12676 D.n12356 D.t3881 7.493
R12677 D.n12336 D.t2591 7.493
R12678 D.n12311 D.t4289 7.493
R12679 D.n12216 D.t2527 7.493
R12680 D.n12198 D.t1952 7.493
R12681 D.n12180 D.t2137 7.493
R12682 D.n12162 D.t4344 7.493
R12683 D.n12144 D.t3084 7.493
R12684 D.n12126 D.t677 7.493
R12685 D.n12108 D.t724 7.493
R12686 D.n12090 D.t2828 7.493
R12687 D.n12072 D.t3143 7.493
R12688 D.n12054 D.t1699 7.493
R12689 D.n12036 D.t98 7.493
R12690 D.n12018 D.t687 7.493
R12691 D.n12000 D.t1393 7.493
R12692 D.n11982 D.t589 7.493
R12693 D.n11964 D.t2199 7.493
R12694 D.n11946 D.t1778 7.493
R12695 D.n11928 D.t224 7.493
R12696 D.n11909 D.t3938 7.493
R12697 D.n11887 D.t20 7.493
R12698 D.n11919 D.t2079 7.493
R12699 D.n11937 D.t3594 7.493
R12700 D.n11955 D.t3477 7.493
R12701 D.n11973 D.t821 7.493
R12702 D.n11991 D.t1054 7.493
R12703 D.n12009 D.t4262 7.493
R12704 D.n12027 D.t2916 7.493
R12705 D.n12045 D.t2479 7.493
R12706 D.n12063 D.t2466 7.493
R12707 D.n12081 D.t1244 7.493
R12708 D.n12099 D.t1199 7.493
R12709 D.n12117 D.t3500 7.493
R12710 D.n12135 D.t2034 7.493
R12711 D.n12153 D.t1155 7.493
R12712 D.n12171 D.t852 7.493
R12713 D.n12189 D.t444 7.493
R12714 D.n12207 D.t1263 7.493
R12715 D.n12229 D.t895 7.493
R12716 D.n11518 D.t2037 7.493
R12717 D.n11538 D.t4032 7.493
R12718 D.n11558 D.t2288 7.493
R12719 D.n11578 D.t2440 7.493
R12720 D.n11598 D.t3274 7.493
R12721 D.n11618 D.t1117 7.493
R12722 D.n11638 D.t2109 7.493
R12723 D.n11658 D.t1335 7.493
R12724 D.n11678 D.t2038 7.493
R12725 D.n11698 D.t3748 7.493
R12726 D.n11718 D.t134 7.493
R12727 D.n11738 D.t532 7.493
R12728 D.n11758 D.t377 7.493
R12729 D.n11778 D.t740 7.493
R12730 D.n11798 D.t4090 7.493
R12731 D.n11818 D.t26 7.493
R12732 D.n11838 D.t539 7.493
R12733 D.n11852 D.t4371 7.493
R12734 D.n11827 D.t2874 7.493
R12735 D.n11807 D.t998 7.493
R12736 D.n11787 D.t3195 7.493
R12737 D.n11767 D.t1549 7.493
R12738 D.n11747 D.t4260 7.493
R12739 D.n11727 D.t3833 7.493
R12740 D.n11707 D.t2112 7.493
R12741 D.n11687 D.t1502 7.493
R12742 D.n11667 D.t2699 7.493
R12743 D.n11647 D.t3455 7.493
R12744 D.n11627 D.t3588 7.493
R12745 D.n11607 D.t4095 7.493
R12746 D.n11587 D.t4223 7.493
R12747 D.n11567 D.t4157 7.493
R12748 D.n11547 D.t3739 7.493
R12749 D.n11527 D.t4252 7.493
R12750 D.n11504 D.t2293 7.493
R12751 D.n11417 D.t4130 7.493
R12752 D.n11399 D.t2174 7.493
R12753 D.n11381 D.t4475 7.493
R12754 D.n11363 D.t2713 7.493
R12755 D.n11345 D.t628 7.493
R12756 D.n11327 D.t4013 7.493
R12757 D.n11309 D.t2178 7.493
R12758 D.n11291 D.t4254 7.493
R12759 D.n11273 D.t4054 7.493
R12760 D.n11255 D.t2977 7.493
R12761 D.n11237 D.t698 7.493
R12762 D.n11219 D.t3837 7.493
R12763 D.n11201 D.t1577 7.493
R12764 D.n11183 D.t2589 7.493
R12765 D.n11165 D.t3909 7.493
R12766 D.n11146 D.t3579 7.493
R12767 D.n11124 D.t1454 7.493
R12768 D.n11156 D.t1712 7.493
R12769 D.n11174 D.t4063 7.493
R12770 D.n11192 D.t3704 7.493
R12771 D.n11210 D.t3087 7.493
R12772 D.n11228 D.t2500 7.493
R12773 D.n11246 D.t477 7.493
R12774 D.n11264 D.t3746 7.493
R12775 D.n11282 D.t2087 7.493
R12776 D.n11300 D.t2336 7.493
R12777 D.n11318 D.t4140 7.493
R12778 D.n11336 D.t3925 7.493
R12779 D.n11354 D.t3716 7.493
R12780 D.n11372 D.t3943 7.493
R12781 D.n11390 D.t3973 7.493
R12782 D.n11408 D.t551 7.493
R12783 D.n11430 D.t4330 7.493
R12784 D.n10795 D.t3218 7.493
R12785 D.n10815 D.t1390 7.493
R12786 D.n10835 D.t1668 7.493
R12787 D.n10855 D.t2912 7.493
R12788 D.n10875 D.t3005 7.493
R12789 D.n10895 D.t1394 7.493
R12790 D.n10915 D.t910 7.493
R12791 D.n10935 D.t431 7.493
R12792 D.n10955 D.t1428 7.493
R12793 D.n10975 D.t1725 7.493
R12794 D.n10995 D.t3114 7.493
R12795 D.n11015 D.t759 7.493
R12796 D.n11035 D.t396 7.493
R12797 D.n11055 D.t1432 7.493
R12798 D.n11075 D.t3366 7.493
R12799 D.n11089 D.t1146 7.493
R12800 D.n11064 D.t2042 7.493
R12801 D.n11044 D.t4214 7.493
R12802 D.n11024 D.t3550 7.493
R12803 D.n11004 D.t2140 7.493
R12804 D.n10984 D.t1198 7.493
R12805 D.n10964 D.t696 7.493
R12806 D.n10944 D.t1430 7.493
R12807 D.n10924 D.t3877 7.493
R12808 D.n10904 D.t1105 7.493
R12809 D.n10884 D.t2007 7.493
R12810 D.n10864 D.t1144 7.493
R12811 D.n10844 D.t2227 7.493
R12812 D.n10824 D.t339 7.493
R12813 D.n10804 D.t1169 7.493
R12814 D.n10781 D.t2446 7.493
R12815 D.n10698 D.t3951 7.493
R12816 D.n10680 D.t2089 7.493
R12817 D.n10662 D.t2272 7.493
R12818 D.n10644 D.t2398 7.493
R12819 D.n10626 D.t2587 7.493
R12820 D.n10608 D.t135 7.493
R12821 D.n10590 D.t4073 7.493
R12822 D.n10572 D.t976 7.493
R12823 D.n10554 D.t1621 7.493
R12824 D.n10536 D.t289 7.493
R12825 D.n10518 D.t916 7.493
R12826 D.n10500 D.t2999 7.493
R12827 D.n10482 D.t2750 7.493
R12828 D.n10463 D.t1703 7.493
R12829 D.n10441 D.t4331 7.493
R12830 D.n10473 D.t4334 7.493
R12831 D.n10491 D.t1228 7.493
R12832 D.n10509 D.t511 7.493
R12833 D.n10527 D.t4037 7.493
R12834 D.n10545 D.t1355 7.493
R12835 D.n10563 D.t2694 7.493
R12836 D.n10581 D.t3288 7.493
R12837 D.n10599 D.t1049 7.493
R12838 D.n10617 D.t2686 7.493
R12839 D.n10635 D.t4329 7.493
R12840 D.n10653 D.t3854 7.493
R12841 D.n10671 D.t4429 7.493
R12842 D.n10689 D.t4298 7.493
R12843 D.n10711 D.t4279 7.493
R12844 D.n10152 D.t1359 7.493
R12845 D.n10172 D.t2160 7.493
R12846 D.n10192 D.t4464 7.493
R12847 D.n10212 D.t490 7.493
R12848 D.n10232 D.t3768 7.493
R12849 D.n10252 D.t4296 7.493
R12850 D.n10272 D.t4449 7.493
R12851 D.n10292 D.t4250 7.493
R12852 D.n10312 D.t1037 7.493
R12853 D.n10332 D.t1251 7.493
R12854 D.n10352 D.t1998 7.493
R12855 D.n10372 D.t3167 7.493
R12856 D.n10392 D.t2995 7.493
R12857 D.n10406 D.t3540 7.493
R12858 D.n10381 D.t2285 7.493
R12859 D.n10361 D.t2076 7.493
R12860 D.n10341 D.t4271 7.493
R12861 D.n10321 D.t4458 7.493
R12862 D.n10301 D.t2643 7.493
R12863 D.n10281 D.t3031 7.493
R12864 D.n10261 D.t2863 7.493
R12865 D.n10241 D.t3135 7.493
R12866 D.n10221 D.t2850 7.493
R12867 D.n10201 D.t3820 7.493
R12868 D.n10181 D.t3257 7.493
R12869 D.n10161 D.t1871 7.493
R12870 D.n10136 D.t1156 7.493
R12871 D.n10059 D.t340 7.493
R12872 D.n10041 D.t1594 7.493
R12873 D.n10023 D.t1730 7.493
R12874 D.n10005 D.t481 7.493
R12875 D.n9987 D.t3590 7.493
R12876 D.n9969 D.t2295 7.493
R12877 D.n9951 D.t925 7.493
R12878 D.n9933 D.t3655 7.493
R12879 D.n9915 D.t4215 7.493
R12880 D.n9897 D.t1029 7.493
R12881 D.n9879 D.t1658 7.493
R12882 D.n9860 D.t3974 7.493
R12883 D.n9838 D.t286 7.493
R12884 D.n9870 D.t2170 7.493
R12885 D.n9888 D.t84 7.493
R12886 D.n9906 D.t1652 7.493
R12887 D.n9924 D.t1301 7.493
R12888 D.n9942 D.t3552 7.493
R12889 D.n9960 D.t1093 7.493
R12890 D.n9978 D.t1888 7.493
R12891 D.n9996 D.t2420 7.493
R12892 D.n10014 D.t2252 7.493
R12893 D.n10032 D.t1949 7.493
R12894 D.n10050 D.t876 7.493
R12895 D.n10071 D.t3152 7.493
R12896 D.n9589 D.t3759 7.493
R12897 D.n9609 D.t2029 7.493
R12898 D.n9629 D.t261 7.493
R12899 D.n9649 D.t1718 7.493
R12900 D.n9669 D.t1026 7.493
R12901 D.n9689 D.t1953 7.493
R12902 D.n9709 D.t781 7.493
R12903 D.n9729 D.t1627 7.493
R12904 D.n9749 D.t1472 7.493
R12905 D.n9769 D.t2681 7.493
R12906 D.n9789 D.t1180 7.493
R12907 D.n9803 D.t3265 7.493
R12908 D.n9778 D.t1914 7.493
R12909 D.n9758 D.t2122 7.493
R12910 D.n9738 D.t1887 7.493
R12911 D.n9718 D.t3562 7.493
R12912 D.n9698 D.t258 7.493
R12913 D.n9678 D.t1734 7.493
R12914 D.n9658 D.t2602 7.493
R12915 D.n9638 D.t164 7.493
R12916 D.n9618 D.t1939 7.493
R12917 D.n9598 D.t4185 7.493
R12918 D.n9573 D.t1797 7.493
R12919 D.n9494 D.t2439 7.493
R12920 D.n9476 D.t4268 7.493
R12921 D.n9458 D.t3233 7.493
R12922 D.n9440 D.t4419 7.493
R12923 D.n9422 D.t3586 7.493
R12924 D.n9404 D.t3197 7.493
R12925 D.n9386 D.t3793 7.493
R12926 D.n9368 D.t1509 7.493
R12927 D.n9350 D.t112 7.493
R12928 D.n9331 D.t2972 7.493
R12929 D.n9309 D.t1462 7.493
R12930 D.n9341 D.t2732 7.493
R12931 D.n9359 D.t2711 7.493
R12932 D.n9377 D.t2770 7.493
R12933 D.n9395 D.t2733 7.493
R12934 D.n9413 D.t3045 7.493
R12935 D.n9431 D.t3062 7.493
R12936 D.n9449 D.t3132 7.493
R12937 D.n9467 D.t2808 7.493
R12938 D.n9485 D.t2840 7.493
R12939 D.n9507 D.t3372 7.493
R12940 D.n9100 D.t4438 7.493
R12941 D.n9120 D.t871 7.493
R12942 D.n9140 D.t1877 7.493
R12943 D.n9160 D.t463 7.493
R12944 D.n9180 D.t3444 7.493
R12945 D.n9200 D.t4357 7.493
R12946 D.n9220 D.t4065 7.493
R12947 D.n9240 D.t4403 7.493
R12948 D.n9260 D.t3491 7.493
R12949 D.n9274 D.t226 7.493
R12950 D.n9249 D.t525 7.493
R12951 D.n9229 D.t3803 7.493
R12952 D.n9209 D.t1081 7.493
R12953 D.n9189 D.t499 7.493
R12954 D.n9169 D.t2411 7.493
R12955 D.n9149 D.t2213 7.493
R12956 D.n9129 D.t3225 7.493
R12957 D.n9109 D.t386 7.493
R12958 D.n9086 D.t528 7.493
R12959 D.n9015 D.t1866 7.493
R12960 D.n8997 D.t2456 7.493
R12961 D.n8979 D.t3662 7.493
R12962 D.n8961 D.t1438 7.493
R12963 D.n8943 D.t3249 7.493
R12964 D.n8925 D.t3374 7.493
R12965 D.n8907 D.t343 7.493
R12966 D.n8888 D.t2291 7.493
R12967 D.n8866 D.t2807 7.493
R12968 D.n8898 D.t3414 7.493
R12969 D.n8916 D.t45 7.493
R12970 D.n8934 D.t2041 7.493
R12971 D.n8952 D.t1317 7.493
R12972 D.n8970 D.t36 7.493
R12973 D.n8988 D.t623 7.493
R12974 D.n9006 D.t1716 7.493
R12975 D.n9028 D.t4183 7.493
R12976 D.n8697 D.t2882 7.493
R12977 D.n8717 D.t4326 7.493
R12978 D.n8737 D.t573 7.493
R12979 D.n8757 D.t1932 7.493
R12980 D.n8777 D.t1010 7.493
R12981 D.n8797 D.t450 7.493
R12982 D.n8817 D.t3796 7.493
R12983 D.n8831 D.t2324 7.493
R12984 D.n8806 D.t2980 7.493
R12985 D.n8786 D.t2946 7.493
R12986 D.n8766 D.t2974 7.493
R12987 D.n8746 D.t3029 7.493
R12988 D.n8726 D.t2775 7.493
R12989 D.n8706 D.t2767 7.493
R12990 D.n8681 D.t92 7.493
R12991 D.n8616 D.t128 7.493
R12992 D.n8598 D.t4413 7.493
R12993 D.n8580 D.t3276 7.493
R12994 D.n8562 D.t3703 7.493
R12995 D.n8544 D.t4444 7.493
R12996 D.n8525 D.t1447 7.493
R12997 D.n8503 D.t4502 7.493
R12998 D.n8535 D.t161 7.493
R12999 D.n8553 D.t2393 7.493
R13000 D.n8571 D.t1962 7.493
R13001 D.n8589 D.t3826 7.493
R13002 D.n8607 D.t2605 7.493
R13003 D.n8628 D.t2884 7.493
R13004 D.n8374 D.t2331 7.493
R13005 D.n8394 D.t1218 7.493
R13006 D.n8414 D.t3192 7.493
R13007 D.n8434 D.t1423 7.493
R13008 D.n8454 D.t1053 7.493
R13009 D.n8468 D.t549 7.493
R13010 D.n8443 D.t685 7.493
R13011 D.n8423 D.t3193 7.493
R13012 D.n8403 D.t882 7.493
R13013 D.n8383 D.t2130 7.493
R13014 D.n8358 D.t3520 7.493
R13015 D.n8291 D.t3075 7.493
R13016 D.n8273 D.t3263 7.493
R13017 D.n8255 D.t1278 7.493
R13018 D.n8236 D.t4267 7.493
R13019 D.n8214 D.t1823 7.493
R13020 D.n8246 D.t3122 7.493
R13021 D.n8264 D.t3054 7.493
R13022 D.n8282 D.t4163 7.493
R13023 D.n8304 D.t4151 7.493
R13024 D.n8125 D.t2455 7.493
R13025 D.n8145 D.t4295 7.493
R13026 D.n8165 D.t2496 7.493
R13027 D.n8179 D.t2538 7.493
R13028 D.n8154 D.t3811 7.493
R13029 D.n8134 D.t2092 7.493
R13030 D.n8111 D.t2724 7.493
R13031 D.n8052 D.t3042 7.493
R13032 D.n8033 D.t1170 7.493
R13033 D.n8011 D.t1343 7.493
R13034 D.n8043 D.t1157 7.493
R13035 D.n8065 D.t1878 7.493
R13036 D.n54 D.t179 7.493
R13037 D.n63 D.t3983 7.493
R13038 D.n72 D.t705 7.493
R13039 D.n81 D.t414 7.493
R13040 D.n90 D.t2885 7.493
R13041 D.n99 D.t254 7.493
R13042 D.n108 D.t3883 7.493
R13043 D.n117 D.t4319 7.493
R13044 D.n126 D.t2954 7.493
R13045 D.n135 D.t1586 7.493
R13046 D.n144 D.t951 7.493
R13047 D.n153 D.t1518 7.493
R13048 D.n162 D.t1632 7.493
R13049 D.n171 D.t2896 7.493
R13050 D.n180 D.t1340 7.493
R13051 D.n189 D.t3110 7.493
R13052 D.n198 D.t3354 7.493
R13053 D.n207 D.t2044 7.493
R13054 D.n216 D.t238 7.493
R13055 D.n225 D.t2762 7.493
R13056 D.n234 D.t661 7.493
R13057 D.n243 D.t4264 7.493
R13058 D.n252 D.t1561 7.493
R13059 D.n261 D.t3831 7.493
R13060 D.n270 D.t3641 7.493
R13061 D.n279 D.t2110 7.493
R13062 D.n288 D.t47 7.493
R13063 D.n297 D.t2318 7.493
R13064 D.n306 D.t3887 7.493
R13065 D.n315 D.t4474 7.493
R13066 D.n324 D.t1044 7.493
R13067 D.n333 D.t2172 7.493
R13068 D.n342 D.t3964 7.493
R13069 D.n351 D.t4006 7.493
R13070 D.n360 D.t4098 7.493
R13071 D.n369 D.t411 7.493
R13072 D.n378 D.t2707 7.493
R13073 D.n387 D.t2084 7.493
R13074 D.n396 D.t2894 7.493
R13075 D.n405 D.t1754 7.493
R13076 D.n414 D.t721 7.493
R13077 D.n423 D.t1485 7.493
R13078 D.n432 D.t274 7.493
R13079 D.n526 D.t4016 7.493
R13080 D.n542 D.t2465 7.493
R13081 D.n1130 D.t2555 7.493
R13082 D.n1116 D.t616 7.493
R13083 D.n1102 D.t2952 7.493
R13084 D.n1088 D.t3959 7.493
R13085 D.n1074 D.t3189 7.493
R13086 D.n1060 D.t4211 7.493
R13087 D.n1046 D.t2638 7.493
R13088 D.n1032 D.t556 7.493
R13089 D.n1018 D.t1785 7.493
R13090 D.n1004 D.t775 7.493
R13091 D.n990 D.t1807 7.493
R13092 D.n976 D.t3044 7.493
R13093 D.n962 D.t1231 7.493
R13094 D.n948 D.t1123 7.493
R13095 D.n934 D.t2060 7.493
R13096 D.n920 D.t2210 7.493
R13097 D.n906 D.t3610 7.493
R13098 D.n892 D.t701 7.493
R13099 D.n878 D.t820 7.493
R13100 D.n864 D.t2780 7.493
R13101 D.n850 D.t1055 7.493
R13102 D.n836 D.t3279 7.493
R13103 D.n822 D.t4307 7.493
R13104 D.n808 D.t1293 7.493
R13105 D.n794 D.t2768 7.493
R13106 D.n780 D.t168 7.493
R13107 D.n766 D.t2478 7.493
R13108 D.n752 D.t1583 7.493
R13109 D.n738 D.t2442 7.493
R13110 D.n724 D.t1608 7.493
R13111 D.n710 D.t2287 7.493
R13112 D.n696 D.t1805 7.493
R13113 D.n682 D.t2102 7.493
R13114 D.n668 D.t3474 7.493
R13115 D.n654 D.t1478 7.493
R13116 D.n640 D.t819 7.493
R13117 D.n626 D.t926 7.493
R13118 D.n612 D.t2114 7.493
R13119 D.n598 D.t2514 7.493
R13120 D.n584 D.t4482 7.493
R13121 D.n570 D.t197 7.493
R13122 D.n556 D.t2184 7.493
R13123 D.n1153 D.t2115 7.493
R13124 D.n1169 D.t990 7.493
R13125 D.n1729 D.t67 7.493
R13126 D.n1715 D.t963 7.493
R13127 D.n1701 D.t2962 7.493
R13128 D.n1687 D.t121 7.493
R13129 D.n1673 D.t4050 7.493
R13130 D.n1659 D.t51 7.493
R13131 D.n1645 D.t783 7.493
R13132 D.n1631 D.t3694 7.493
R13133 D.n1617 D.t1976 7.493
R13134 D.n1603 D.t3506 7.493
R13135 D.n1589 D.t3256 7.493
R13136 D.n1575 D.t2881 7.493
R13137 D.n1561 D.t235 7.493
R13138 D.n1547 D.t364 7.493
R13139 D.n1533 D.t3907 7.493
R13140 D.n1519 D.t596 7.493
R13141 D.n1505 D.t2839 7.493
R13142 D.n1491 D.t126 7.493
R13143 D.n1477 D.t2003 7.493
R13144 D.n1463 D.t3470 7.493
R13145 D.n1449 D.t2031 7.493
R13146 D.n1435 D.t505 7.493
R13147 D.n1421 D.t1637 7.493
R13148 D.n1407 D.t2419 7.493
R13149 D.n1393 D.t4191 7.493
R13150 D.n1379 D.t1232 7.493
R13151 D.n1365 D.t1732 7.493
R13152 D.n1351 D.t948 7.493
R13153 D.n1337 D.t4386 7.493
R13154 D.n1323 D.t1721 7.493
R13155 D.n1309 D.t2914 7.493
R13156 D.n1295 D.t1418 7.493
R13157 D.n1281 D.t4043 7.493
R13158 D.n1267 D.t3137 7.493
R13159 D.n1253 D.t3521 7.493
R13160 D.n1239 D.t3271 7.493
R13161 D.n1225 D.t4420 7.493
R13162 D.n1211 D.t2221 7.493
R13163 D.n1197 D.t4244 7.493
R13164 D.n1183 D.t2347 7.493
R13165 D.n1752 D.t2973 7.493
R13166 D.n1768 D.t346 7.493
R13167 D.n2300 D.t1014 7.493
R13168 D.n2286 D.t1855 7.493
R13169 D.n2272 D.t3512 7.493
R13170 D.n2258 D.t144 7.493
R13171 D.n2244 D.t4184 7.493
R13172 D.n2230 D.t170 7.493
R13173 D.n2216 D.t4146 7.493
R13174 D.n2202 D.t3932 7.493
R13175 D.n2188 D.t325 7.493
R13176 D.n2174 D.t3633 7.493
R13177 D.n2160 D.t720 7.493
R13178 D.n2146 D.t710 7.493
R13179 D.n2132 D.t1132 7.493
R13180 D.n2118 D.t276 7.493
R13181 D.n2104 D.t4476 7.493
R13182 D.n2090 D.t373 7.493
R13183 D.n2076 D.t4454 7.493
R13184 D.n2062 D.t99 7.493
R13185 D.n2048 D.t3680 7.493
R13186 D.n2034 D.t48 7.493
R13187 D.n2020 D.t3756 7.493
R13188 D.n2006 D.t2900 7.493
R13189 D.n1992 D.t1779 7.493
R13190 D.n1978 D.t1477 7.493
R13191 D.n1964 D.t2695 7.493
R13192 D.n1950 D.t840 7.493
R13193 D.n1936 D.t2242 7.493
R13194 D.n1922 D.t59 7.493
R13195 D.n1908 D.t2097 7.493
R13196 D.n1894 D.t3894 7.493
R13197 D.n1880 D.t307 7.493
R13198 D.n1866 D.t2735 7.493
R13199 D.n1852 D.t2286 7.493
R13200 D.n1838 D.t3036 7.493
R13201 D.n1824 D.t131 7.493
R13202 D.n1810 D.t2970 7.493
R13203 D.n1796 D.t3639 7.493
R13204 D.n1782 D.t4387 7.493
R13205 D.n2323 D.t1708 7.493
R13206 D.n2339 D.t885 7.493
R13207 D.n2843 D.t1545 7.493
R13208 D.n2829 D.t402 7.493
R13209 D.n2815 D.t1036 7.493
R13210 D.n2801 D.t3823 7.493
R13211 D.n2787 D.t3229 7.493
R13212 D.n2773 D.t77 7.493
R13213 D.n2759 D.t3139 7.493
R13214 D.n2745 D.t4481 7.493
R13215 D.n2731 D.t884 7.493
R13216 D.n2717 D.t957 7.493
R13217 D.n2703 D.t3865 7.493
R13218 D.n2689 D.t2181 7.493
R13219 D.n2675 D.t2426 7.493
R13220 D.n2661 D.t3264 7.493
R13221 D.n2647 D.t32 7.493
R13222 D.n2633 D.t1810 7.493
R13223 D.n2619 D.t3352 7.493
R13224 D.n2605 D.t2313 7.493
R13225 D.n2591 D.t2936 7.493
R13226 D.n2577 D.t177 7.493
R13227 D.n2563 D.t780 7.493
R13228 D.n2549 D.t3869 7.493
R13229 D.n2535 D.t186 7.493
R13230 D.n2521 D.t664 7.493
R13231 D.n2507 D.t2085 7.493
R13232 D.n2493 D.t2370 7.493
R13233 D.n2479 D.t1313 7.493
R13234 D.n2465 D.t1556 7.493
R13235 D.n2451 D.t3375 7.493
R13236 D.n2437 D.t2422 7.493
R13237 D.n2423 D.t1260 7.493
R13238 D.n2409 D.t1312 7.493
R13239 D.n2395 D.t2476 7.493
R13240 D.n2381 D.t34 7.493
R13241 D.n2367 D.t1841 7.493
R13242 D.n2353 D.t1508 7.493
R13243 D.n2866 D.t3757 7.493
R13244 D.n2882 D.t504 7.493
R13245 D.n3358 D.t1601 7.493
R13246 D.n3344 D.t4356 7.493
R13247 D.n3330 D.t2211 7.493
R13248 D.n3316 D.t1554 7.493
R13249 D.n3302 D.t614 7.493
R13250 D.n3288 D.t2338 7.493
R13251 D.n3274 D.t4423 7.493
R13252 D.n3260 D.t320 7.493
R13253 D.n3246 D.t2617 7.493
R13254 D.n3232 D.t2345 7.493
R13255 D.n3218 D.t3103 7.493
R13256 D.n3204 D.t2601 7.493
R13257 D.n3190 D.t3409 7.493
R13258 D.n3176 D.t3852 7.493
R13259 D.n3162 D.t522 7.493
R13260 D.n3148 D.t1611 7.493
R13261 D.n3134 D.t1560 7.493
R13262 D.n3120 D.t3876 7.493
R13263 D.n3106 D.t4439 7.493
R13264 D.n3092 D.t70 7.493
R13265 D.n3078 D.t3011 7.493
R13266 D.n3064 D.t1382 7.493
R13267 D.n3050 D.t1240 7.493
R13268 D.n3036 D.t3002 7.493
R13269 D.n3022 D.t1625 7.493
R13270 D.n3008 D.t1440 7.493
R13271 D.n2994 D.t3928 7.493
R13272 D.n2980 D.t2959 7.493
R13273 D.n2966 D.t4349 7.493
R13274 D.n2952 D.t498 7.493
R13275 D.n2938 D.t4197 7.493
R13276 D.n2924 D.t2404 7.493
R13277 D.n2910 D.t3618 7.493
R13278 D.n2896 D.t2025 7.493
R13279 D.n3382 D.t2811 7.493
R13280 D.n3398 D.t2666 7.493
R13281 D.n3846 D.t808 7.493
R13282 D.n3832 D.t4281 7.493
R13283 D.n3818 D.t182 7.493
R13284 D.n3804 D.t207 7.493
R13285 D.n3790 D.t1947 7.493
R13286 D.n3776 D.t3807 7.493
R13287 D.n3762 D.t2942 7.493
R13288 D.n3748 D.t613 7.493
R13289 D.n3734 D.t3597 7.493
R13290 D.n3720 D.t868 7.493
R13291 D.n3706 D.t4309 7.493
R13292 D.n3692 D.t585 7.493
R13293 D.n3678 D.t3388 7.493
R13294 D.n3664 D.t2155 7.493
R13295 D.n3650 D.t2376 7.493
R13296 D.n3636 D.t4418 7.493
R13297 D.n3622 D.t1316 7.493
R13298 D.n3608 D.t1551 7.493
R13299 D.n3594 D.t109 7.493
R13300 D.n3580 D.t3525 7.493
R13301 D.n3566 D.t4345 7.493
R13302 D.n3552 D.t3205 7.493
R13303 D.n3538 D.t3237 7.493
R13304 D.n3524 D.t3853 7.493
R13305 D.n3510 D.t3220 7.493
R13306 D.n3496 D.t1740 7.493
R13307 D.n3482 D.t3056 7.493
R13308 D.n3468 D.t2949 7.493
R13309 D.n3454 D.t399 7.493
R13310 D.n3440 D.t2871 7.493
R13311 D.n3426 D.t178 7.493
R13312 D.n3412 D.t2817 7.493
R13313 D.n3870 D.t1620 7.493
R13314 D.n3886 D.t458 7.493
R13315 D.n4306 D.t3071 7.493
R13316 D.n4292 D.t4030 7.493
R13317 D.n4278 D.t3954 7.493
R13318 D.n4264 D.t4242 7.493
R13319 D.n4250 D.t148 7.493
R13320 D.n4236 D.t2484 7.493
R13321 D.n4222 D.t3332 7.493
R13322 D.n4208 D.t3472 7.493
R13323 D.n4194 D.t1524 7.493
R13324 D.n4180 D.t3719 7.493
R13325 D.n4166 D.t3602 7.493
R13326 D.n4152 D.t2261 7.493
R13327 D.n4138 D.t2854 7.493
R13328 D.n4124 D.t1437 7.493
R13329 D.n4110 D.t813 7.493
R13330 D.n4096 D.t4245 7.493
R13331 D.n4082 D.t3186 7.493
R13332 D.n4068 D.t2329 7.493
R13333 D.n4054 D.t1933 7.493
R13334 D.n4040 D.t3806 7.493
R13335 D.n4026 D.t1499 7.493
R13336 D.n4012 D.t1789 7.493
R13337 D.n3998 D.t1200 7.493
R13338 D.n3984 D.t201 7.493
R13339 D.n3970 D.t260 7.493
R13340 D.n3956 D.t1097 7.493
R13341 D.n3942 D.t4383 7.493
R13342 D.n3928 D.t265 7.493
R13343 D.n3914 D.t390 7.493
R13344 D.n3900 D.t1956 7.493
R13345 D.n4330 D.t1885 7.493
R13346 D.n4346 D.t4361 7.493
R13347 D.n4738 D.t4337 7.493
R13348 D.n4724 D.t375 7.493
R13349 D.n4710 D.t962 7.493
R13350 D.n4696 D.t4232 7.493
R13351 D.n4682 D.t101 7.493
R13352 D.n4668 D.t3557 7.493
R13353 D.n4654 D.t50 7.493
R13354 D.n4640 D.t2243 7.493
R13355 D.n4626 D.t2990 7.493
R13356 D.n4612 D.t3082 7.493
R13357 D.n4598 D.t2729 7.493
R13358 D.n4584 D.t2511 7.493
R13359 D.n4570 D.t4314 7.493
R13360 D.n4556 D.t2278 7.493
R13361 D.n4542 D.t2905 7.493
R13362 D.n4528 D.t4025 7.493
R13363 D.n4514 D.t3600 7.493
R13364 D.n4500 D.t4167 7.493
R13365 D.n4486 D.t1680 7.493
R13366 D.n4472 D.t4070 7.493
R13367 D.n4458 D.t533 7.493
R13368 D.n4444 D.t4121 7.493
R13369 D.n4430 D.t2413 7.493
R13370 D.n4416 D.t3980 7.493
R13371 D.n4402 D.t1669 7.493
R13372 D.n4388 D.t1271 7.493
R13373 D.n4374 D.t4134 7.493
R13374 D.n4360 D.t1092 7.493
R13375 D.n4762 D.t2993 7.493
R13376 D.n4778 D.t97 7.493
R13377 D.n5142 D.t3960 7.493
R13378 D.n5128 D.t3196 7.493
R13379 D.n5114 D.t1818 7.493
R13380 D.n5100 D.t3858 7.493
R13381 D.n5086 D.t2610 7.493
R13382 D.n5072 D.t1496 7.493
R13383 D.n5058 D.t171 7.493
R13384 D.n5044 D.t1408 7.493
R13385 D.n5030 D.t3429 7.493
R13386 D.n5016 D.t4291 7.493
R13387 D.n5002 D.t253 7.493
R13388 D.n4988 D.t3418 7.493
R13389 D.n4974 D.t1130 7.493
R13390 D.n4960 D.t2124 7.493
R13391 D.n4946 D.t4370 7.493
R13392 D.n4932 D.t2649 7.493
R13393 D.n4918 D.t1527 7.493
R13394 D.n4904 D.t4216 7.493
R13395 D.n4890 D.t1698 7.493
R13396 D.n4876 D.t1514 7.493
R13397 D.n4862 D.t2772 7.493
R13398 D.n4848 D.t2700 7.493
R13399 D.n4834 D.t1474 7.493
R13400 D.n4820 D.t2867 7.493
R13401 D.n4806 D.t3660 7.493
R13402 D.n4792 D.t452 7.493
R13403 D.n5166 D.t2778 7.493
R13404 D.n5182 D.t2363 7.493
R13405 D.n5518 D.t4220 7.493
R13406 D.n5504 D.t1993 7.493
R13407 D.n5490 D.t401 7.493
R13408 D.n5476 D.t1164 7.493
R13409 D.n5462 D.t3822 7.493
R13410 D.n5448 D.t2427 7.493
R13411 D.n5434 D.t71 7.493
R13412 D.n5420 D.t3398 7.493
R13413 D.n5406 D.t1687 7.493
R13414 D.n5392 D.t3767 7.493
R13415 D.n5378 D.t2024 7.493
R13416 D.n5364 D.t3004 7.493
R13417 D.n5350 D.t3442 7.493
R13418 D.n5336 D.t2490 7.493
R13419 D.n5322 D.t3331 7.493
R13420 D.n5308 D.t1943 7.493
R13421 D.n5294 D.t2308 7.493
R13422 D.n5280 D.t3697 7.493
R13423 D.n5266 D.t263 7.493
R13424 D.n5252 D.t2457 7.493
R13425 D.n5238 D.t4131 7.493
R13426 D.n5224 D.t1192 7.493
R13427 D.n5210 D.t1465 7.493
R13428 D.n5196 D.t2529 7.493
R13429 D.n5542 D.t1590 7.493
R13430 D.n5558 D.t2869 7.493
R13431 D.n5866 D.t2158 7.493
R13432 D.n5852 D.t3810 7.493
R13433 D.n5838 D.t3172 7.493
R13434 D.n5824 D.t586 7.493
R13435 D.n5810 D.t1553 7.493
R13436 D.n5796 D.t3321 7.493
R13437 D.n5782 D.t3702 7.493
R13438 D.n5768 D.t3117 7.493
R13439 D.n5754 D.t1792 7.493
R13440 D.n5740 D.t1548 7.493
R13441 D.n5726 D.t1628 7.493
R13442 D.n5712 D.t4064 7.493
R13443 D.n5698 D.t319 7.493
R13444 D.n5684 D.t3559 7.493
R13445 D.n5670 D.t3608 7.493
R13446 D.n5656 D.t3751 7.493
R13447 D.n5642 D.t3554 7.493
R13448 D.n5628 D.t2230 7.493
R13449 D.n5614 D.t8 7.493
R13450 D.n5600 D.t3345 7.493
R13451 D.n5586 D.t1375 7.493
R13452 D.n5572 D.t1559 7.493
R13453 D.n5890 D.t2035 7.493
R13454 D.n5906 D.t24 7.493
R13455 D.n6186 D.t1563 7.493
R13456 D.n6172 D.t909 7.493
R13457 D.n6158 D.t4322 7.493
R13458 D.n6144 D.t1959 7.493
R13459 D.n6130 D.t2330 7.493
R13460 D.n6116 D.t4508 7.493
R13461 D.n6102 D.t4071 7.493
R13462 D.n6088 D.t4412 7.493
R13463 D.n6074 D.t1580 7.493
R13464 D.n6060 D.t210 7.493
R13465 D.n6046 D.t3358 7.493
R13466 D.n6032 D.t3168 7.493
R13467 D.n6018 D.t755 7.493
R13468 D.n6004 D.t1970 7.493
R13469 D.n5990 D.t2684 7.493
R13470 D.n5976 D.t2086 7.493
R13471 D.n5962 D.t639 7.493
R13472 D.n5948 D.t3808 7.493
R13473 D.n5934 D.t3968 7.493
R13474 D.n5920 D.t543 7.493
R13475 D.n6210 D.t3801 7.493
R13476 D.n6226 D.t227 7.493
R13477 D.n6478 D.t491 7.493
R13478 D.n6464 D.t3380 7.493
R13479 D.n6450 D.t4026 7.493
R13480 D.n6436 D.t272 7.493
R13481 D.n6422 D.t4206 7.493
R13482 D.n6408 D.t1318 7.493
R13483 D.n6394 D.t1567 7.493
R13484 D.n6380 D.t2561 7.493
R13485 D.n6366 D.t23 7.493
R13486 D.n6352 D.t2009 7.493
R13487 D.n6338 D.t3207 7.493
R13488 D.n6324 D.t3302 7.493
R13489 D.n6310 D.t2740 7.493
R13490 D.n6296 D.t1241 7.493
R13491 D.n6282 D.t3428 7.493
R13492 D.n6268 D.t1675 7.493
R13493 D.n6254 D.t1930 7.493
R13494 D.n6240 D.t4492 7.493
R13495 D.n6502 D.t267 7.493
R13496 D.n6518 D.t3108 7.493
R13497 D.n6742 D.t2125 7.493
R13498 D.n6728 D.t3078 7.493
R13499 D.n6714 D.t1945 7.493
R13500 D.n6700 D.t897 7.493
R13501 D.n6686 D.t4009 7.493
R13502 D.n6672 D.t1151 7.493
R13503 D.n6658 D.t3176 7.493
R13504 D.n6644 D.t2670 7.493
R13505 D.n6630 D.t2748 7.493
R13506 D.n6616 D.t3298 7.493
R13507 D.n6602 D.t2424 7.493
R13508 D.n6588 D.t3947 7.493
R13509 D.n6574 D.t1023 7.493
R13510 D.n6560 D.t3238 7.493
R13511 D.n6546 D.t3350 7.493
R13512 D.n6532 D.t2312 7.493
R13513 D.n6766 D.t849 7.493
R13514 D.n6782 D.t2081 7.493
R13515 D.n6978 D.t3818 7.493
R13516 D.n6964 D.t4382 7.493
R13517 D.n6950 D.t2105 7.493
R13518 D.n6936 D.t3381 7.493
R13519 D.n6922 D.t94 7.493
R13520 D.n6908 D.t2606 7.493
R13521 D.n6894 D.t2459 7.493
R13522 D.n6880 D.t3019 7.493
R13523 D.n6866 D.t1254 7.493
R13524 D.n6852 D.t1891 7.493
R13525 D.n6838 D.t829 7.493
R13526 D.n6824 D.t1500 7.493
R13527 D.n6810 D.t1179 7.493
R13528 D.n6796 D.t2852 7.493
R13529 D.n7002 D.t4176 7.493
R13530 D.n7018 D.t1354 7.493
R13531 D.n7186 D.t3529 7.493
R13532 D.n7172 D.t3221 7.493
R13533 D.n7158 D.t2473 7.493
R13534 D.n7144 D.t3154 7.493
R13535 D.n7130 D.t2373 7.493
R13536 D.n7116 D.t3199 7.493
R13537 D.n7102 D.t3880 7.493
R13538 D.n7088 D.t771 7.493
R13539 D.n7074 D.t1798 7.493
R13540 D.n7060 D.t1076 7.493
R13541 D.n7046 D.t943 7.493
R13542 D.n7032 D.t159 7.493
R13543 D.n7210 D.t1173 7.493
R13544 D.n7226 D.t2800 7.493
R13545 D.n7366 D.t4204 7.493
R13546 D.n7352 D.t215 7.493
R13547 D.n7338 D.t977 7.493
R13548 D.n7324 D.t2392 7.493
R13549 D.n7310 D.t2728 7.493
R13550 D.n7296 D.t3473 7.493
R13551 D.n7282 D.t547 7.493
R13552 D.n7268 D.t264 7.493
R13553 D.n7254 D.t1831 7.493
R13554 D.n7240 D.t2432 7.493
R13555 D.n7390 D.t3649 7.493
R13556 D.n7406 D.t3341 7.493
R13557 D.n7518 D.t1243 7.493
R13558 D.n7504 D.t2790 7.493
R13559 D.n7490 D.t1682 7.493
R13560 D.n7476 D.t1417 7.493
R13561 D.n7462 D.t4500 7.493
R13562 D.n7448 D.t2267 7.493
R13563 D.n7434 D.t3776 7.493
R13564 D.n7420 D.t3573 7.493
R13565 D.n7542 D.t645 7.493
R13566 D.n7558 D.t3638 7.493
R13567 D.n7642 D.t3612 7.493
R13568 D.n7628 D.t3896 7.493
R13569 D.n7614 D.t2322 7.493
R13570 D.n7600 D.t3041 7.493
R13571 D.n7586 D.t2702 7.493
R13572 D.n7572 D.t1409 7.493
R13573 D.n7666 D.t3399 7.493
R13574 D.n7682 D.t1140 7.493
R13575 D.n7738 D.t2897 7.493
R13576 D.n7724 D.t1741 7.493
R13577 D.n7710 D.t866 7.493
R13578 D.n7696 D.t3915 7.493
R13579 D.n7761 D.t797 7.493
R13580 D.n7777 D.t3307 7.493
R13581 D.n7805 D.t4378 7.493
R13582 D.n7791 D.t1750 7.493
R13583 D.n7853 D.t4164 7.099
R13584 D.n7817 D.t406 7.099
R13585 D.n7838 D.t2405 7.099
R13586 D.n7828 D.t2218 7.099
R13587 D.n449 D.t3667 7.099
R13588 D.n440 D.t2090 7.099
R13589 D.n31 D.t4117 7.099
R13590 D.n7958 D.t1796 7.099
R13591 D.n7943 D.t2675 7.099
R13592 D.n14063 D.t2447 7.099
R13593 D.n14045 D.t4046 7.099
R13594 D.n14027 D.t350 7.099
R13595 D.n14009 D.t3769 7.099
R13596 D.n13991 D.t2789 7.099
R13597 D.n13973 D.t4283 7.099
R13598 D.n13955 D.t4416 7.099
R13599 D.n13937 D.t3652 7.099
R13600 D.n13919 D.t103 7.099
R13601 D.n13901 D.t2968 7.099
R13602 D.n13883 D.t4263 7.099
R13603 D.n13865 D.t142 7.099
R13604 D.n13847 D.t2512 7.099
R13605 D.n13829 D.t3161 7.099
R13606 D.n13811 D.t3737 7.099
R13607 D.n13793 D.t1994 7.099
R13608 D.n13775 D.t1880 7.099
R13609 D.n13757 D.t3873 7.099
R13610 D.n13739 D.t602 7.099
R13611 D.n13721 D.t2550 7.099
R13612 D.n13703 D.t2819 7.099
R13613 D.n13684 D.t3592 7.099
R13614 D.n13694 D.t4397 7.099
R13615 D.n13712 D.t4087 7.099
R13616 D.n13730 D.t1771 7.099
R13617 D.n13748 D.t3555 7.099
R13618 D.n13766 D.t3063 7.099
R13619 D.n13784 D.t3648 7.099
R13620 D.n13802 D.t1183 7.099
R13621 D.n13820 D.t29 7.099
R13622 D.n13838 D.t4365 7.099
R13623 D.n13856 D.t2388 7.099
R13624 D.n13874 D.t1348 7.099
R13625 D.n13892 D.t769 7.099
R13626 D.n13910 D.t3340 7.099
R13627 D.n13928 D.t1870 7.099
R13628 D.n13946 D.t88 7.099
R13629 D.n13964 D.t1746 7.099
R13630 D.n13982 D.t1020 7.099
R13631 D.n14000 D.t1534 7.099
R13632 D.n14018 D.t3860 7.099
R13633 D.n14036 D.t603 7.099
R13634 D.n14054 D.t1681 7.099
R13635 D.n14076 D.t4467 7.099
R13636 D.n13209 D.t1960 7.099
R13637 D.n13229 D.t3404 7.099
R13638 D.n13249 D.t1476 7.099
R13639 D.n13269 D.t1122 7.099
R13640 D.n13289 D.t1269 7.099
R13641 D.n13309 D.t2000 7.099
R13642 D.n13329 D.t462 7.099
R13643 D.n13349 D.t1488 7.099
R13644 D.n13369 D.t1996 7.099
R13645 D.n13389 D.t3944 7.099
R13646 D.n13409 D.t4255 7.099
R13647 D.n13429 D.t1453 7.099
R13648 D.n13449 D.t2264 7.099
R13649 D.n13469 D.t3784 7.099
R13650 D.n13489 D.t4367 7.099
R13651 D.n13509 D.t2545 7.099
R13652 D.n13529 D.t1109 7.099
R13653 D.n13549 D.t2468 7.099
R13654 D.n13569 D.t3971 7.099
R13655 D.n13589 D.t2450 7.099
R13656 D.n13609 D.t1555 7.099
R13657 D.n13598 D.t3377 7.099
R13658 D.n13578 D.t1825 7.099
R13659 D.n13558 D.t3094 7.099
R13660 D.n13538 D.t3953 7.099
R13661 D.n13518 D.t2431 7.099
R13662 D.n13498 D.t1516 7.099
R13663 D.n13478 D.t3616 7.099
R13664 D.n13458 D.t3142 7.099
R13665 D.n13438 D.t3373 7.099
R13666 D.n13418 D.t3204 7.099
R13667 D.n13398 D.t2875 7.099
R13668 D.n13378 D.t1936 7.099
R13669 D.n13358 D.t1202 7.099
R13670 D.n13338 D.t38 7.099
R13671 D.n13318 D.t4456 7.099
R13672 D.n13298 D.t4374 7.099
R13673 D.n13278 D.t3422 7.099
R13674 D.n13258 D.t3454 7.099
R13675 D.n13238 D.t4067 7.099
R13676 D.n13218 D.t4209 7.099
R13677 D.n13193 D.t2517 7.099
R13678 D.n13100 D.t2510 7.099
R13679 D.n13082 D.t1950 7.099
R13680 D.n13064 D.t2300 7.099
R13681 D.n13046 D.t1767 7.099
R13682 D.n13028 D.t15 7.099
R13683 D.n13010 D.t4136 7.099
R13684 D.n12992 D.t1617 7.099
R13685 D.n12974 D.t1035 7.099
R13686 D.n12956 D.t1764 7.099
R13687 D.n12938 D.t2501 7.099
R13688 D.n12920 D.t2637 7.099
R13689 D.n12902 D.t2157 7.099
R13690 D.n12884 D.t622 7.099
R13691 D.n12866 D.t441 7.099
R13692 D.n12848 D.t2815 7.099
R13693 D.n12830 D.t4343 7.099
R13694 D.n12812 D.t2940 7.099
R13695 D.n12794 D.t2094 7.099
R13696 D.n12776 D.t2718 7.099
R13697 D.n12757 D.t4228 7.099
R13698 D.n12767 D.t1860 7.099
R13699 D.n12785 D.t806 7.099
R13700 D.n12803 D.t285 7.099
R13701 D.n12821 D.t1938 7.099
R13702 D.n12839 D.t133 7.099
R13703 D.n12857 D.t4243 7.099
R13704 D.n12875 D.t3304 7.099
R13705 D.n12893 D.t2248 7.099
R13706 D.n12911 D.t306 7.099
R13707 D.n12929 D.t2886 7.099
R13708 D.n12947 D.t4320 7.099
R13709 D.n12965 D.t3578 7.099
R13710 D.n12983 D.t2801 7.099
R13711 D.n13001 D.t3014 7.099
R13712 D.n13019 D.t3651 7.099
R13713 D.n13037 D.t480 7.099
R13714 D.n13055 D.t1737 7.099
R13715 D.n13073 D.t923 7.099
R13716 D.n13091 D.t3369 7.099
R13717 D.n13112 D.t4099 7.099
R13718 D.n12326 D.t2004 7.099
R13719 D.n12346 D.t3656 7.099
R13720 D.n12366 D.t3496 7.099
R13721 D.n12386 D.t4404 7.099
R13722 D.n12406 D.t3116 7.099
R13723 D.n12426 D.t4364 7.099
R13724 D.n12446 D.t4348 7.099
R13725 D.n12466 D.t4436 7.099
R13726 D.n12486 D.t3772 7.099
R13727 D.n12506 D.t3886 7.099
R13728 D.n12526 D.t1613 7.099
R13729 D.n12546 D.t4177 7.099
R13730 D.n12566 D.t2600 7.099
R13731 D.n12586 D.t2354 7.099
R13732 D.n12606 D.t3729 7.099
R13733 D.n12626 D.t2661 7.099
R13734 D.n12646 D.t4002 7.099
R13735 D.n12666 D.t1912 7.099
R13736 D.n12686 D.t865 7.099
R13737 D.n12675 D.t1833 7.099
R13738 D.n12655 D.t1867 7.099
R13739 D.n12635 D.t2741 7.099
R13740 D.n12615 D.t4415 7.099
R13741 D.n12595 D.t2931 7.099
R13742 D.n12575 D.t863 7.099
R13743 D.n12555 D.t1136 7.099
R13744 D.n12535 D.t4479 7.099
R13745 D.n12515 D.t4346 7.099
R13746 D.n12495 D.t3848 7.099
R13747 D.n12475 D.t1856 7.099
R13748 D.n12455 D.t3646 7.099
R13749 D.n12435 D.t1176 7.099
R13750 D.n12415 D.t249 7.099
R13751 D.n12395 D.t1504 7.099
R13752 D.n12375 D.t3723 7.099
R13753 D.n12355 D.t1050 7.099
R13754 D.n12335 D.t2028 7.099
R13755 D.n12310 D.t2244 7.099
R13756 D.n12215 D.t2837 7.099
R13757 D.n12197 D.t1626 7.099
R13758 D.n12179 D.t1470 7.099
R13759 D.n12161 D.t252 7.099
R13760 D.n12143 D.t1203 7.099
R13761 D.n12125 D.t1571 7.099
R13762 D.n12107 D.t590 7.099
R13763 D.n12089 D.t1475 7.099
R13764 D.n12071 D.t1365 7.099
R13765 D.n12053 D.t2335 7.099
R13766 D.n12035 D.t1817 7.099
R13767 D.n12017 D.t3518 7.099
R13768 D.n11999 D.t2185 7.099
R13769 D.n11981 D.t2231 7.099
R13770 D.n11963 D.t811 7.099
R13771 D.n11945 D.t2519 7.099
R13772 D.n11927 D.t3933 7.099
R13773 D.n11908 D.t1367 7.099
R13774 D.n11918 D.t1119 7.099
R13775 D.n11936 D.t3355 7.099
R13776 D.n11954 D.t2816 7.099
R13777 D.n11972 D.t1242 7.099
R13778 D.n11990 D.t2319 7.099
R13779 D.n12008 D.t188 7.099
R13780 D.n12026 D.t3289 7.099
R13781 D.n12044 D.t2929 7.099
R13782 D.n12062 D.t2784 7.099
R13783 D.n12080 D.t1196 7.099
R13784 D.n12098 D.t110 7.099
R13785 D.n12116 D.t1783 7.099
R13786 D.n12134 D.t1006 7.099
R13787 D.n12152 D.t2608 7.099
R13788 D.n12170 D.t3318 7.099
R13789 D.n12188 D.t4280 7.099
R13790 D.n12206 D.t4259 7.099
R13791 D.n12228 D.t1768 7.099
R13792 D.n11517 D.t2752 7.099
R13793 D.n11537 D.t1197 7.099
R13794 D.n11557 D.t150 7.099
R13795 D.n11577 D.t1004 7.099
R13796 D.n11597 D.t1787 7.099
R13797 D.n11617 D.t3261 7.099
R13798 D.n11637 D.t1257 7.099
R13799 D.n11657 D.t495 7.099
R13800 D.n11677 D.t1967 7.099
R13801 D.n11697 D.t106 7.099
R13802 D.n11717 D.t374 7.099
R13803 D.n11737 D.t275 7.099
R13804 D.n11757 D.t3532 7.099
R13805 D.n11777 D.t2668 7.099
R13806 D.n11797 D.t2375 7.099
R13807 D.n11817 D.t3644 7.099
R13808 D.n11837 D.t13 7.099
R13809 D.n11826 D.t2945 7.099
R13810 D.n11806 D.t4145 7.099
R13811 D.n11786 D.t187 7.099
R13812 D.n11766 D.t1356 7.099
R13813 D.n11746 D.t4497 7.099
R13814 D.n11726 D.t3874 7.099
R13815 D.n11706 D.t3981 7.099
R13816 D.n11686 D.t2891 7.099
R13817 D.n11666 D.t3136 7.099
R13818 D.n11646 D.t2922 7.099
R13819 D.n11626 D.t4443 7.099
R13820 D.n11606 D.t3866 7.099
R13821 D.n11586 D.t4441 7.099
R13822 D.n11566 D.t4153 7.099
R13823 D.n11546 D.t870 7.099
R13824 D.n11526 D.t1923 7.099
R13825 D.n11503 D.t691 7.099
R13826 D.n11416 D.t633 7.099
R13827 D.n11398 D.t4393 7.099
R13828 D.n11380 D.t4457 7.099
R13829 D.n11362 D.t3433 7.099
R13830 D.n11344 D.t2892 7.099
R13831 D.n11326 D.t4277 7.099
R13832 D.n11308 D.t768 7.099
R13833 D.n11290 D.t2547 7.099
R13834 D.n11272 D.t4035 7.099
R13835 D.n11254 D.t237 7.099
R13836 D.n11236 D.t588 7.099
R13837 D.n11218 D.t1872 7.099
R13838 D.n11200 D.t2810 7.099
R13839 D.n11182 D.t2201 7.099
R13840 D.n11164 D.t541 7.099
R13841 D.n11145 D.t774 7.099
R13842 D.n11155 D.t2333 7.099
R13843 D.n11173 D.t1975 7.099
R13844 D.n11191 D.t663 7.099
R13845 D.n11209 D.t2408 7.099
R13846 D.n11227 D.t583 7.099
R13847 D.n11245 D.t618 7.099
R13848 D.n11263 D.t3211 7.099
R13849 D.n11281 D.t2380 7.099
R13850 D.n11299 D.t2228 7.099
R13851 D.n11317 D.t973 7.099
R13852 D.n11335 D.t3248 7.099
R13853 D.n11353 D.t1429 7.099
R13854 D.n11371 D.t996 7.099
R13855 D.n11389 D.t911 7.099
R13856 D.n11407 D.t1299 7.099
R13857 D.n11429 D.t1531 7.099
R13858 D.n10794 D.t233 7.099
R13859 D.n10814 D.t999 7.099
R13860 D.n10834 D.t1444 7.099
R13861 D.n10854 D.t3955 7.099
R13862 D.n10874 D.t1174 7.099
R13863 D.n10894 D.t940 7.099
R13864 D.n10914 D.t824 7.099
R13865 D.n10934 D.t208 7.099
R13866 D.n10954 D.t739 7.099
R13867 D.n10974 D.t703 7.099
R13868 D.n10994 D.t192 7.099
R13869 D.n11014 D.t379 7.099
R13870 D.n11034 D.t1640 7.099
R13871 D.n11054 D.t3985 7.099
R13872 D.n11074 D.t3083 7.099
R13873 D.n11063 D.t86 7.099
R13874 D.n11043 D.t4058 7.099
R13875 D.n11023 D.t1661 7.099
R13876 D.n11003 D.t2460 7.099
R13877 D.n10983 D.t1987 7.099
R13878 D.n10963 D.t1337 7.099
R13879 D.n10943 D.t4506 7.099
R13880 D.n10923 D.t2203 7.099
R13881 D.n10903 D.t4042 7.099
R13882 D.n10883 D.t1013 7.099
R13883 D.n10863 D.t1910 7.099
R13884 D.n10843 D.t519 7.099
R13885 D.n10823 D.t4126 7.099
R13886 D.n10803 D.t465 7.099
R13887 D.n10780 D.t3339 7.099
R13888 D.n10697 D.t1819 7.099
R13889 D.n10679 D.t900 7.099
R13890 D.n10661 D.t1986 7.099
R13891 D.n10643 D.t1008 7.099
R13892 D.n10625 D.t2116 7.099
R13893 D.n10607 D.t731 7.099
R13894 D.n10589 D.t2320 7.099
R13895 D.n10571 D.t1532 7.099
R13896 D.n10553 D.t1619 7.099
R13897 D.n10535 D.t4401 7.099
R13898 D.n10517 D.t3747 7.099
R13899 D.n10499 D.t1622 7.099
R13900 D.n10481 D.t2592 7.099
R13901 D.n10462 D.t2120 7.099
R13902 D.n10472 D.t2813 7.099
R13903 D.n10490 D.t3696 7.099
R13904 D.n10508 D.t1977 7.099
R13905 D.n10526 D.t3917 7.099
R13906 D.n10544 D.t3030 7.099
R13907 D.n10562 D.t3001 7.099
R13908 D.n10580 D.t559 7.099
R13909 D.n10598 D.t1641 7.099
R13910 D.n10616 D.t801 7.099
R13911 D.n10634 D.t4078 7.099
R13912 D.n10652 D.t3275 7.099
R13913 D.n10670 D.t4452 7.099
R13914 D.n10688 D.t4241 7.099
R13915 D.n10710 D.t2619 7.099
R13916 D.n10151 D.t2161 7.099
R13917 D.n10171 D.t4433 7.099
R13918 D.n10191 D.t3505 7.099
R13919 D.n10211 D.t4017 7.099
R13920 D.n10231 D.t2186 7.099
R13921 D.n10251 D.t1688 7.099
R13922 D.n10271 D.t717 7.099
R13923 D.n10291 D.t2530 7.099
R13924 D.n10311 D.t4023 7.099
R13925 D.n10331 D.t3134 7.099
R13926 D.n10351 D.t762 7.099
R13927 D.n10371 D.t438 7.099
R13928 D.n10391 D.t4019 7.099
R13929 D.n10380 D.t413 7.099
R13930 D.n10360 D.t1064 7.099
R13931 D.n10340 D.t2678 7.099
R13932 D.n10320 D.t2941 7.099
R13933 D.n10300 D.t2371 7.099
R13934 D.n10280 D.t2127 7.099
R13935 D.n10260 D.t1868 7.099
R13936 D.n10240 D.t955 7.099
R13937 D.n10220 D.t344 7.099
R13938 D.n10200 D.t3191 7.099
R13939 D.n10180 D.t1217 7.099
R13940 D.n10160 D.t2515 7.099
R13941 D.n10135 D.t1063 7.099
R13942 D.n10058 D.t199 7.099
R13943 D.n10040 D.t2552 7.099
R13944 D.n10022 D.t1926 7.099
R13945 D.n10004 D.t277 7.099
R13946 D.n9986 D.t722 7.099
R13947 D.n9968 D.t913 7.099
R13948 D.n9950 D.t453 7.099
R13949 D.n9932 D.t2325 7.099
R13950 D.n9914 D.t679 7.099
R13951 D.n9896 D.t932 7.099
R13952 D.n9878 D.t3130 7.099
R13953 D.n9859 D.t1929 7.099
R13954 D.n9869 D.t2751 7.099
R13955 D.n9887 D.t4115 7.099
R13956 D.n9905 D.t326 7.099
R13957 D.n9923 D.t2415 7.099
R13958 D.n9941 D.t2194 7.099
R13959 D.n9959 D.t4027 7.099
R13960 D.n9977 D.t2542 7.099
R13961 D.n9995 D.t765 7.099
R13962 D.n10013 D.t1696 7.099
R13963 D.n10031 D.t3517 7.099
R13964 D.n10049 D.t2301 7.099
R13965 D.n10070 D.t1733 7.099
R13966 D.n9588 D.t4303 7.099
R13967 D.n9608 D.t468 7.099
R13968 D.n9628 D.t597 7.099
R13969 D.n9648 D.t989 7.099
R13970 D.n9668 D.t2107 7.099
R13971 D.n9688 D.t2304 7.099
R13972 D.n9708 D.t3969 7.099
R13973 D.n9728 D.t654 7.099
R13974 D.n9748 D.t1314 7.099
R13975 D.n9768 D.t1309 7.099
R13976 D.n9788 D.t1361 7.099
R13977 D.n9777 D.t2950 7.099
R13978 D.n9757 D.t749 7.099
R13979 D.n9737 D.t970 7.099
R13980 D.n9717 D.t4471 7.099
R13981 D.n9697 D.t735 7.099
R13982 D.n9677 D.t204 7.099
R13983 D.n9657 D.t1346 7.099
R13984 D.n9637 D.t933 7.099
R13985 D.n9617 D.t571 7.099
R13986 D.n9597 D.t4269 7.099
R13987 D.n9572 D.t2658 7.099
R13988 D.n9493 D.t1129 7.099
R13989 D.n9475 D.t702 7.099
R13990 D.n9457 D.t2063 7.099
R13991 D.n9439 D.t4010 7.099
R13992 D.n9421 D.t2173 7.099
R13993 D.n9403 D.t1376 7.099
R13994 D.n9385 D.t708 7.099
R13995 D.n9367 D.t2068 7.099
R13996 D.n9349 D.t4014 7.099
R13997 D.n9330 D.t1380 7.099
R13998 D.n9340 D.t2026 7.099
R13999 D.n9358 D.t1185 7.099
R14000 D.n9376 D.t1662 7.099
R14001 D.n9394 D.t1385 7.099
R14002 D.n9412 D.t1163 7.099
R14003 D.n9430 D.t3930 7.099
R14004 D.n9448 D.t485 7.099
R14005 D.n9466 D.t1273 7.099
R14006 D.n9484 D.t1265 7.099
R14007 D.n9506 D.t3614 7.099
R14008 D.n9099 D.t3847 7.099
R14009 D.n9119 D.t395 7.099
R14010 D.n9139 D.t1568 7.099
R14011 D.n9159 D.t1918 7.099
R14012 D.n9179 D.t1389 7.099
R14013 D.n9199 D.t362 7.099
R14014 D.n9219 D.t689 7.099
R14015 D.n9239 D.t1908 7.099
R14016 D.n9259 D.t809 7.099
R14017 D.n9248 D.t3989 7.099
R14018 D.n9228 D.t2260 7.099
R14019 D.n9208 D.t1974 7.099
R14020 D.n9188 D.t40 7.099
R14021 D.n9168 D.t714 7.099
R14022 D.n9148 D.t1684 7.099
R14023 D.n9128 D.t791 7.099
R14024 D.n9108 D.t3458 7.099
R14025 D.n9085 D.t1262 7.099
R14026 D.n9014 D.t4468 7.099
R14027 D.n8996 D.t1634 7.099
R14028 D.n8978 D.t503 7.099
R14029 D.n8960 D.t2578 7.099
R14030 D.n8942 D.t2088 7.099
R14031 D.n8924 D.t220 7.099
R14032 D.n8906 D.t2018 7.099
R14033 D.n8887 D.t1875 7.099
R14034 D.n8897 D.t887 7.099
R14035 D.n8915 D.t2154 7.099
R14036 D.n8933 D.t3993 7.099
R14037 D.n8951 D.t2052 7.099
R14038 D.n8969 D.t904 7.099
R14039 D.n8987 D.t605 7.099
R14040 D.n9005 D.t3924 7.099
R14041 D.n9027 D.t741 7.099
R14042 D.n8696 D.t3488 7.099
R14043 D.n8716 D.t61 7.099
R14044 D.n8736 D.t2055 7.099
R14045 D.n8756 D.t4000 7.099
R14046 D.n8776 D.t2159 7.099
R14047 D.n8796 D.t1372 7.099
R14048 D.n8816 D.t3353 7.099
R14049 D.n8805 D.t734 7.099
R14050 D.n8785 D.t805 7.099
R14051 D.n8765 D.t920 7.099
R14052 D.n8745 D.t945 7.099
R14053 D.n8725 D.t2594 7.099
R14054 D.n8705 D.t881 7.099
R14055 D.n8680 D.t3786 7.099
R14056 D.n8615 D.t3601 7.099
R14057 D.n8597 D.t408 7.099
R14058 D.n8579 D.t846 7.099
R14059 D.n8561 D.t1615 7.099
R14060 D.n8543 D.t1593 7.099
R14061 D.n8524 D.t3303 7.099
R14062 D.n8534 D.t798 7.099
R14063 D.n8552 D.t2314 7.099
R14064 D.n8570 D.t1161 7.099
R14065 D.n8588 D.t1342 7.099
R14066 D.n8606 D.t3492 7.099
R14067 D.n8627 D.t2616 7.099
R14068 D.n8373 D.t2245 7.099
R14069 D.n8393 D.t1542 7.099
R14070 D.n8413 D.t2341 7.099
R14071 D.n8433 D.t2454 7.099
R14072 D.n8453 D.t1636 7.099
R14073 D.n8442 D.t3240 7.099
R14074 D.n8422 D.t1700 7.099
R14075 D.n8402 D.t423 7.099
R14076 D.n8382 D.t1042 7.099
R14077 D.n8357 D.t4448 7.099
R14078 D.n8290 D.t3867 7.099
R14079 D.n8272 D.t52 7.099
R14080 D.n8254 D.t2047 7.099
R14081 D.n8235 D.t3890 7.099
R14082 D.n8245 D.t3501 7.099
R14083 D.n8263 D.t536 7.099
R14084 D.n8281 D.t3513 7.099
R14085 D.n8303 D.t2743 7.099
R14086 D.n8124 D.t1158 7.099
R14087 D.n8144 D.t928 7.099
R14088 D.n8164 D.t1401 7.099
R14089 D.n8153 D.t4096 7.099
R14090 D.n8133 D.t1283 7.099
R14091 D.n8110 D.t830 7.099
R14092 D.n8051 D.t3570 7.099
R14093 D.n8032 D.t3919 7.099
R14094 D.n8042 D.t3717 7.099
R14095 D.n8064 D.t772 7.099
R14096 D.n53 D.t651 7.099
R14097 D.n62 D.t125 7.099
R14098 D.n71 D.t28 7.099
R14099 D.n80 D.t4116 7.099
R14100 D.n89 D.t3329 7.099
R14101 D.n98 D.t3668 7.099
R14102 D.n107 D.t1368 7.099
R14103 D.n116 D.t837 7.099
R14104 D.n125 D.t149 7.099
R14105 D.n134 D.t562 7.099
R14106 D.n143 D.t3292 7.099
R14107 D.n152 D.t1653 7.099
R14108 D.n161 D.t649 7.099
R14109 D.n170 D.t1168 7.099
R14110 D.n179 D.t2401 7.099
R14111 D.n188 D.t745 7.099
R14112 D.n197 D.t1142 7.099
R14113 D.n206 D.t4282 7.099
R14114 D.n215 D.t2957 7.099
R14115 D.n224 D.t1738 7.099
R14116 D.n233 D.t1441 7.099
R14117 D.n242 D.t2271 7.099
R14118 D.n251 D.t3920 7.099
R14119 D.n260 D.t1591 7.099
R14120 D.n269 D.t3228 7.099
R14121 D.n278 D.t4196 7.099
R14122 D.n287 D.t4435 7.099
R14123 D.n296 D.t1755 7.099
R14124 D.n305 D.t1801 7.099
R14125 D.n314 D.t1024 7.099
R14126 D.n323 D.t213 7.099
R14127 D.n332 D.t1569 7.099
R14128 D.n341 D.t832 7.099
R14129 D.n350 D.t3287 7.099
R14130 D.n359 D.t3278 7.099
R14131 D.n368 D.t66 7.099
R14132 D.n377 D.t3393 7.099
R14133 D.n386 D.t2342 7.099
R14134 D.n395 D.t4052 7.099
R14135 D.n404 D.t750 7.099
R14136 D.n413 D.t3239 7.099
R14137 D.n422 D.t3966 7.099
R14138 D.n431 D.t3392 7.099
R14139 D.n525 D.t4304 7.099
R14140 D.n541 D.t4106 7.099
R14141 D.n513 D.t3734 7.099
R14142 D.n1129 D.t1068 7.099
R14143 D.n1115 D.t3802 7.099
R14144 D.n1101 D.t1012 7.099
R14145 D.n1087 D.t1793 7.099
R14146 D.n1073 D.t1041 7.099
R14147 D.n1059 D.t4462 7.099
R14148 D.n1045 D.t3126 7.099
R14149 D.n1031 D.t4432 7.099
R14150 D.n1017 D.t1574 7.099
R14151 D.n1003 D.t74 7.099
R14152 D.n989 D.t3507 7.099
R14153 D.n975 D.t1691 7.099
R14154 D.n961 D.t3434 7.099
R14155 D.n947 D.t2937 7.099
R14156 D.n933 D.t1116 7.099
R14157 D.n919 D.t1459 7.099
R14158 D.n905 D.t3621 7.099
R14159 D.n891 D.t2564 7.099
R14160 D.n877 D.t4422 7.099
R14161 D.n863 D.t4379 7.099
R14162 D.n849 D.t3683 7.099
R14163 D.n835 D.t1404 7.099
R14164 D.n821 D.t3227 7.099
R14165 D.n807 D.t2268 7.099
R14166 D.n793 D.t1791 7.099
R14167 D.n779 D.t180 7.099
R14168 D.n765 D.t3752 7.099
R14169 D.n751 D.t4188 7.099
R14170 D.n737 D.t472 7.099
R14171 D.n723 D.t3320 7.099
R14172 D.n709 D.t3593 7.099
R14173 D.n695 D.t2834 7.099
R14174 D.n681 D.t1410 7.099
R14175 D.n667 D.t4137 7.099
R14176 D.n653 D.t1736 7.099
R14177 D.n639 D.t419 7.099
R14178 D.n625 D.t454 7.099
R14179 D.n611 D.t1040 7.099
R14180 D.n597 D.t295 7.099
R14181 D.n583 D.t1498 7.099
R14182 D.n569 D.t1814 7.099
R14183 D.n555 D.t3902 7.099
R14184 D.n1152 D.t114 7.099
R14185 D.n1168 D.t1420 7.099
R14186 D.n1143 D.t4168 7.099
R14187 D.n1728 D.t972 7.099
R14188 D.n1714 D.t4072 7.099
R14189 D.n1700 D.t1325 7.099
R14190 D.n1686 D.t1984 7.099
R14191 D.n1672 D.t2697 7.099
R14192 D.n1658 D.t834 7.099
R14193 D.n1644 D.t4186 7.099
R14194 D.n1630 D.t2193 7.099
R14195 D.n1616 D.t3484 7.099
R14196 D.n1602 D.t2315 7.099
R14197 D.n1588 D.t3916 7.099
R14198 D.n1574 D.t288 7.099
R14199 D.n1560 D.t577 7.099
R14200 D.n1546 D.t3572 7.099
R14201 D.n1532 D.t1834 7.099
R14202 D.n1518 D.t231 7.099
R14203 D.n1504 D.t1017 7.099
R14204 D.n1490 D.t1790 7.099
R14205 D.n1476 D.t3511 7.099
R14206 D.n1462 D.t3895 7.099
R14207 D.n1448 D.t2806 7.099
R14208 D.n1434 D.t3115 7.099
R14209 D.n1420 D.t785 7.099
R14210 D.n1406 D.t1406 7.099
R14211 D.n1392 D.t1980 7.099
R14212 D.n1378 D.t635 7.099
R14213 D.n1364 D.t969 7.099
R14214 D.n1350 D.t1072 7.099
R14215 D.n1336 D.t3254 7.099
R14216 D.n1322 D.t1208 7.099
R14217 D.n1308 D.t3284 7.099
R14218 D.n1294 D.t105 7.099
R14219 D.n1280 D.t3502 7.099
R14220 D.n1266 D.t1159 7.099
R14221 D.n1252 D.t3640 7.099
R14222 D.n1238 D.t1341 7.099
R14223 D.n1224 D.t407 7.099
R14224 D.n1210 D.t1679 7.099
R14225 D.n1196 D.t1723 7.099
R14226 D.n1182 D.t3834 7.099
R14227 D.n1751 D.t4049 7.099
R14228 D.n1767 D.t3898 7.099
R14229 D.n1742 D.t4162 7.099
R14230 D.n2299 D.t931 7.099
R14231 D.n2285 D.t1905 7.099
R14232 D.n2271 D.t1659 7.099
R14233 D.n2257 D.t214 7.099
R14234 D.n2243 D.t1028 7.099
R14235 D.n2229 D.t2360 7.099
R14236 D.n2215 D.t3493 7.099
R14237 D.n2201 D.t2641 7.099
R14238 D.n2187 D.t2971 7.099
R14239 D.n2173 D.t3842 7.099
R14240 D.n2159 D.t4484 7.099
R14241 D.n2145 D.t17 7.099
R14242 D.n2131 D.t3580 7.099
R14243 D.n2117 D.t4171 7.099
R14244 D.n2103 D.t3541 7.099
R14245 D.n2089 D.t4069 7.099
R14246 D.n2075 D.t1059 7.099
R14247 D.n2061 D.t1557 7.099
R14248 D.n2047 D.t991 7.099
R14249 D.n2033 D.t1001 7.099
R14250 D.n2019 D.t4118 7.099
R14251 D.n2005 D.t4125 7.099
R14252 D.n1991 D.t4147 7.099
R14253 D.n1977 D.t3124 7.099
R14254 D.n1963 D.t3272 7.099
R14255 D.n1949 D.t1820 7.099
R14256 D.n1935 D.t2689 7.099
R14257 D.n1921 D.t3664 7.099
R14258 D.n1907 D.t1744 7.099
R14259 D.n1893 D.t1812 7.099
R14260 D.n1879 D.t1019 7.099
R14261 D.n1865 D.t917 7.099
R14262 D.n1851 D.t1277 7.099
R14263 D.n1837 D.t944 7.099
R14264 D.n1823 D.t3711 7.099
R14265 D.n1809 D.t1526 7.099
R14266 D.n1795 D.t60 7.099
R14267 D.n1781 D.t3516 7.099
R14268 D.n2322 D.t754 7.099
R14269 D.n2338 D.t1633 7.099
R14270 D.n2313 D.t4011 7.099
R14271 D.n2842 D.t4335 7.099
R14272 D.n2828 D.t2709 7.099
R14273 D.n2814 D.t1308 7.099
R14274 D.n2800 D.t890 7.099
R14275 D.n2786 D.t2757 7.099
R14276 D.n2772 D.t1892 7.099
R14277 D.n2758 D.t1295 7.099
R14278 D.n2744 D.t671 7.099
R14279 D.n2730 D.t4359 7.099
R14280 D.n2716 D.t637 7.099
R14281 D.n2702 D.t189 7.099
R14282 D.n2688 D.t2620 7.099
R14283 D.n2674 D.t4159 7.099
R14284 D.n2660 D.t4181 7.099
R14285 D.n2646 D.t3685 7.099
R14286 D.n2632 D.t1566 7.099
R14287 D.n2618 D.t1886 7.099
R14288 D.n2604 D.t22 7.099
R14289 D.n2590 D.t1034 7.099
R14290 D.n2576 D.t1753 7.099
R14291 D.n2562 D.t3230 7.099
R14292 D.n2548 D.t1899 7.099
R14293 D.n2534 D.t3127 7.099
R14294 D.n2520 D.t4045 7.099
R14295 D.n2506 D.t886 7.099
R14296 D.n2492 D.t1616 7.099
R14297 D.n2478 D.t1852 7.099
R14298 D.n2464 D.t4284 7.099
R14299 D.n2450 D.t966 7.099
R14300 D.n2436 D.t3994 7.099
R14301 D.n2422 D.t535 7.099
R14302 D.n2408 D.t2050 7.099
R14303 D.n2394 D.t3770 7.099
R14304 D.n2380 D.t56 7.099
R14305 D.n2366 D.t436 7.099
R14306 D.n2352 D.t3889 7.099
R14307 D.n2865 D.t3213 7.099
R14308 D.n2881 D.t3362 7.099
R14309 D.n2856 D.t1103 7.099
R14310 D.n3357 D.t3077 7.099
R14311 D.n3343 D.t3990 7.099
R14312 D.n3329 D.t914 7.099
R14313 D.n3315 D.t2910 7.099
R14314 D.n3301 D.t162 7.099
R14315 D.n3287 D.t3735 7.099
R14316 D.n3273 D.t2672 7.099
R14317 D.n3259 D.t2281 7.099
R14318 D.n3245 D.t3760 7.099
R14319 D.n3231 D.t2491 7.099
R14320 D.n3217 D.t1286 7.099
R14321 D.n3203 D.t1944 7.099
R14322 D.n3189 D.t3323 7.099
R14323 D.n3175 D.t4005 7.099
R14324 D.n3161 D.t2870 7.099
R14325 D.n3147 D.t2603 7.099
R14326 D.n3133 D.t1602 7.099
R14327 D.n3119 D.t2149 7.099
R14328 D.n3105 D.t861 7.099
R14329 D.n3091 D.t1087 7.099
R14330 D.n3077 D.t542 7.099
R14331 D.n3063 D.t1770 7.099
R14332 D.n3049 D.t4123 7.099
R14333 D.n3035 D.t2558 7.099
R14334 D.n3021 D.t3407 7.099
R14335 D.n3007 D.t79 7.099
R14336 D.n2993 D.t1047 7.099
R14337 D.n2979 D.t1973 7.099
R14338 D.n2965 D.t46 7.099
R14339 D.n2951 D.t2582 7.099
R14340 D.n2937 D.t1466 7.099
R14341 D.n2923 D.t486 7.099
R14342 D.n2909 D.t3402 7.099
R14343 D.n2895 D.t1635 7.099
R14344 D.n3381 D.t410 7.099
R14345 D.n3397 D.t3232 7.099
R14346 D.n3372 D.t2015 7.099
R14347 D.n3845 D.t760 7.099
R14348 D.n3831 D.t2708 7.099
R14349 D.n3817 D.t3125 7.099
R14350 D.n3803 D.t2833 7.099
R14351 D.n3789 D.t251 7.099
R14352 D.n3775 D.t4293 7.099
R14353 D.n3761 D.t1836 7.099
R14354 D.n3747 D.t2583 7.099
R14355 D.n3733 D.t54 7.099
R14356 D.n3719 D.t3817 7.099
R14357 D.n3705 D.t3293 7.099
R14358 D.n3691 D.t2101 7.099
R14359 D.n3677 D.t2747 7.099
R14360 D.n3663 D.t2725 7.099
R14361 D.n3649 D.t4278 7.099
R14362 D.n3635 D.t157 7.099
R14363 D.n3621 D.t810 7.099
R14364 D.n3607 D.t4338 7.099
R14365 D.n3593 D.t160 7.099
R14366 D.n3579 D.t1250 7.099
R14367 D.n3565 D.t2010 7.099
R14368 D.n3551 D.t221 7.099
R14369 D.n3537 D.t3789 7.099
R14370 D.n3523 D.t366 7.099
R14371 D.n3509 D.t3101 7.099
R14372 D.n3495 D.t2499 7.099
R14373 D.n3481 D.t184 7.099
R14374 D.n3467 D.t1597 7.099
R14375 D.n3453 D.t1378 7.099
R14376 D.n3439 D.t403 7.099
R14377 D.n3425 D.t348 7.099
R14378 D.n3411 D.t2522 7.099
R14379 D.n3869 D.t2058 7.099
R14380 D.n3885 D.t2593 7.099
R14381 D.n3860 D.t2384 7.099
R14382 D.n4305 D.t3268 7.099
R14383 D.n4291 D.t1191 7.099
R14384 D.n4277 D.t3012 7.099
R14385 D.n4263 D.t2525 7.099
R14386 D.n4249 D.t631 7.099
R14387 D.n4235 D.t3359 7.099
R14388 D.n4221 D.t448 7.099
R14389 D.n4207 D.t1213 7.099
R14390 D.n4193 D.t152 7.099
R14391 D.n4179 D.t1497 7.099
R14392 D.n4165 D.t2349 7.099
R14393 D.n4151 D.t2472 7.099
R14394 D.n4137 D.t500 7.099
R14395 D.n4123 D.t1238 7.099
R14396 D.n4109 D.t4084 7.099
R14397 D.n4095 D.t2633 7.099
R14398 D.n4081 D.t4392 7.099
R14399 D.n4067 D.t3028 7.099
R14400 D.n4053 D.t3956 7.099
R14401 D.n4039 D.t690 7.099
R14402 D.n4025 D.t1821 7.099
R14403 D.n4011 D.t1066 7.099
R14404 D.n3997 D.t368 7.099
R14405 D.n3983 D.t2842 7.099
R14406 D.n3969 D.t2418 7.099
R14407 D.n3955 D.t3945 7.099
R14408 D.n3941 D.t447 7.099
R14409 D.n3927 D.t2165 7.099
R14410 D.n3913 D.t2299 7.099
R14411 D.n3899 D.t4003 7.099
R14412 D.n4329 D.t2573 7.099
R14413 D.n4345 D.t912 7.099
R14414 D.n4320 D.t3976 7.099
R14415 D.n4737 D.t191 7.099
R14416 D.n4723 D.t1558 7.099
R14417 D.n4709 D.t699 7.099
R14418 D.n4695 D.t141 7.099
R14419 D.n4681 D.t1913 7.099
R14420 D.n4667 D.t4389 7.099
R14421 D.n4653 D.t3844 7.099
R14422 D.n4639 D.t429 7.099
R14423 D.n4625 D.t75 7.099
R14424 D.n4611 D.t4205 7.099
R14425 D.n4597 D.t1412 7.099
R14426 D.n4583 D.t3424 7.099
R14427 D.n4569 D.t3622 7.099
R14428 D.n4555 D.t1351 7.099
R14429 D.n4541 D.t1584 7.099
R14430 D.n4527 D.t1099 7.099
R14431 D.n4513 D.t3076 7.099
R14432 D.n4499 D.t2070 7.099
R14433 D.n4485 D.t1724 7.099
R14434 D.n4471 D.t2904 7.099
R14435 D.n4457 D.t2437 7.099
R14436 D.n4443 D.t594 7.099
R14437 D.n4429 D.t3018 7.099
R14438 D.n4415 D.t2802 7.099
R14439 D.n4401 D.t1481 7.099
R14440 D.n4387 D.t2964 7.099
R14441 D.n4373 D.t2368 7.099
R14442 D.n4359 D.t2095 7.099
R14443 D.n4761 D.t718 7.099
R14444 D.n4777 D.t1439 7.099
R14445 D.n4752 D.t580 7.099
R14446 D.n5141 D.t566 7.099
R14447 D.n5127 D.t1148 7.099
R14448 D.n5113 D.t2169 7.099
R14449 D.n5099 D.t4485 7.099
R14450 D.n5085 D.t72 7.099
R14451 D.n5071 D.t3281 7.099
R14452 D.n5057 D.t1539 7.099
R14453 D.n5043 D.t4047 7.099
R14454 D.n5029 D.t2316 7.099
R14455 D.n5015 D.t3583 7.099
R14456 D.n5001 D.t3394 7.099
R14457 D.n4987 D.t3533 7.099
R14458 D.n4973 D.t2234 7.099
R14459 D.n4959 D.t3437 7.099
R14460 D.n4945 D.t3699 7.099
R14461 D.n4931 D.t1339 7.099
R14462 D.n4917 D.t63 7.099
R14463 D.n4903 D.t1147 7.099
R14464 D.n4889 D.t3138 7.099
R14465 D.n4875 D.t1463 7.099
R14466 D.n4861 D.t2588 7.099
R14467 D.n4847 D.t1284 7.099
R14468 D.n4833 D.t1381 7.099
R14469 D.n4819 D.t767 7.099
R14470 D.n4805 D.t2777 7.099
R14471 D.n4791 D.t4240 7.099
R14472 D.n5165 D.t3440 7.099
R14473 D.n5181 D.t3328 7.099
R14474 D.n5156 D.t3382 7.099
R14475 D.n5517 D.t2284 7.099
R14476 D.n5503 D.t627 7.099
R14477 D.n5489 D.t2074 7.099
R14478 D.n5475 D.t308 7.099
R14479 D.n5461 D.t4305 7.099
R14480 D.n5447 D.t751 7.099
R14481 D.n5433 D.t2569 7.099
R14482 D.n5419 D.t2859 7.099
R14483 D.n5405 D.t3526 7.099
R14484 D.n5391 D.t2016 7.099
R14485 D.n5377 D.t2887 7.099
R14486 D.n5363 D.t3657 7.099
R14487 D.n5349 D.t591 7.099
R14488 D.n5335 D.t576 7.099
R14489 D.n5321 D.t3942 7.099
R14490 D.n5307 D.t1847 7.099
R14491 D.n5293 D.t146 7.099
R14492 D.n5279 D.t4085 7.099
R14493 D.n5265 D.t3875 7.099
R14494 D.n5251 D.t658 7.099
R14495 D.n5237 D.t3524 7.099
R14496 D.n5223 D.t938 7.099
R14497 D.n5209 D.t2565 7.099
R14498 D.n5195 D.t3497 7.099
R14499 D.n5541 D.t166 7.099
R14500 D.n5557 D.t1784 7.099
R14501 D.n5532 D.t3156 7.099
R14502 D.n5865 D.t1189 7.099
R14503 D.n5851 D.t389 7.099
R14504 D.n5837 D.t2283 7.099
R14505 D.n5823 D.t1124 7.099
R14506 D.n5809 D.t4038 7.099
R14507 D.n5795 D.t2719 7.099
R14508 D.n5781 D.t4353 7.099
R14509 D.n5767 D.t3495 7.099
R14510 D.n5753 D.t382 7.099
R14511 D.n5739 D.t1154 7.099
R14512 D.n5725 D.t3530 7.099
R14513 D.n5711 D.t4488 7.099
R14514 D.n5697 D.t3544 7.099
R14515 D.n5683 D.t3560 7.099
R14516 D.n5669 D.t983 7.099
R14517 D.n5655 D.t299 7.099
R14518 D.n5641 D.t2611 7.099
R14519 D.n5627 D.t4446 7.099
R14520 D.n5613 D.t2327 7.099
R14521 D.n5599 D.t1644 7.099
R14522 D.n5585 D.t230 7.099
R14523 D.n5571 D.t1302 7.099
R14524 D.n5889 D.t1898 7.099
R14525 D.n5905 D.t3647 7.099
R14526 D.n5880 D.t4315 7.099
R14527 D.n6185 D.t3548 7.099
R14528 D.n6171 D.t3862 7.099
R14529 D.n6157 D.t2134 7.099
R14530 D.n6143 D.t2406 7.099
R14531 D.n6129 D.t1224 7.099
R14532 D.n6115 D.t1252 7.099
R14533 D.n6101 D.t4219 7.099
R14534 D.n6087 D.t1300 7.099
R14535 D.n6073 D.t1907 7.099
R14536 D.n6059 D.t2636 7.099
R14537 D.n6045 D.t352 7.099
R14538 D.n6031 D.t190 7.099
R14539 D.n6017 D.t3064 7.099
R14540 D.n6003 D.t3542 7.099
R14541 D.n5989 D.t123 7.099
R14542 D.n5975 D.t512 7.099
R14543 D.n5961 D.t4024 7.099
R14544 D.n5947 D.t2207 7.099
R14545 D.n5933 D.t2714 7.099
R14546 D.n5919 D.t2961 7.099
R14547 D.n6209 D.t4182 7.099
R14548 D.n6225 D.t4175 7.099
R14549 D.n6200 D.t3744 7.099
R14550 D.n6477 D.t3093 7.099
R14551 D.n6463 D.t2989 7.099
R14552 D.n6449 D.t2498 7.099
R14553 D.n6435 D.t3371 7.099
R14554 D.n6421 D.t1639 7.099
R14555 D.n6407 D.t290 7.099
R14556 D.n6393 D.t4012 7.099
R14557 D.n6379 D.t2696 7.099
R14558 D.n6365 D.t3173 7.099
R14559 D.n6351 D.t816 7.099
R14560 D.n6337 D.t2664 7.099
R14561 D.n6323 D.t4372 7.099
R14562 D.n6309 D.t1060 7.099
R14563 D.n6295 D.t3686 7.099
R14564 D.n6281 D.t1166 7.099
R14565 D.n6267 D.t2386 7.099
R14566 D.n6253 D.t347 7.099
R14567 D.n6239 D.t153 7.099
R14568 D.n6501 D.t2253 7.099
R14569 D.n6517 D.t1942 7.099
R14570 D.n6492 D.t80 7.099
R14571 D.n6741 D.t4226 7.099
R14572 D.n6727 D.t3445 7.099
R14573 D.n6713 D.t3832 7.099
R14574 D.n6699 D.t2832 7.099
R14575 D.n6685 D.t2108 7.099
R14576 D.n6671 D.t250 7.099
R14577 D.n6657 D.t113 7.099
R14578 D.n6643 D.t1843 7.099
R14579 D.n6629 D.t3659 7.099
R14580 D.n6615 D.t1279 7.099
R14581 D.n6601 D.t3048 7.099
R14582 D.n6587 D.t3324 7.099
R14583 D.n6573 D.t950 7.099
R14584 D.n6559 D.t2862 7.099
R14585 D.n6545 D.t1631 7.099
R14586 D.n6531 D.t3179 7.099
R14587 D.n6765 D.t3308 7.099
R14588 D.n6781 D.t1603 7.099
R14589 D.n6756 D.t3798 7.099
R14590 D.n6977 D.t4222 7.099
R14591 D.n6963 D.t1305 7.099
R14592 D.n6949 D.t2804 7.099
R14593 D.n6935 D.t4301 7.099
R14594 D.n6921 D.t2475 7.099
R14595 D.n6907 D.t239 7.099
R14596 D.n6893 D.t1515 7.099
R14597 D.n6879 D.t55 7.099
R14598 D.n6865 D.t3872 7.099
R14599 D.n6851 D.t3294 7.099
R14600 D.n6837 D.t778 7.099
R14601 D.n6823 D.t122 7.099
R14602 D.n6809 D.t3118 7.099
R14603 D.n6795 D.t4341 7.099
R14604 D.n7001 D.t3342 7.099
R14605 D.n7017 D.t2860 7.099
R14606 D.n6992 D.t2251 7.099
R14607 D.n7185 D.t1550 7.099
R14608 D.n7171 D.t3295 7.099
R14609 D.n7157 D.t4199 7.099
R14610 D.n7143 D.t4400 7.099
R14611 D.n7129 D.t3698 7.099
R14612 D.n7115 D.t449 7.099
R14613 D.n7101 D.t3913 7.099
R14614 D.n7087 D.t151 7.099
R14615 D.n7073 D.t3775 7.099
R14616 D.n7059 D.t2350 7.099
R14617 D.n7045 D.t3539 7.099
R14618 D.n7031 D.t482 7.099
R14619 D.n7209 D.t3623 7.099
R14620 D.n7225 D.t3632 7.099
R14621 D.n7200 D.t464 7.099
R14622 D.n7365 D.t2209 7.099
R14623 D.n7351 D.t3750 7.099
R14624 D.n7337 D.t4120 7.099
R14625 D.n7323 D.t3357 7.099
R14626 D.n7309 D.t1958 7.099
R14627 D.n7295 D.t3845 7.099
R14628 D.n7281 D.t1306 7.099
R14629 D.n7267 D.t87 7.099
R14630 D.n7253 D.t3605 7.099
R14631 D.n7239 D.t1413 7.099
R14632 D.n7389 D.t3243 7.099
R14633 D.n7405 D.t4483 7.099
R14634 D.n7380 D.t3922 7.099
R14635 D.n7517 D.t1971 7.099
R14636 D.n7503 D.t2560 7.099
R14637 D.n7489 D.t3379 7.099
R14638 D.n7475 D.t3113 7.099
R14639 D.n7461 D.t873 7.099
R14640 D.n7447 D.t1540 7.099
R14641 D.n7433 D.t1143 7.099
R14642 D.n7419 D.t2306 7.099
R14643 D.n7541 D.t3527 7.099
R14644 D.n7557 D.t626 7.099
R14645 D.n7532 D.t3499 7.099
R14646 D.n7641 D.t3791 7.099
R14647 D.n7627 D.t398 7.099
R14648 D.n7613 D.t3452 7.099
R14649 D.n7599 D.t4421 7.099
R14650 D.n7585 D.t3926 7.099
R14651 D.n7571 D.t2570 7.099
R14652 D.n7665 D.t4332 7.099
R14653 D.n7681 D.t2992 7.099
R14654 D.n7656 D.t1069 7.099
R14655 D.n7737 D.t1707 7.099
R14656 D.n7723 D.t1011 7.099
R14657 D.n7709 D.t3589 7.099
R14658 D.n7695 D.t1043 7.099
R14659 D.n7760 D.t2723 7.099
R14660 D.n7776 D.t35 7.099
R14661 D.n7751 D.t974 7.099
R14662 D.n7804 D.t1255 7.099
R14663 D.n7790 D.t1267 7.099
R14664 D.n454 D.t3731 7.065
R14665 D.n7821 D.t1739 7.065
R14666 D.n7893 D.t3260 7.065
R14667 D.n7977 D.t10 7.065
R14668 D.n13660 D.t138 7.065
R14669 D.n13625 D.t3710 7.065
R14670 D.n12737 D.t3247 7.065
R14671 D.n12702 D.t1934 7.065
R14672 D.n11888 D.t4351 7.065
R14673 D.n11853 D.t4478 7.065
R14674 D.n11125 D.t1391 7.065
R14675 D.n11090 D.t2574 7.065
R14676 D.n10442 D.t2903 7.065
R14677 D.n10407 D.t3105 7.065
R14678 D.n9839 D.t2224 7.065
R14679 D.n9804 D.t4040 7.065
R14680 D.n9310 D.t2572 7.065
R14681 D.n9275 D.t330 7.065
R14682 D.n8867 D.t656 7.065
R14683 D.n8832 D.t439 7.065
R14684 D.n8504 D.t3033 7.065
R14685 D.n8469 D.t470 7.065
R14686 D.n8215 D.t1677 7.065
R14687 D.n8180 D.t4362 7.065
R14688 D.n8012 D.t638 7.065
R14689 D.n503 D.t1505 7.038
R14690 D.n7854 D.t826 7.037
R14691 D.n7818 D.t212 7.037
R14692 D.n7931 D.t3563 7.037
R14693 D.n14091 D.t388 7.037
R14694 D.n13178 D.t2722 7.037
R14695 D.n13121 D.t4179 7.037
R14696 D.n12295 D.t3411 7.037
R14697 D.n12243 D.t1297 7.037
R14698 D.n11491 D.t1207 7.037
R14699 D.n11444 D.t2407 7.037
R14700 D.n10768 D.t2706 7.037
R14701 D.n10725 D.t1979 7.037
R14702 D.n10120 D.t3003 7.037
R14703 D.n10079 D.t2604 7.037
R14704 D.n9557 D.t2266 7.037
R14705 D.n9521 D.t4355 7.037
R14706 D.n9073 D.t2445 7.037
R14707 D.n9042 D.t3283 7.037
R14708 D.n8665 D.t1426 7.037
R14709 D.n8636 D.t1606 7.037
R14710 D.n8342 D.t4198 7.037
R14711 D.n8318 D.t3504 7.037
R14712 D.n8098 D.t1457 7.037
R14713 D.n8079 D.t2645 7.037
R14714 D.n7910 D.t2663 7.037
R14715 D.n514 D.t1896 7.037
R14716 D.n1144 D.t279 7.037
R14717 D.n1743 D.t3166 7.037
R14718 D.n2314 D.t4217 7.037
R14719 D.n2857 D.t2164 7.037
R14720 D.n3373 D.t2071 7.037
R14721 D.n3861 D.t492 7.037
R14722 D.n4321 D.t2126 7.037
R14723 D.n4753 D.t2494 7.037
R14724 D.n5157 D.t1647 7.037
R14725 D.n5533 D.t3482 7.037
R14726 D.n5881 D.t2822 7.037
R14727 D.n6201 D.t3463 7.037
R14728 D.n6493 D.t3792 7.037
R14729 D.n6757 D.t2705 7.037
R14730 D.n6993 D.t1530 7.037
R14731 D.n7201 D.t1266 7.037
R14732 D.n7381 D.t2416 7.037
R14733 D.n7533 D.t73 7.037
R14734 D.n7657 D.t1581 7.037
R14735 D.n7752 D.t280 7.037
R14736 D.n532 D.t1274 7.031
R14737 D.n1159 D.t934 7.031
R14738 D.n1758 D.t766 7.031
R14739 D.n2329 D.t937 7.031
R14740 D.n2872 D.t1642 7.031
R14741 D.n3388 D.t2204 7.031
R14742 D.n3876 D.t2379 7.031
R14743 D.n4336 D.t3096 7.031
R14744 D.n4768 D.t2691 7.031
R14745 D.n5172 D.t2890 7.031
R14746 D.n5548 D.t2534 7.031
R14747 D.n5896 D.t1815 7.031
R14748 D.n6216 D.t550 7.031
R14749 D.n6508 D.t4503 7.031
R14750 D.n6772 D.t1048 7.031
R14751 D.n7008 D.t2843 7.031
R14752 D.n7216 D.t222 7.031
R14753 D.n7396 D.t2436 7.031
R14754 D.n7548 D.t3794 7.031
R14755 D.n7672 D.t552 7.031
R14756 D.n7767 D.t3585 7.031
R14757 D.n7859 D.t202 7.031
R14758 D.n7836 D.t2584 7.007
R14759 D.n7826 D.t140 7.007
R14760 D.n446 D.t569 7.007
R14761 D.n437 D.t3389 7.007
R14762 D.n29 D.t2715 7.007
R14763 D.n7956 D.t681 7.007
R14764 D.n7941 D.t669 7.007
R14765 D.n14060 D.t2628 7.007
R14766 D.n14042 D.t1941 7.007
R14767 D.n14024 D.t216 7.007
R14768 D.n14006 D.t567 7.007
R14769 D.n13988 D.t1719 7.007
R14770 D.n13970 D.t860 7.007
R14771 D.n13952 D.t2298 7.007
R14772 D.n13934 D.t469 7.007
R14773 D.n13916 D.t624 7.007
R14774 D.n13898 D.t3338 7.007
R14775 D.n13880 D.t3619 7.007
R14776 D.n13862 D.t4490 7.007
R14777 D.n13844 D.t1816 7.007
R14778 D.n13826 D.t3347 7.007
R14779 D.n13808 D.t2358 7.007
R14780 D.n13790 D.t704 7.007
R14781 D.n13772 D.t248 7.007
R14782 D.n13754 D.t1303 7.007
R14783 D.n13736 D.t255 7.007
R14784 D.n13718 D.t2310 7.007
R14785 D.n13700 D.t3236 7.007
R14786 D.n13681 D.t3020 7.007
R14787 D.n13692 D.t2121 7.007
R14788 D.n13710 D.t1758 7.007
R14789 D.n13728 D.t2182 7.007
R14790 D.n13746 D.t3701 7.007
R14791 D.n13764 D.t18 7.007
R14792 D.n13782 D.t3888 7.007
R14793 D.n13800 D.t2975 7.007
R14794 D.n13818 D.t478 7.007
R14795 D.n13836 D.t3415 7.007
R14796 D.n13854 D.t4408 7.007
R14797 D.n13872 D.t3547 7.007
R14798 D.n13890 D.t1711 7.007
R14799 D.n13908 D.t4465 7.007
R14800 D.n13926 D.t2162 7.007
R14801 D.n13944 D.t3999 7.007
R14802 D.n13962 D.t1326 7.007
R14803 D.n13980 D.t915 7.007
R14804 D.n13998 D.t648 7.007
R14805 D.n14016 D.t3037 7.007
R14806 D.n14034 D.t3046 7.007
R14807 D.n14052 D.t2857 7.007
R14808 D.n14074 D.t1673 7.007
R14809 D.n13206 D.t479 7.007
R14810 D.n13226 D.t2045 7.007
R14811 D.n13246 D.t700 7.007
R14812 D.n13266 D.t2061 7.007
R14813 D.n13286 D.t4007 7.007
R14814 D.n13306 D.t2562 7.007
R14815 D.n13326 D.t1374 7.007
R14816 D.n13346 D.t706 7.007
R14817 D.n13366 D.t2065 7.007
R14818 D.n13386 D.t1848 7.007
R14819 D.n13406 D.t578 7.007
R14820 D.n13426 D.t2535 7.007
R14821 D.n13446 D.t1280 7.007
R14822 D.n13466 D.t2461 7.007
R14823 D.n13486 D.t1665 7.007
R14824 D.n13506 D.t3006 7.007
R14825 D.n13526 D.t3918 7.007
R14826 D.n13546 D.t1623 7.007
R14827 D.n13566 D.t4493 7.007
R14828 D.n13586 D.t1704 7.007
R14829 D.n13606 D.t855 7.007
R14830 D.n13596 D.t4020 7.007
R14831 D.n13576 D.t3421 7.007
R14832 D.n13556 D.t65 7.007
R14833 D.n13536 D.t1383 7.007
R14834 D.n13516 D.t2866 7.007
R14835 D.n13496 D.t1403 7.007
R14836 D.n13476 D.t2255 7.007
R14837 D.n13456 D.t4133 7.007
R14838 D.n13436 D.t4075 7.007
R14839 D.n13416 D.t461 7.007
R14840 D.n13396 D.t3940 7.007
R14841 D.n13376 D.t1731 7.007
R14842 D.n13356 D.t1595 7.007
R14843 D.n13336 D.t1614 7.007
R14844 D.n13316 D.t845 7.007
R14845 D.n13296 D.t2598 7.007
R14846 D.n13276 D.t2758 7.007
R14847 D.n13256 D.t960 7.007
R14848 D.n13236 D.t1963 7.007
R14849 D.n13216 D.t3827 7.007
R14850 D.n13191 D.t3598 7.007
R14851 D.n13097 D.t2803 7.007
R14852 D.n13079 D.t632 7.007
R14853 D.n13061 D.t393 7.007
R14854 D.n13043 D.t1565 7.007
R14855 D.n13025 D.t1917 7.007
R14856 D.n13007 D.t1452 7.007
R14857 D.n12989 D.t241 7.007
R14858 D.n12971 D.t727 7.007
R14859 D.n12953 D.t1906 7.007
R14860 D.n12935 D.t1315 7.007
R14861 D.n12917 D.t1327 7.007
R14862 D.n12899 D.t3026 7.007
R14863 D.n12881 D.t2701 7.007
R14864 D.n12863 D.t2020 7.007
R14865 D.n12845 D.t3949 7.007
R14866 D.n12827 D.t3051 7.007
R14867 D.n12809 D.t763 7.007
R14868 D.n12791 D.t466 7.007
R14869 D.n12773 D.t3626 7.007
R14870 D.n12754 D.t2040 7.007
R14871 D.n12765 D.t3086 7.007
R14872 D.n12783 D.t193 7.007
R14873 D.n12801 D.t3740 7.007
R14874 D.n12819 D.t1482 7.007
R14875 D.n12837 D.t2369 7.007
R14876 D.n12855 D.t3835 7.007
R14877 D.n12873 D.t2667 7.007
R14878 D.n12891 D.t4352 7.007
R14879 D.n12909 D.t3779 7.007
R14880 D.n12927 D.t4079 7.007
R14881 D.n12945 D.t2241 7.007
R14882 D.n12963 D.t2030 7.007
R14883 D.n12981 D.t4 7.007
R14884 D.n12999 D.t2340 7.007
R14885 D.n13017 D.t1521 7.007
R14886 D.n13035 D.t353 7.007
R14887 D.n13053 D.t3494 7.007
R14888 D.n13071 D.t3536 7.007
R14889 D.n13089 D.t814 7.007
R14890 D.n13110 D.t417 7.007
R14891 D.n12323 D.t1427 7.007
R14892 D.n12343 D.t3208 7.007
R14893 D.n12363 D.t1672 7.007
R14894 D.n12383 D.t502 7.007
R14895 D.n12403 D.t2577 7.007
R14896 D.n12423 D.t1851 7.007
R14897 D.n12443 D.t317 7.007
R14898 D.n12463 D.t1985 7.007
R14899 D.n12483 D.t531 7.007
R14900 D.n12503 D.t2651 7.007
R14901 D.n12523 D.t1287 7.007
R14902 D.n12543 D.t2629 7.007
R14903 D.n12563 D.t3995 7.007
R14904 D.n12583 D.t1656 7.007
R14905 D.n12603 D.t2480 7.007
R14906 D.n12623 D.t939 7.007
R14907 D.n12643 D.t3024 7.007
R14908 D.n12663 D.t530 7.007
R14909 D.n12683 D.t3013 7.007
R14910 D.n12673 D.t4055 7.007
R14911 D.n12653 D.t2879 7.007
R14912 D.n12633 D.t1486 7.007
R14913 D.n12613 D.t488 7.007
R14914 D.n12593 D.t2563 7.007
R14915 D.n12573 D.t3901 7.007
R14916 D.n12553 D.t2798 7.007
R14917 D.n12533 D.t1920 7.007
R14918 D.n12513 D.t683 7.007
R14919 D.n12493 D.t2206 7.007
R14920 D.n12473 D.t2151 7.007
R14921 D.n12453 D.t3991 7.007
R14922 D.n12433 D.t2046 7.007
R14923 D.n12413 D.t49 7.007
R14924 D.n12393 D.t425 7.007
R14925 D.n12373 D.t3546 7.007
R14926 D.n12353 D.t3483 7.007
R14927 D.n12333 D.t3305 7.007
R14928 D.n12308 D.t497 7.007
R14929 D.n12212 D.t3891 7.007
R14930 D.n12194 D.t3893 7.007
R14931 D.n12176 D.t58 7.007
R14932 D.n12158 D.t2053 7.007
R14933 D.n12140 D.t3996 7.007
R14934 D.n12122 D.t2557 7.007
R14935 D.n12104 D.t3899 7.007
R14936 D.n12086 D.t64 7.007
R14937 D.n12068 D.t236 7.007
R14938 D.n12050 D.t1761 7.007
R14939 D.n12032 D.t1102 7.007
R14940 D.n12014 D.t918 7.007
R14941 D.n11996 D.t3658 7.007
R14942 D.n11978 D.t3217 7.007
R14943 D.n11960 D.t2113 7.007
R14944 D.n11942 D.t1310 7.007
R14945 D.n11924 D.t3158 7.007
R14946 D.n11905 D.t3344 7.007
R14947 D.n11916 D.t1873 7.007
R14948 D.n11934 D.t2417 7.007
R14949 D.n11952 D.t1246 7.007
R14950 D.n11970 D.t3467 7.007
R14951 D.n11988 D.t2983 7.007
R14952 D.n12006 D.t3391 7.007
R14953 D.n12024 D.t2365 7.007
R14954 D.n12042 D.t2653 7.007
R14955 D.n12060 D.t1879 7.007
R14956 D.n12078 D.t1643 7.007
R14957 D.n12096 D.t800 7.007
R14958 D.n12114 D.t891 7.007
R14959 D.n12132 D.t952 7.007
R14960 D.n12150 D.t506 7.007
R14961 D.n12168 D.t3515 7.007
R14962 D.n12186 D.t3958 7.007
R14963 D.n12204 D.t2005 7.007
R14964 D.n12226 D.t3677 7.007
R14965 D.n11514 D.t21 7.007
R14966 D.n11534 D.t1528 7.007
R14967 D.n11554 D.t946 7.007
R14968 D.n11574 D.t921 7.007
R14969 D.n11594 D.t1612 7.007
R14970 D.n11614 D.t1435 7.007
R14971 D.n11634 D.t629 7.007
R14972 D.n11654 D.t3742 7.007
R14973 D.n11674 D.t4229 7.007
R14974 D.n11694 D.t2674 7.007
R14975 D.n11714 D.t1519 7.007
R14976 D.n11734 D.t203 7.007
R14977 D.n11754 D.t2836 7.007
R14978 D.n11774 D.t4015 7.007
R14979 D.n11794 D.t338 7.007
R14980 D.n11814 D.t2219 7.007
R14981 D.n11834 D.t2150 7.007
R14982 D.n11824 D.t247 7.007
R14983 D.n11804 D.t165 7.007
R14984 D.n11784 D.t4152 7.007
R14985 D.n11764 D.t3863 7.007
R14986 D.n11744 D.t2409 7.007
R14987 D.n11724 D.t979 7.007
R14988 D.n11704 D.t2196 7.007
R14989 D.n11684 D.t3538 7.007
R14990 D.n11664 D.t33 7.007
R14991 D.n11644 D.t954 7.007
R14992 D.n11624 D.t331 7.007
R14993 D.n11604 D.t874 7.007
R14994 D.n11584 D.t1546 7.007
R14995 D.n11564 D.t1084 7.007
R14996 D.n11544 D.t3799 7.007
R14997 D.n11524 D.t4399 7.007
R14998 D.n11501 D.t2742 7.007
R14999 D.n11413 D.t4414 7.007
R15000 D.n11395 D.t296 7.007
R15001 D.n11377 D.t1582 7.007
R15002 D.n11359 D.t2334 7.007
R15003 D.n11341 D.t6 7.007
R15004 D.n11323 D.t1828 7.007
R15005 D.n11305 D.t2036 7.007
R15006 D.n11287 D.t2487 7.007
R15007 D.n11269 D.t598 7.007
R15008 D.n11251 D.t424 7.007
R15009 D.n11233 D.t3214 7.007
R15010 D.n11215 D.t218 7.007
R15011 D.n11197 D.t1925 7.007
R15012 D.n11179 D.t4324 7.007
R15013 D.n11161 D.t1223 7.007
R15014 D.n11142 D.t1749 7.007
R15015 D.n11153 D.t4388 7.007
R15016 D.n11171 D.t2779 7.007
R15017 D.n11189 D.t815 7.007
R15018 D.n11207 D.t1127 7.007
R15019 D.n11225 D.t4469 7.007
R15020 D.n11243 D.t4077 7.007
R15021 D.n11261 D.t4258 7.007
R15022 D.n11279 D.t4325 7.007
R15023 D.n11297 D.t4193 7.007
R15024 D.n11315 D.t764 7.007
R15025 D.n11333 D.t1695 7.007
R15026 D.n11351 D.t416 7.007
R15027 D.n11369 D.t1038 7.007
R15028 D.n11387 D.t3449 7.007
R15029 D.n11405 D.t3446 7.007
R15030 D.n11427 D.t1648 7.007
R15031 D.n10791 D.t1968 7.007
R15032 D.n10811 D.t426 7.007
R15033 D.n10831 D.t1701 7.007
R15034 D.n10851 D.t777 7.007
R15035 D.n10871 D.t3988 7.007
R15036 D.n10891 D.t565 7.007
R15037 D.n10911 D.t3088 7.007
R15038 D.n10931 D.t2640 7.007
R15039 D.n10951 D.t313 7.007
R15040 D.n10971 D.t4128 7.007
R15041 D.n10991 D.t305 7.007
R15042 D.n11011 D.t460 7.007
R15043 D.n11031 D.t383 7.007
R15044 D.n11051 D.t2624 7.007
R15045 D.n11071 D.t4406 7.007
R15046 D.n11061 D.t333 7.007
R15047 D.n11041 D.t2635 7.007
R15048 D.n11021 D.t195 7.007
R15049 D.n11001 D.t3571 7.007
R15050 D.n10981 D.t1598 7.007
R15051 D.n10961 D.t784 7.007
R15052 D.n10941 D.t818 7.007
R15053 D.n10921 D.t1894 7.007
R15054 D.n10901 D.t2489 7.007
R15055 D.n10881 D.t941 7.007
R15056 D.n10861 D.t534 7.007
R15057 D.n10841 D.t3241 7.007
R15058 D.n10821 D.t4051 7.007
R15059 D.n10801 D.t3368 7.007
R15060 D.n10778 D.t1781 7.007
R15061 D.n10694 D.t4127 7.007
R15062 D.n10676 D.t507 7.007
R15063 D.n10658 D.t953 7.007
R15064 D.n10640 D.t888 7.007
R15065 D.n10622 D.t4194 7.007
R15066 D.n10604 D.t4172 7.007
R15067 D.n10586 D.t1674 7.007
R15068 D.n10568 D.t3581 7.007
R15069 D.n10550 D.t4195 7.007
R15070 D.n10532 D.t2787 7.007
R15071 D.n10514 D.t1373 7.007
R15072 D.n10496 D.t11 7.007
R15073 D.n10478 D.t3528 7.007
R15074 D.n10459 D.t1900 7.007
R15075 D.n10470 D.t327 7.007
R15076 D.n10488 D.t4487 7.007
R15077 D.n10506 D.t3561 7.007
R15078 D.n10524 D.t3849 7.007
R15079 D.n10542 D.t2549 7.007
R15080 D.n10560 D.t1788 7.007
R15081 D.n10578 D.t270 7.007
R15082 D.n10596 D.t2650 7.007
R15083 D.n10614 D.t2736 7.007
R15084 D.n10632 D.t1245 7.007
R15085 D.n10650 D.t1256 7.007
R15086 D.n10668 D.t3636 7.007
R15087 D.n10686 D.t2216 7.007
R15088 D.n10708 D.t927 7.007
R15089 D.n10148 D.t1624 7.007
R15090 D.n10168 D.t1237 7.007
R15091 D.n10188 D.t875 7.007
R15092 D.n10208 D.t1229 7.007
R15093 D.n10228 D.t3490 7.007
R15094 D.n10248 D.t892 7.007
R15095 D.n10268 D.t1840 7.007
R15096 D.n10288 D.t2477 7.007
R15097 D.n10308 D.t867 7.007
R15098 D.n10328 D.t1450 7.007
R15099 D.n10348 D.t3713 7.007
R15100 D.n10368 D.t41 7.007
R15101 D.n10388 D.t167 7.007
R15102 D.n10378 D.t4431 7.007
R15103 D.n10358 D.t725 7.007
R15104 D.n10338 D.t1842 7.007
R15105 D.n10318 D.t1296 7.007
R15106 D.n10298 D.t3691 7.007
R15107 D.n10278 D.t4200 7.007
R15108 D.n10258 D.t3566 7.007
R15109 D.n10238 D.t4221 7.007
R15110 D.n10218 D.t2716 7.007
R15111 D.n10198 D.t3456 7.007
R15112 D.n10178 D.t3219 7.007
R15113 D.n10158 D.t3595 7.007
R15114 D.n10133 D.t287 7.007
R15115 D.n10055 D.t2956 7.007
R15116 D.n10037 D.t799 7.007
R15117 D.n10019 D.t2129 7.007
R15118 D.n10001 D.t292 7.007
R15119 D.n9983 D.t329 7.007
R15120 D.n9965 D.t1145 7.007
R15121 D.n9947 D.t158 7.007
R15122 D.n9929 D.t2262 7.007
R15123 D.n9911 D.t314 7.007
R15124 D.n9893 D.t1471 7.007
R15125 D.n9875 D.t2835 7.007
R15126 D.n9856 D.t4407 7.007
R15127 D.n9867 D.t742 7.007
R15128 D.n9885 D.t1338 7.007
R15129 D.n9903 D.t4336 7.007
R15130 D.n9921 D.t4294 7.007
R15131 D.n9939 D.t4274 7.007
R15132 D.n9957 D.t2481 7.007
R15133 D.n9975 D.t1849 7.007
R15134 D.n9993 D.t524 7.007
R15135 D.n10011 D.t3805 7.007
R15136 D.n10029 D.t4141 7.007
R15137 D.n10047 D.t3927 7.007
R15138 D.n10068 D.t1204 7.007
R15139 D.n9585 D.t2238 7.007
R15140 D.n9605 D.t3187 7.007
R15141 D.n9625 D.t3266 7.007
R15142 D.n9645 D.t3438 7.007
R15143 D.n9665 D.t4257 7.007
R15144 D.n9685 D.t4174 7.007
R15145 D.n9705 D.t3838 7.007
R15146 D.n9725 D.t4044 7.007
R15147 D.n9745 D.t4207 7.007
R15148 D.n9765 D.t2403 7.007
R15149 D.n9785 D.t335 7.007
R15150 D.n9775 D.t2687 7.007
R15151 D.n9755 D.t2002 7.007
R15152 D.n9735 D.t898 7.007
R15153 D.n9715 D.t3182 7.007
R15154 D.n9695 D.t2509 7.007
R15155 D.n9675 D.t174 7.007
R15156 D.n9655 D.t1152 7.007
R15157 D.n9635 D.t3693 7.007
R15158 D.n9615 D.t3178 7.007
R15159 D.n9595 D.t2021 7.007
R15160 D.n9570 D.t57 7.007
R15161 D.n9490 D.t2240 7.007
R15162 D.n9472 D.t1448 7.007
R15163 D.n9454 D.t2464 7.007
R15164 D.n9436 D.t2513 7.007
R15165 D.n9418 D.t2296 7.007
R15166 D.n9400 D.t688 7.007
R15167 D.n9382 D.t1464 7.007
R15168 D.n9364 D.t2471 7.007
R15169 D.n9346 D.t1227 7.007
R15170 D.n9327 D.t328 7.007
R15171 D.n9338 D.t3821 7.007
R15172 D.n9356 D.t196 7.007
R15173 D.n9374 D.t1990 7.007
R15174 D.n9392 D.t1057 7.007
R15175 D.n9410 D.t1421 7.007
R15176 D.n9428 D.t2731 7.007
R15177 D.n9446 D.t2876 7.007
R15178 D.n9464 D.t2851 7.007
R15179 D.n9482 D.t2898 7.007
R15180 D.n9504 D.t1096 7.007
R15181 D.n9096 D.t4236 7.007
R15182 D.n9116 D.t2704 7.007
R15183 D.n9136 D.t1469 7.007
R15184 D.n9156 D.t1757 7.007
R15185 D.n9176 D.t2083 7.007
R15186 D.n9196 D.t827 7.007
R15187 D.n9216 D.t2759 7.007
R15188 D.n9236 D.t2075 7.007
R15189 D.n9256 D.t3049 7.007
R15190 D.n9246 D.t1806 7.007
R15191 D.n9226 D.t4233 7.007
R15192 D.n9206 D.t3469 7.007
R15193 D.n9186 D.t2848 7.007
R15194 D.n9166 D.t2613 7.007
R15195 D.n9146 D.t223 7.007
R15196 D.n9126 D.t1070 7.007
R15197 D.n9106 D.t284 7.007
R15198 D.n9083 D.t3457 7.007
R15199 D.n9011 D.t2630 7.007
R15200 D.n8993 D.t4166 7.007
R15201 D.n8975 D.t3145 7.007
R15202 D.n8957 D.t4092 7.007
R15203 D.n8939 D.t4256 7.007
R15204 D.n8921 D.t2654 7.007
R15205 D.n8903 D.t76 7.007
R15206 D.n8884 D.t2395 7.007
R15207 D.n8895 D.t1709 7.007
R15208 D.n8913 D.t2495 7.007
R15209 D.n8931 D.t1350 7.007
R15210 D.n8949 D.t1331 7.007
R15211 D.n8967 D.t3884 7.007
R15212 D.n8985 D.t3202 7.007
R15213 D.n9003 D.t4384 7.007
R15214 D.n9025 D.t2394 7.007
R15215 D.n8693 D.t3053 7.007
R15216 D.n8713 D.t1416 7.007
R15217 D.n8733 D.t2385 7.007
R15218 D.n8753 D.t2503 7.007
R15219 D.n8773 D.t1715 7.007
R15220 D.n8793 D.t3846 7.007
R15221 D.n8813 D.t2292 7.007
R15222 D.n8803 D.t3023 7.007
R15223 D.n8783 D.t445 7.007
R15224 D.n8763 D.t2622 7.007
R15225 D.n8743 D.t3337 7.007
R15226 D.n8723 D.t256 7.007
R15227 D.n8703 D.t2761 7.007
R15228 D.n8678 D.t3606 7.007
R15229 D.n8612 D.t1027 7.007
R15230 D.n8594 D.t2688 7.007
R15231 D.n8576 D.t1275 7.007
R15232 D.n8558 D.t2671 7.007
R15233 D.n8540 D.t975 7.007
R15234 D.n8521 D.t3061 7.007
R15235 D.n8532 D.t1073 7.007
R15236 D.n8550 D.t3174 7.007
R15237 D.n8568 D.t2727 7.007
R15238 D.n8586 D.t3128 7.007
R15239 D.n8604 D.t2872 7.007
R15240 D.n8625 D.t1282 7.007
R15241 D.n8370 D.t935 7.007
R15242 D.n8390 D.t2660 7.007
R15243 D.n8410 D.t2825 7.007
R15244 D.n8430 D.t3413 7.007
R15245 D.n8450 D.t2453 7.007
R15246 D.n8440 D.t155 7.007
R15247 D.n8420 D.t3804 7.007
R15248 D.n8400 D.t1086 7.007
R15249 D.n8380 D.t1353 7.007
R15250 D.n8355 D.t2069 7.007
R15251 D.n8287 D.t3439 7.007
R15252 D.n8269 D.t994 7.007
R15253 D.n8251 D.t2142 7.007
R15254 D.n8232 D.t2749 7.007
R15255 D.n8243 D.t2944 7.007
R15256 D.n8261 D.t42 7.007
R15257 D.n8279 D.t1883 7.007
R15258 D.n8301 D.t372 7.007
R15259 D.n8121 D.t1897 7.007
R15260 D.n8141 D.t1610 7.007
R15261 D.n8161 D.t2978 7.007
R15262 D.n8151 D.t1710 7.007
R15263 D.n8131 D.t3090 7.007
R15264 D.n8108 D.t2911 7.007
R15265 D.n8048 D.t2188 7.007
R15266 D.n8029 D.t412 7.007
R15267 D.n8040 D.t2717 7.007
R15268 D.n8062 D.t1162 7.007
R15269 D.n51 D.t2924 7.007
R15270 D.n60 D.t3450 7.007
R15271 D.n69 D.t1289 7.007
R15272 D.n78 D.t3068 7.007
R15273 D.n87 D.t269 7.007
R15274 D.n96 D.t850 7.007
R15275 D.n105 D.t2133 7.007
R15276 D.n114 D.t1134 7.007
R15277 D.n123 D.t232 7.007
R15278 D.n132 D.t1895 7.007
R15279 D.n141 D.t1543 7.007
R15280 D.n150 D.t615 7.007
R15281 D.n159 D.t136 7.007
R15282 D.n168 D.t370 7.007
R15283 D.n177 D.t3653 7.007
R15284 D.n186 D.t2821 7.007
R15285 D.n195 D.t3312 7.007
R15286 D.n204 D.t555 7.007
R15287 D.n213 D.t1762 7.007
R15288 D.n222 D.t385 7.007
R15289 D.n231 D.t354 7.007
R15290 D.n240 D.t129 7.007
R15291 D.n249 D.t3148 7.007
R15292 D.n258 D.t4093 7.007
R15293 D.n267 D.t997 7.007
R15294 D.n276 D.t1387 7.007
R15295 D.n285 D.t2273 7.007
R15296 D.n294 D.t1927 7.007
R15297 D.n303 D.t2091 7.007
R15298 D.n312 D.t451 7.007
R15299 D.n321 D.t2533 7.007
R15300 D.n330 D.t903 7.007
R15301 D.n339 D.t761 7.007
R15302 D.n348 D.t665 7.007
R15303 D.n357 D.t1692 7.007
R15304 D.n366 D.t1397 7.007
R15305 D.n375 D.t1536 7.007
R15306 D.n384 D.t3170 7.007
R15307 D.n393 D.t1320 7.007
R15308 D.n402 D.t1091 7.007
R15309 D.n411 D.t262 7.007
R15310 D.n420 D.t1884 7.007
R15311 D.n429 D.t1702 7.007
R15312 D.n530 D.t1760 7.007
R15313 D.n522 D.t3226 7.007
R15314 D.n538 D.t2809 7.007
R15315 D.n1126 D.t1077 7.007
R15316 D.n1112 D.t2932 7.007
R15317 D.n1098 D.t175 7.007
R15318 D.n1084 D.t1344 7.007
R15319 D.n1070 D.t3234 7.007
R15320 D.n1056 D.t1080 7.007
R15321 D.n1042 D.t3674 7.007
R15322 D.n1028 D.t584 7.007
R15323 D.n1014 D.t2443 7.007
R15324 D.n1000 D.t2520 7.007
R15325 D.n986 D.t278 7.007
R15326 D.n972 D.t1111 7.007
R15327 D.n958 D.t961 7.007
R15328 D.n944 D.t1752 7.007
R15329 D.n930 D.t120 7.007
R15330 D.n916 D.t793 7.007
R15331 D.n902 D.t4498 7.007
R15332 D.n888 D.t1272 7.007
R15333 D.n874 D.t2791 7.007
R15334 D.n860 D.t2652 7.007
R15335 D.n846 D.t817 7.007
R15336 D.n832 D.t1298 7.007
R15337 D.n818 D.t1125 7.007
R15338 D.n804 D.t4288 7.007
R15339 D.n790 D.t4473 7.007
R15340 D.n776 D.t3609 7.007
R15341 D.n762 D.t3910 7.007
R15342 D.n748 D.t1666 7.007
R15343 D.n734 D.t2528 7.007
R15344 D.n720 D.t1618 7.007
R15345 D.n706 D.t713 7.007
R15346 D.n692 D.t1578 7.007
R15347 D.n678 D.t1683 7.007
R15348 D.n664 D.t2307 7.007
R15349 D.n650 D.t788 7.007
R15350 D.n636 D.t1082 7.007
R15351 D.n622 D.t2726 7.007
R15352 D.n608 D.t668 7.007
R15353 D.n594 D.t3432 7.007
R15354 D.n580 D.t2412 7.007
R15355 D.n566 D.t2797 7.007
R15356 D.n552 D.t2214 7.007
R15357 D.n1157 D.t2673 7.007
R15358 D.n1149 D.t2925 7.007
R15359 D.n1165 D.t173 7.007
R15360 D.n1725 D.t2428 7.007
R15361 D.n1711 D.t2541 7.007
R15362 D.n1697 D.t1186 7.007
R15363 D.n1683 D.t2899 7.007
R15364 D.n1669 D.t3535 7.007
R15365 D.n1655 D.t1247 7.007
R15366 D.n1641 D.t3066 7.007
R15367 D.n1627 D.t2507 7.007
R15368 D.n1613 D.t3410 7.007
R15369 D.n1599 D.t2212 7.007
R15370 D.n1585 D.t3692 7.007
R15371 D.n1571 D.t2148 7.007
R15372 D.n1557 D.t1854 7.007
R15373 D.n1543 D.t732 7.007
R15374 D.n1529 D.t2609 7.007
R15375 D.n1515 D.t2976 7.007
R15376 D.n1501 D.t137 7.007
R15377 D.n1487 D.t1328 7.007
R15378 D.n1473 D.t3689 7.007
R15379 D.n1459 D.t1074 7.007
R15380 D.n1445 D.t3864 7.007
R15381 D.n1431 D.t1007 7.007
R15382 D.n1417 D.t2425 7.007
R15383 D.n1403 D.t756 7.007
R15384 D.n1389 D.t25 7.007
R15385 D.n1375 D.t2889 7.007
R15386 D.n1361 D.t4138 7.007
R15387 D.n1347 D.t545 7.007
R15388 D.n1333 D.t1706 7.007
R15389 D.n1319 D.t738 7.007
R15390 D.n1305 D.t3929 7.007
R15391 D.n1291 D.t209 7.007
R15392 D.n1277 D.t484 7.007
R15393 D.n1263 D.t3133 7.007
R15394 D.n1249 D.t291 7.007
R15395 D.n1235 D.t2841 7.007
R15396 D.n1221 D.t2721 7.007
R15397 D.n1207 D.t3157 7.007
R15398 D.n1193 D.t3745 7.007
R15399 D.n1179 D.t2823 7.007
R15400 D.n1756 D.t1106 7.007
R15401 D.n1748 D.t2849 7.007
R15402 D.n1764 D.t3885 7.007
R15403 D.n2296 D.t1490 7.007
R15404 D.n2282 D.t1579 7.007
R15405 D.n2268 D.t959 7.007
R15406 D.n2254 D.t2880 7.007
R15407 D.n2240 D.t2082 7.007
R15408 D.n2226 D.t3009 7.007
R15409 D.n2212 D.t4308 7.007
R15410 D.n2198 D.t3816 7.007
R15411 D.n2184 D.t3687 7.007
R15412 D.n2170 D.t4402 7.007
R15413 D.n2156 D.t4189 7.007
R15414 D.n2142 D.t825 7.007
R15415 D.n2128 D.t400 7.007
R15416 D.n2114 D.t1253 7.007
R15417 D.n2100 D.t2236 7.007
R15418 D.n2086 D.t2532 7.007
R15419 D.n2072 D.t1222 7.007
R15420 D.n2058 D.t2951 7.007
R15421 D.n2044 D.t4111 7.007
R15422 D.n2030 D.t1177 7.007
R15423 D.n2016 D.t3035 7.007
R15424 D.n2002 D.t301 7.007
R15425 D.n1988 D.t3489 7.007
R15426 D.n1974 D.t2744 7.007
R15427 D.n1960 D.t981 7.007
R15428 D.n1946 D.t3349 7.007
R15429 D.n1932 D.t2200 7.007
R15430 D.n1918 D.t2198 7.007
R15431 D.n1904 D.t206 7.007
R15432 D.n1890 D.t4034 7.007
R15433 D.n1876 D.t1345 7.007
R15434 D.n1862 D.t1600 7.007
R15435 D.n1848 D.t2756 7.007
R15436 D.n1834 D.t3931 7.007
R15437 D.n1820 D.t2438 7.007
R15438 D.n1806 D.t257 7.007
R15439 D.n1792 D.t1400 7.007
R15440 D.n1778 D.t1651 7.007
R15441 D.n2327 D.t3970 7.007
R15442 D.n2319 D.t1889 7.007
R15443 D.n2335 D.t2655 7.007
R15444 D.n2839 D.t666 7.007
R15445 D.n2825 D.t836 7.007
R15446 D.n2811 D.t2396 7.007
R15447 D.n2797 D.t922 7.007
R15448 D.n2783 D.t595 7.007
R15449 D.n2769 D.t2963 7.007
R15450 D.n2755 D.t4154 7.007
R15451 D.n2741 D.t3038 7.007
R15452 D.n2727 D.t2846 7.007
R15453 D.n2713 D.t3986 7.007
R15454 D.n2699 D.t2163 7.007
R15455 D.n2685 D.t3348 7.007
R15456 D.n2671 D.t3129 7.007
R15457 D.n2657 D.t1585 7.007
R15458 D.n2643 D.t2502 7.007
R15459 D.n2629 D.t1529 7.007
R15460 D.n2615 D.t841 7.007
R15461 D.n2601 D.t2984 7.007
R15462 D.n2587 D.t3201 7.007
R15463 D.n2573 D.t391 7.007
R15464 D.n2559 D.t4317 7.007
R15465 D.n2545 D.t2451 7.007
R15466 D.n2531 D.t3387 7.007
R15467 D.n2517 D.t1178 7.007
R15468 D.n2503 D.t2374 7.007
R15469 D.n2489 D.t604 7.007
R15470 D.n2475 D.t2648 7.007
R15471 D.n2461 D.t2138 7.007
R15472 D.n2447 D.t2544 7.007
R15473 D.n2433 D.t2143 7.007
R15474 D.n2419 D.t3839 7.007
R15475 D.n2405 D.t993 7.007
R15476 D.n2391 D.t2868 7.007
R15477 D.n2377 D.t3553 7.007
R15478 D.n2363 D.t2917 7.007
R15479 D.n2349 D.t1095 7.007
R15480 D.n2870 D.t2710 7.007
R15481 D.n2862 D.t4411 7.007
R15482 D.n2878 D.t0 7.007
R15483 D.n3354 D.t3164 7.007
R15484 D.n3340 D.t1826 7.007
R15485 D.n3326 D.t1456 7.007
R15486 D.n3312 D.t1215 7.007
R15487 D.n3298 D.t3335 7.007
R15488 D.n3284 D.t776 7.007
R15489 D.n3270 D.t332 7.007
R15490 D.n3256 D.t4224 7.007
R15491 D.n3242 D.t4313 7.007
R15492 D.n3228 D.t3112 7.007
R15493 D.n3214 D.t2765 7.007
R15494 D.n3200 D.t546 7.007
R15495 D.n3186 D.t4261 7.007
R15496 D.n3172 D.t1830 7.007
R15497 D.n3158 D.t3946 7.007
R15498 D.n3144 D.t1230 7.007
R15499 D.n3130 D.t2389 7.007
R15500 D.n3116 D.t2059 7.007
R15501 D.n3102 D.t643 7.007
R15502 D.n3088 D.t2934 7.007
R15503 D.n3074 D.t3326 7.007
R15504 D.n3060 D.t942 7.007
R15505 D.n3046 D.t2792 7.007
R15506 D.n3032 D.t670 7.007
R15507 D.n3018 D.t1924 7.007
R15508 D.n3004 D.t2302 7.007
R15509 D.n2990 D.t2226 7.007
R15510 D.n2976 D.t3476 7.007
R15511 D.n2962 D.t378 7.007
R15512 D.n2948 D.t4459 7.007
R15513 D.n2934 D.t116 7.007
R15514 D.n2920 D.t4427 7.007
R15515 D.n2906 D.t323 7.007
R15516 D.n2892 D.t3267 7.007
R15517 D.n3386 D.t2618 7.007
R15518 D.n3378 D.t4094 7.007
R15519 D.n3394 D.t1062 7.007
R15520 D.n3842 D.t4158 7.007
R15521 D.n3828 D.t1773 7.007
R15522 D.n3814 D.t1434 7.007
R15523 D.n3800 D.t5 7.007
R15524 D.n3786 D.t2351 7.007
R15525 D.n3772 D.t3906 7.007
R15526 D.n3758 D.t995 7.007
R15527 D.n3744 D.t2864 7.007
R15528 D.n3730 D.t4160 7.007
R15529 D.n3716 D.t4499 7.007
R15530 D.n3702 D.t163 7.007
R15531 D.n3688 D.t3519 7.007
R15532 D.n3674 D.t4318 7.007
R15533 D.n3660 D.t3255 7.007
R15534 D.n3646 D.t2935 7.007
R15535 D.n3632 D.t234 7.007
R15536 D.n3618 D.t1442 7.007
R15537 D.n3604 D.t847 7.007
R15538 D.n3590 D.t3471 7.007
R15539 D.n3576 D.t770 7.007
R15540 D.n3562 D.t2596 7.007
R15541 D.n3548 D.t2774 7.007
R15542 D.n3534 D.t4227 7.007
R15543 D.n3520 D.t1120 7.007
R15544 D.n3506 D.t3718 7.007
R15545 D.n3492 D.t2907 7.007
R15546 D.n3478 D.t3290 7.007
R15547 D.n3464 D.t2096 7.007
R15548 D.n3450 D.t686 7.007
R15549 D.n3436 D.t1931 7.007
R15550 D.n3422 D.t281 7.007
R15551 D.n3408 D.t2690 7.007
R15552 D.n3874 D.t3141 7.007
R15553 D.n3866 D.t1415 7.007
R15554 D.n3882 D.t3140 7.007
R15555 D.n4302 D.t1370 7.007
R15556 D.n4288 D.t1369 7.007
R15557 D.n4274 D.t2861 7.007
R15558 D.n4260 D.t1398 7.007
R15559 D.n4246 D.t1422 7.007
R15560 D.n4232 D.t2202 7.007
R15561 D.n4218 D.t1756 7.007
R15562 D.n4204 D.t4445 7.007
R15563 D.n4190 D.t790 7.007
R15564 D.n4176 D.t369 7.007
R15565 D.n4162 D.t2217 7.007
R15566 D.n4148 D.t4097 7.007
R15567 D.n4134 D.t2013 7.007
R15568 D.n4120 D.t719 7.007
R15569 D.n4106 D.t4234 7.007
R15570 D.n4092 D.t1479 7.007
R15571 D.n4078 D.t1433 7.007
R15572 D.n4064 D.t1776 7.007
R15573 D.n4050 D.t2269 7.007
R15574 D.n4036 D.t3475 7.007
R15575 D.n4022 D.t4132 7.007
R15576 D.n4008 D.t2913 7.007
R15577 D.n3994 D.t3259 7.007
R15578 D.n3980 D.t37 7.007
R15579 D.n3966 D.t3941 7.007
R15580 D.n3952 D.t62 7.007
R15581 D.n3938 D.t4156 7.007
R15582 D.n3924 D.t2505 7.007
R15583 D.n3910 D.t2339 7.007
R15584 D.n3896 D.t695 7.007
R15585 D.n4334 D.t245 7.007
R15586 D.n4326 D.t4451 7.007
R15587 D.n4342 D.t1138 7.007
R15588 D.n4734 D.t1362 7.007
R15589 D.n4720 D.t4447 7.007
R15590 D.n4706 D.t3453 7.007
R15591 D.n4692 D.t2377 7.007
R15592 D.n4678 D.t2147 7.007
R15593 D.n4664 D.t2685 7.007
R15594 D.n4650 D.t610 7.007
R15595 D.n4636 D.t3356 7.007
R15596 D.n4622 D.t1588 7.007
R15597 D.n4608 D.t1139 7.007
R15598 D.n4594 D.t527 7.007
R15599 D.n4580 D.t4480 7.007
R15600 D.n4566 D.t3177 7.007
R15601 D.n4552 D.t4088 7.007
R15602 D.n4538 D.t4081 7.007
R15603 D.n4524 D.t1645 7.007
R15604 D.n4510 D.t2901 7.007
R15605 D.n4496 D.t1332 7.007
R15606 D.n4482 D.t1407 7.007
R15607 D.n4468 D.t243 7.007
R15608 D.n4454 D.t3251 7.007
R15609 D.n4440 D.t1864 7.007
R15610 D.n4426 D.t3921 7.007
R15611 D.n4412 D.t516 7.007
R15612 D.n4398 D.t432 7.007
R15613 D.n4384 D.t147 7.007
R15614 D.n4370 D.t2043 7.007
R15615 D.n4356 D.t2265 7.007
R15616 D.n4766 D.t634 7.007
R15617 D.n4758 D.t1748 7.007
R15618 D.n4774 D.t986 7.007
R15619 D.n5138 D.t2146 7.007
R15620 D.n5124 D.t3095 7.007
R15621 D.n5110 D.t4390 7.007
R15622 D.n5096 D.t1713 7.007
R15623 D.n5082 D.t823 7.007
R15624 D.n5068 D.t2232 7.007
R15625 D.n5054 D.t1079 7.007
R15626 D.n5040 D.t2737 7.007
R15627 D.n5026 D.t1769 7.007
R15628 D.n5012 D.t2249 7.007
R15629 D.n4998 D.t787 7.007
R15630 D.n4984 D.t315 7.007
R15631 D.n4970 D.t1992 7.007
R15632 D.n4956 D.t2208 7.007
R15633 D.n4942 D.t1115 7.007
R15634 D.n4928 D.t2909 7.007
R15635 D.n4914 D.t3708 7.007
R15636 D.n4900 D.t1901 7.007
R15637 D.n4886 D.t3397 7.007
R15638 D.n4872 D.t3235 7.007
R15639 D.n4858 D.t355 7.007
R15640 D.n4844 D.t1392 7.007
R15641 D.n4830 D.t4428 7.007
R15642 D.n4816 D.t435 7.007
R15643 D.n4802 D.t3607 7.007
R15644 D.n4788 D.t82 7.007
R15645 D.n5170 D.t2001 7.007
R15646 D.n5162 D.t345 7.007
R15647 D.n5178 D.t2981 7.007
R15648 D.n5514 D.t1291 7.007
R15649 D.n5500 D.t4350 7.007
R15650 D.n5486 D.t2546 7.007
R15651 D.n5472 D.t3730 7.007
R15652 D.n5458 D.t2786 7.007
R15653 D.n5444 D.t2355 7.007
R15654 D.n5430 D.t1249 7.007
R15655 D.n5416 D.t1946 7.007
R15656 D.n5402 D.t304 7.007
R15657 D.n5388 D.t3376 7.007
R15658 D.n5374 D.t3481 7.007
R15659 D.n5360 D.t2387 7.007
R15660 D.n5346 D.t3809 7.007
R15661 D.n5332 D.t1000 7.007
R15662 D.n5318 D.t2755 7.007
R15663 D.n5304 D.t3972 7.007
R15664 D.n5290 D.t796 7.007
R15665 D.n5276 D.t682 7.007
R15666 D.n5262 D.t673 7.007
R15667 D.n5248 D.t2176 7.007
R15668 D.n5234 D.t1009 7.007
R15669 D.n5220 D.t3700 7.007
R15670 D.n5206 D.t753 7.007
R15671 D.n5192 D.t1802 7.007
R15672 D.n5546 D.t4425 7.007
R15673 D.n5538 D.t802 7.007
R15674 D.n5554 D.t3175 7.007
R15675 D.n5862 D.t1881 7.007
R15676 D.n5848 D.t4083 7.007
R15677 D.n5834 D.t2011 7.007
R15678 D.n5820 D.t3010 7.007
R15679 D.n5806 D.t3099 7.007
R15680 D.n5792 D.t442 7.007
R15681 D.n5778 D.t730 7.007
R15682 D.n5764 D.t1804 7.007
R15683 D.n5750 D.t1061 7.007
R15684 D.n5736 D.t3032 7.007
R15685 D.n5722 D.t2939 7.007
R15686 D.n5708 D.t3180 7.007
R15687 D.n5694 D.t908 7.007
R15688 D.n5680 D.t833 7.007
R15689 D.n5666 D.t1957 7.007
R15690 D.n5652 D.t3778 7.007
R15691 D.n5638 D.t455 7.007
R15692 D.n5624 D.t1322 7.007
R15693 D.n5610 D.t1175 7.007
R15694 D.n5596 D.t2119 7.007
R15695 D.n5582 D.t3212 7.007
R15696 D.n5568 D.t4180 7.007
R15697 D.n5894 D.t1022 7.007
R15698 D.n5886 D.t4041 7.007
R15699 D.n5902 D.t2220 7.007
R15700 D.n6182 D.t1654 7.007
R15701 D.n6168 D.t1587 7.007
R15702 D.n6154 D.t1098 7.007
R15703 D.n6140 D.t4369 7.007
R15704 D.n6126 D.t2067 7.007
R15705 D.n6112 D.t3722 7.007
R15706 D.n6098 D.t2921 7.007
R15707 D.n6084 D.t3650 7.007
R15708 D.n6070 D.t967 7.007
R15709 D.n6056 D.t4417 7.007
R15710 D.n6042 D.t3503 7.007
R15711 D.n6028 D.t3309 7.007
R15712 D.n6014 D.t3408 7.007
R15713 D.n6000 D.t3565 7.007
R15714 D.n5986 D.t3447 7.007
R15715 D.n5972 D.t4410 7.007
R15716 D.n5958 D.t3022 7.007
R15717 D.n5944 D.t1235 7.007
R15718 D.n5930 D.t409 7.007
R15719 D.n5916 D.t538 7.007
R15720 D.n6214 D.t473 7.007
R15721 D.n6206 D.t2229 7.007
R15722 D.n6222 D.t4391 7.007
R15723 D.n6474 D.t3435 7.007
R15724 D.n6460 D.t3625 7.007
R15725 D.n6446 D.t1114 7.007
R15726 D.n6432 D.t3855 7.007
R15727 D.n6418 D.t1141 7.007
R15728 D.n6404 D.t4272 7.007
R15729 D.n6390 D.t2830 7.007
R15730 D.n6376 D.t650 7.007
R15731 D.n6362 D.t930 7.007
R15732 D.n6348 D.t3343 7.007
R15733 D.n6334 D.t3790 7.007
R15734 D.n6320 D.t3576 7.007
R15735 D.n6306 D.t1090 7.007
R15736 D.n6292 D.t862 7.007
R15737 D.n6278 D.t1319 7.007
R15738 D.n6264 D.t4273 7.007
R15739 D.n6250 D.t2057 7.007
R15740 D.n6236 D.t3937 7.007
R15741 D.n6506 D.t2818 7.007
R15742 D.n6498 D.t3131 7.007
R15743 D.n6514 D.t601 7.007
R15744 D.n6738 D.t723 7.007
R15745 D.n6724 D.t2575 7.007
R15746 D.n6710 D.t1835 7.007
R15747 D.n6696 D.t3878 7.007
R15748 D.n6682 D.t1195 7.007
R15749 D.n6668 D.t4299 7.007
R15750 D.n6654 D.t2048 7.007
R15751 D.n6640 D.t2893 7.007
R15752 D.n6626 D.t4340 7.007
R15753 D.n6612 D.t3314 7.007
R15754 D.n6598 D.t509 7.007
R15755 D.n6584 D.t1989 7.007
R15756 D.n6570 D.t1487 7.007
R15757 D.n6556 D.t3620 7.007
R15758 D.n6542 D.t489 7.007
R15759 D.n6528 D.t3330 7.007
R15760 D.n6770 D.t1285 7.007
R15761 D.n6762 D.t2923 7.007
R15762 D.n6778 D.t2390 7.007
R15763 D.n6974 D.t3430 7.007
R15764 D.n6960 D.t430 7.007
R15765 D.n6946 D.t3666 7.007
R15766 D.n6932 D.t2290 7.007
R15767 D.n6918 D.t39 7.007
R15768 D.n6904 D.t1592 7.007
R15769 D.n6890 D.t2753 7.007
R15770 D.n6876 D.t228 7.007
R15771 D.n6862 D.t992 7.007
R15772 D.n6848 D.t3162 7.007
R15773 D.n6834 D.t4107 7.007
R15774 D.n6820 D.t619 7.007
R15775 D.n6806 D.t1483 7.007
R15776 D.n6792 D.t318 7.007
R15777 D.n7006 D.t1443 7.007
R15778 D.n6998 D.t2449 7.007
R15779 D.n7014 D.t2965 7.007
R15780 D.n7182 D.t3285 7.007
R15781 D.n7168 D.t4048 7.007
R15782 D.n7154 D.t1596 7.007
R15783 D.n7140 D.t856 7.007
R15784 D.n7126 D.t1431 7.007
R15785 D.n7112 D.t2878 7.007
R15786 D.n7098 D.t3111 7.007
R15787 D.n7084 D.t3645 7.007
R15788 D.n7070 D.t1396 7.007
R15789 D.n7056 D.t3825 7.007
R15790 D.n7042 D.t1384 7.007
R15791 D.n7028 D.t3982 7.007
R15792 D.n7214 D.t3914 7.007
R15793 D.n7206 D.t2895 7.007
R15794 D.n7222 D.t9 7.007
R15795 D.n7362 D.t4466 7.007
R15796 D.n7348 D.t2982 7.007
R15797 D.n7334 D.t2827 7.007
R15798 D.n7320 D.t1304 7.007
R15799 D.n7306 D.t2738 7.007
R15800 D.n7292 D.t4453 7.007
R15801 D.n7278 D.t2183 7.007
R15802 D.n7264 D.t2521 7.007
R15803 D.n7250 D.t3727 7.007
R15804 D.n7236 D.t2556 7.007
R15805 D.n7394 D.t1786 7.007
R15806 D.n7386 D.t89 7.007
R15807 D.n7402 D.t4310 7.007
R15808 D.n7514 D.t1745 7.007
R15809 D.n7500 D.t1630 7.007
R15810 D.n7486 D.t1714 7.007
R15811 D.n7472 D.t2615 7.007
R15812 D.n7458 D.t2346 7.007
R15813 D.n7444 D.t3299 7.007
R15814 D.n7430 D.t2595 7.007
R15815 D.n7416 D.t2657 7.007
R15816 D.n7546 D.t2156 7.007
R15817 D.n7538 D.t2926 7.007
R15818 D.n7554 D.t611 7.007
R15819 D.n7638 D.t4316 7.007
R15820 D.n7624 D.t1121 7.007
R15821 D.n7610 D.t4333 7.007
R15822 D.n7596 D.t1874 7.007
R15823 D.n7582 D.t869 7.007
R15824 D.n7568 D.t2746 7.007
R15825 D.n7670 D.t2263 7.007
R15826 D.n7662 D.t1937 7.007
R15827 D.n7678 D.t3783 7.007
R15828 D.n7734 D.t1126 7.007
R15829 D.n7720 D.t807 7.007
R15830 D.n7706 D.t4368 7.007
R15831 D.n7692 D.t283 7.007
R15832 D.n7765 D.t3079 7.007
R15833 D.n7757 D.t3250 7.007
R15834 D.n7773 D.t3736 7.007
R15835 D.n7801 D.t4082 7.007
R15836 D.n7787 D.t2796 7.007
R15837 D.n7820 D.t2745 7.007
R15838 D.n7857 D.t982 7.007
R15839 D.n531 D.t3774 6.598
R15840 D.n1158 D.t3479 6.598
R15841 D.n1757 D.t2553 6.598
R15842 D.n2328 D.t311 6.598
R15843 D.n2871 D.t392 6.598
R15844 D.n3387 D.t4113 6.598
R15845 D.n3875 D.t880 6.598
R15846 D.n4335 D.t667 6.598
R15847 D.n4767 D.t1686 6.598
R15848 D.n5171 D.t1402 6.598
R15849 D.n5547 D.t3892 6.598
R15850 D.n5895 D.t1671 6.598
R15851 D.n6215 D.t1564 6.598
R15852 D.n6507 D.t4004 6.598
R15853 D.n6771 D.t2098 6.598
R15854 D.n7007 D.t902 6.598
R15855 D.n7215 D.t712 6.598
R15856 D.n7395 D.t879 6.598
R15857 D.n7547 D.t322 6.598
R15858 D.n7671 D.t387 6.598
R15859 D.n7766 D.t4230 6.598
R15860 D.n7858 D.t1473 6.598
R15861 D.n503 D.t443 6.568
R15862 D.n7894 D.t630 6.564
R15863 D.n7978 D.t3624 6.564
R15864 D.n13661 D.t4321 6.564
R15865 D.n13626 D.t1552 6.564
R15866 D.n12738 D.t1137 6.564
R15867 D.n12703 D.t4091 6.564
R15868 D.n11889 D.t3663 6.564
R15869 D.n11854 D.t2997 6.564
R15870 D.n11126 D.t1352 6.564
R15871 D.n11091 D.t575 6.564
R15872 D.n10443 D.t2906 6.564
R15873 D.n10408 D.t3828 6.564
R15874 D.n9840 D.t1547 6.564
R15875 D.n9805 D.t2853 6.564
R15876 D.n9311 D.t2362 6.564
R15877 D.n9276 D.t242 6.564
R15878 D.n8868 D.t1850 6.564
R15879 D.n8833 D.t3788 6.564
R15880 D.n8505 D.t4150 6.564
R15881 D.n8470 D.t1965 6.564
R15882 D.n8216 D.t4119 6.564
R15883 D.n8181 D.t3695 6.564
R15884 D.n8013 D.t1071 6.564
R15885 D.n7822 D.t1507 6.564
R15886 D.n454 D.t697 6.528
R15887 D.n7852 D.t127 6.524
R15888 D.n7819 D.t3961 6.524
R15889 D.n7929 D.t1751 6.524
R15890 D.n14089 D.t2676 6.524
R15891 D.n13179 D.t434 6.524
R15892 D.n13122 D.t2080 6.524
R15893 D.n12296 D.t1523 6.524
R15894 D.n12241 D.t2328 6.524
R15895 D.n11492 D.t878 6.524
R15896 D.n11442 D.t2523 6.524
R15897 D.n10769 D.t1909 6.524
R15898 D.n10723 D.t587 6.524
R15899 D.n10121 D.t2064 6.524
R15900 D.n10080 D.t1904 6.524
R15901 D.n9558 D.t515 6.524
R15902 D.n9519 D.t2056 6.524
R15903 D.n9074 D.t4237 6.524
R15904 D.n9040 D.t457 6.524
R15905 D.n8666 D.t321 6.524
R15906 D.n8637 D.t4202 6.524
R15907 D.n8343 D.t1233 6.524
R15908 D.n8316 D.t298 6.524
R15909 D.n8099 D.t2399 6.524
R15910 D.n8077 D.t198 6.524
R15911 D.n7911 D.t183 6.524
R15912 D.n515 D.t1261 6.524
R15913 D.n1145 D.t1292 6.524
R15914 D.n1744 D.t1839 6.524
R15915 D.n2315 D.t2141 6.524
R15916 D.n2858 D.t3258 6.524
R15917 D.n3374 D.t3431 6.524
R15918 D.n3862 D.t3319 6.524
R15919 D.n4322 D.t4463 6.524
R15920 D.n4754 D.t1766 6.524
R15921 D.n5158 D.t2739 6.524
R15922 D.n5534 D.t371 6.524
R15923 D.n5882 D.t3252 6.524
R15924 D.n6202 D.t2233 6.524
R15925 D.n6494 D.t1629 6.524
R15926 D.n6758 D.t3360 6.524
R15927 D.n6994 D.t3905 6.524
R15928 D.n7202 D.t752 6.524
R15929 D.n7382 D.t2734 6.524
R15930 D.n7534 D.t3165 6.524
R15931 D.n7658 D.t2771 6.524
R15932 D.n7753 D.t709 6.524
R15933 D.n7846 D.n7843 0.344
R15934 D.n3371 D.n3370 0.327
R15935 D.n3859 D.n3858 0.327
R15936 D.n4319 D.n4318 0.327
R15937 D.n4751 D.n4750 0.327
R15938 D.n5155 D.n5154 0.327
R15939 D.n5531 D.n5530 0.327
R15940 D.n5879 D.n5878 0.327
R15941 D.n6199 D.n6198 0.327
R15942 D.n6491 D.n6490 0.327
R15943 D.n6755 D.n6754 0.327
R15944 D.n6991 D.n6990 0.327
R15945 D.n7199 D.n7198 0.327
R15946 D.n7379 D.n7378 0.327
R15947 D.n7531 D.n7530 0.327
R15948 D.n7655 D.n7654 0.327
R15949 D.n508 D.n507 0.31
R15950 D.n7846 D.n7845 0.225
R15951 D.n520 D.n519 0.225
R15952 D.n1147 D.n1146 0.225
R15953 D.n1746 D.n1745 0.225
R15954 D.n2317 D.n2316 0.225
R15955 D.n2860 D.n2859 0.225
R15956 D.n3376 D.n3375 0.225
R15957 D.n3864 D.n3863 0.225
R15958 D.n4324 D.n4323 0.225
R15959 D.n4756 D.n4755 0.225
R15960 D.n5160 D.n5159 0.225
R15961 D.n5536 D.n5535 0.225
R15962 D.n5884 D.n5883 0.225
R15963 D.n6204 D.n6203 0.225
R15964 D.n6496 D.n6495 0.225
R15965 D.n6760 D.n6759 0.225
R15966 D.n6996 D.n6995 0.225
R15967 D.n7204 D.n7203 0.225
R15968 D.n7384 D.n7383 0.225
R15969 D.n7536 D.n7535 0.225
R15970 D.n7660 D.n7659 0.225
R15971 D.n7755 D.n7754 0.225
R15972 D.n7848 D.n7847 0.225
R15973 D.n14080 D.n14079 0.21
R15974 D.n13201 D.n13200 0.21
R15975 D.n13116 D.n13115 0.21
R15976 D.n12318 D.n12317 0.21
R15977 D.n11509 D.n11508 0.21
R15978 D.n10786 D.n10785 0.21
R15979 D.n10143 D.n10142 0.21
R15980 D.n10074 D.n10073 0.21
R15981 D.n9580 D.n9579 0.21
R15982 D.n9091 D.n9090 0.21
R15983 D.n8688 D.n8687 0.21
R15984 D.n8631 D.n8630 0.21
R15985 D.n8365 D.n8364 0.21
R15986 D.n8116 D.n8115 0.21
R15987 D.n7951 D.n7950 0.21
R15988 D.n7920 D.n7919 0.205
R15989 D.n7891 D.n7890 0.192
R15990 D.n7898 D.n7897 0.174
R15991 D.n7922 D.n7921 0.163
R15992 D.n7862 D.n7861 0.144
R15993 D.n7988 D.n7987 0.143
R15994 D.n13679 D.n13645 0.143
R15995 D.n13679 D.n13678 0.143
R15996 D.n13636 D.n13173 0.143
R15997 D.n13636 D.n13635 0.143
R15998 D.n12752 D.n12722 0.143
R15999 D.n12752 D.n12751 0.143
R16000 D.n12713 D.n12290 0.143
R16001 D.n12713 D.n12712 0.143
R16002 D.n11903 D.n11873 0.143
R16003 D.n11903 D.n11902 0.143
R16004 D.n11864 D.n11487 0.143
R16005 D.n11864 D.n11863 0.143
R16006 D.n11140 D.n11110 0.143
R16007 D.n11140 D.n11139 0.143
R16008 D.n11101 D.n10764 0.143
R16009 D.n11101 D.n11100 0.143
R16010 D.n10457 D.n10427 0.143
R16011 D.n10457 D.n10456 0.143
R16012 D.n10418 D.n10115 0.143
R16013 D.n10418 D.n10417 0.143
R16014 D.n9854 D.n9824 0.143
R16015 D.n9854 D.n9853 0.143
R16016 D.n9815 D.n9552 0.143
R16017 D.n9815 D.n9814 0.143
R16018 D.n9325 D.n9295 0.143
R16019 D.n9325 D.n9324 0.143
R16020 D.n9286 D.n9069 0.143
R16021 D.n9286 D.n9285 0.143
R16022 D.n8882 D.n8852 0.143
R16023 D.n8882 D.n8881 0.143
R16024 D.n8843 D.n8660 0.143
R16025 D.n8843 D.n8842 0.143
R16026 D.n8519 D.n8489 0.143
R16027 D.n8519 D.n8518 0.143
R16028 D.n8480 D.n8337 0.143
R16029 D.n8480 D.n8479 0.143
R16030 D.n8230 D.n8200 0.143
R16031 D.n8230 D.n8229 0.143
R16032 D.n8191 D.n8094 0.143
R16033 D.n8191 D.n8190 0.143
R16034 D.n8027 D.n7997 0.143
R16035 D.n8027 D.n8026 0.143
R16036 D.n7988 D.n7923 0.143
R16037 D.n7902 D.n7901 0.143
R16038 D.n11498 D.n11488 0.14
R16039 D.n10775 D.n10765 0.14
R16040 D.n9080 D.n9070 0.14
R16041 D.n8105 D.n8095 0.14
R16042 D.n7900 D.n7898 0.133
R16043 D.n14142 D.n14141 0.133
R16044 D.n13169 D.n13168 0.133
R16045 D.n12286 D.n12285 0.133
R16046 D.n11483 D.n11482 0.133
R16047 D.n10760 D.n10759 0.133
R16048 D.n10111 D.n10110 0.133
R16049 D.n9548 D.n9547 0.133
R16050 D.n9065 D.n9064 0.133
R16051 D.n8656 D.n8655 0.133
R16052 D.n8333 D.n8332 0.133
R16053 D.n8090 D.n8089 0.133
R16054 D.n14086 D.n14083 0.131
R16055 D.n14095 D.n14094 0.131
R16056 D.n12238 D.n12234 0.131
R16057 D.n12247 D.n12246 0.131
R16058 D.n11439 D.n11435 0.131
R16059 D.n11448 D.n11447 0.131
R16060 D.n10720 D.n10716 0.131
R16061 D.n10729 D.n10728 0.131
R16062 D.n9516 D.n9512 0.131
R16063 D.n9525 D.n9524 0.131
R16064 D.n9037 D.n9033 0.131
R16065 D.n9046 D.n9045 0.131
R16066 D.n8313 D.n8309 0.131
R16067 D.n8322 D.n8321 0.131
R16068 D.n8074 D.n8070 0.131
R16069 D.n8083 D.n8082 0.131
R16070 D.n7937 D.n7936 0.123
R16071 D.n13187 D.n13186 0.123
R16072 D.n12304 D.n12303 0.123
R16073 D.n10129 D.n10128 0.123
R16074 D.n9566 D.n9565 0.123
R16075 D.n8674 D.n8673 0.123
R16076 D.n8351 D.n8350 0.123
R16077 D.n13127 D.n13126 0.115
R16078 D.n11496 D.n11495 0.115
R16079 D.n10773 D.n10772 0.115
R16080 D.n10085 D.n10084 0.115
R16081 D.n9078 D.n9077 0.115
R16082 D.n8642 D.n8641 0.115
R16083 D.n8103 D.n8102 0.115
R16084 D.n7862 D.n7850 0.115
R16085 D.n13623 D.n13614 0.113
R16086 D.n12700 D.n12691 0.113
R16087 D.n11851 D.n11842 0.113
R16088 D.n11088 D.n11079 0.113
R16089 D.n10405 D.n10396 0.113
R16090 D.n9802 D.n9793 0.113
R16091 D.n9273 D.n9264 0.113
R16092 D.n8830 D.n8821 0.113
R16093 D.n8467 D.n8458 0.113
R16094 D.n8178 D.n8169 0.113
R16095 D.n7973 D.n7964 0.113
R16096 D.n7883 D.n1141 0.111
R16097 D.n7882 D.n1740 0.111
R16098 D.n7881 D.n2311 0.111
R16099 D.n7880 D.n2854 0.111
R16100 D.n7879 D.n3369 0.111
R16101 D.n7878 D.n3857 0.111
R16102 D.n7877 D.n4317 0.111
R16103 D.n7876 D.n4749 0.111
R16104 D.n7875 D.n5153 0.111
R16105 D.n7874 D.n5529 0.111
R16106 D.n7873 D.n5877 0.111
R16107 D.n7872 D.n6197 0.111
R16108 D.n7871 D.n6489 0.111
R16109 D.n7870 D.n6753 0.111
R16110 D.n7869 D.n6989 0.111
R16111 D.n7868 D.n7197 0.111
R16112 D.n7867 D.n7377 0.111
R16113 D.n7866 D.n7529 0.111
R16114 D.n7865 D.n7653 0.111
R16115 D.n7864 D.n7749 0.111
R16116 D.n7863 D.n7816 0.11
R16117 D.n7938 D.n7925 0.109
R16118 D.n14071 D.n14068 0.109
R16119 D.n13188 D.n13175 0.109
R16120 D.n12305 D.n12292 0.109
R16121 D.n12223 D.n12220 0.109
R16122 D.n11424 D.n11421 0.109
R16123 D.n10705 D.n10702 0.109
R16124 D.n10130 D.n10117 0.109
R16125 D.n9567 D.n9554 0.109
R16126 D.n9501 D.n9498 0.109
R16127 D.n9022 D.n9019 0.109
R16128 D.n8675 D.n8662 0.109
R16129 D.n8352 D.n8339 0.109
R16130 D.n8298 D.n8295 0.109
R16131 D.n8059 D.n8056 0.109
R16132 D.n7887 D.n7885 0.109
R16133 D.n7950 D.n7947 0.109
R16134 D.n13200 D.n13197 0.109
R16135 D.n12317 D.n12314 0.109
R16136 D.n10142 D.n10139 0.109
R16137 D.n9579 D.n9576 0.109
R16138 D.n8687 D.n8684 0.109
R16139 D.n8364 D.n8361 0.109
R16140 D.n13642 D.n13641 0.105
R16141 D.n12719 D.n12718 0.105
R16142 D.n11870 D.n11869 0.105
R16143 D.n11107 D.n11106 0.105
R16144 D.n10424 D.n10423 0.105
R16145 D.n9821 D.n9820 0.105
R16146 D.n9292 D.n9291 0.105
R16147 D.n8849 D.n8848 0.105
R16148 D.n8486 D.n8485 0.105
R16149 D.n8197 D.n8196 0.105
R16150 D.n7994 D.n7993 0.105
R16151 D.n13644 D.n13643 0.105
R16152 D.n12721 D.n12720 0.105
R16153 D.n11872 D.n11871 0.105
R16154 D.n11109 D.n11108 0.105
R16155 D.n10426 D.n10425 0.105
R16156 D.n9823 D.n9822 0.105
R16157 D.n9294 D.n9293 0.105
R16158 D.n8851 D.n8850 0.105
R16159 D.n8488 D.n8487 0.105
R16160 D.n8199 D.n8198 0.105
R16161 D.n7996 D.n7995 0.105
R16162 D.n7928 D.n7927 0.102
R16163 D.n14093 D.n14092 0.102
R16164 D.n14088 D.n14087 0.102
R16165 D.n13181 D.n13180 0.102
R16166 D.n12298 D.n12297 0.102
R16167 D.n12245 D.n12244 0.102
R16168 D.n12240 D.n12239 0.102
R16169 D.n11446 D.n11445 0.102
R16170 D.n11441 D.n11440 0.102
R16171 D.n10727 D.n10726 0.102
R16172 D.n10722 D.n10721 0.102
R16173 D.n10123 D.n10122 0.102
R16174 D.n9560 D.n9559 0.102
R16175 D.n9523 D.n9522 0.102
R16176 D.n9518 D.n9517 0.102
R16177 D.n9044 D.n9043 0.102
R16178 D.n9039 D.n9038 0.102
R16179 D.n8668 D.n8667 0.102
R16180 D.n8345 D.n8344 0.102
R16181 D.n8320 D.n8319 0.102
R16182 D.n8315 D.n8314 0.102
R16183 D.n8081 D.n8080 0.102
R16184 D.n8076 D.n8075 0.102
R16185 D.n7913 D.n7912 0.102
R16186 D.n7919 D.n7904 0.101
R16187 D.n13666 D.n13665 0.096
R16188 D.n518 D.n517 0.092
R16189 D.n10 D.n9 0.092
R16190 D.n508 D.n505 0.091
R16191 D.n7884 D.n511 0.085
R16192 D.n14086 D.n14085 0.084
R16193 D.n13185 D.n13184 0.084
R16194 D.n12302 D.n12301 0.084
R16195 D.n12238 D.n12237 0.084
R16196 D.n11439 D.n11438 0.084
R16197 D.n10720 D.n10719 0.084
R16198 D.n10127 D.n10126 0.084
R16199 D.n9564 D.n9563 0.084
R16200 D.n9516 D.n9515 0.084
R16201 D.n9037 D.n9036 0.084
R16202 D.n8672 D.n8671 0.084
R16203 D.n8349 D.n8348 0.084
R16204 D.n8313 D.n8312 0.084
R16205 D.n8074 D.n8073 0.084
R16206 D.n7935 D.n7934 0.084
R16207 D.n456 D.n455 0.079
R16208 D.n14072 D.n14071 0.078
R16209 D.n13203 D.n13188 0.078
R16210 D.n13108 D.n13107 0.078
R16211 D.n12320 D.n12305 0.078
R16212 D.n12224 D.n12223 0.078
R16213 D.n11511 D.n11498 0.078
R16214 D.n11425 D.n11424 0.078
R16215 D.n10788 D.n10775 0.078
R16216 D.n10706 D.n10705 0.078
R16217 D.n10145 D.n10130 0.078
R16218 D.n10066 D.n10065 0.078
R16219 D.n9582 D.n9567 0.078
R16220 D.n9502 D.n9501 0.078
R16221 D.n9093 D.n9080 0.078
R16222 D.n9023 D.n9022 0.078
R16223 D.n8690 D.n8675 0.078
R16224 D.n8623 D.n8622 0.078
R16225 D.n8367 D.n8352 0.078
R16226 D.n8299 D.n8298 0.078
R16227 D.n8118 D.n8105 0.078
R16228 D.n8060 D.n8059 0.078
R16229 D.n7953 D.n7938 0.078
R16230 D.n7861 D.n7860 0.077
R16231 D.n7833 D.n7823 0.077
R16232 D.n13124 D.n13123 0.077
R16233 D.n13119 D.n13118 0.077
R16234 D.n11494 D.n11493 0.077
R16235 D.n10771 D.n10770 0.077
R16236 D.n10082 D.n10081 0.077
R16237 D.n10077 D.n10076 0.077
R16238 D.n9076 D.n9075 0.077
R16239 D.n8639 D.n8638 0.077
R16240 D.n8634 D.n8633 0.077
R16241 D.n8101 D.n8100 0.077
R16242 D.n3 D.n2 0.075
R16243 D.n24 D.n16 0.075
R16244 D.n13613 D.n13603 0.074
R16245 D.n13593 D.n13583 0.074
R16246 D.n13573 D.n13563 0.074
R16247 D.n13553 D.n13543 0.074
R16248 D.n13533 D.n13523 0.074
R16249 D.n13513 D.n13503 0.074
R16250 D.n13493 D.n13483 0.074
R16251 D.n13473 D.n13463 0.074
R16252 D.n13453 D.n13443 0.074
R16253 D.n13433 D.n13423 0.074
R16254 D.n13413 D.n13403 0.074
R16255 D.n13393 D.n13383 0.074
R16256 D.n13373 D.n13363 0.074
R16257 D.n13353 D.n13343 0.074
R16258 D.n13333 D.n13323 0.074
R16259 D.n13313 D.n13303 0.074
R16260 D.n13293 D.n13283 0.074
R16261 D.n13273 D.n13263 0.074
R16262 D.n13253 D.n13243 0.074
R16263 D.n13233 D.n13223 0.074
R16264 D.n12690 D.n12680 0.074
R16265 D.n12670 D.n12660 0.074
R16266 D.n12650 D.n12640 0.074
R16267 D.n12630 D.n12620 0.074
R16268 D.n12610 D.n12600 0.074
R16269 D.n12590 D.n12580 0.074
R16270 D.n12570 D.n12560 0.074
R16271 D.n12550 D.n12540 0.074
R16272 D.n12530 D.n12520 0.074
R16273 D.n12510 D.n12500 0.074
R16274 D.n12490 D.n12480 0.074
R16275 D.n12470 D.n12460 0.074
R16276 D.n12450 D.n12440 0.074
R16277 D.n12430 D.n12420 0.074
R16278 D.n12410 D.n12400 0.074
R16279 D.n12390 D.n12380 0.074
R16280 D.n12370 D.n12360 0.074
R16281 D.n12350 D.n12340 0.074
R16282 D.n11841 D.n11831 0.074
R16283 D.n11821 D.n11811 0.074
R16284 D.n11801 D.n11791 0.074
R16285 D.n11781 D.n11771 0.074
R16286 D.n11761 D.n11751 0.074
R16287 D.n11741 D.n11731 0.074
R16288 D.n11721 D.n11711 0.074
R16289 D.n11701 D.n11691 0.074
R16290 D.n11681 D.n11671 0.074
R16291 D.n11661 D.n11651 0.074
R16292 D.n11641 D.n11631 0.074
R16293 D.n11621 D.n11611 0.074
R16294 D.n11601 D.n11591 0.074
R16295 D.n11581 D.n11571 0.074
R16296 D.n11561 D.n11551 0.074
R16297 D.n11541 D.n11531 0.074
R16298 D.n11078 D.n11068 0.074
R16299 D.n11058 D.n11048 0.074
R16300 D.n11038 D.n11028 0.074
R16301 D.n11018 D.n11008 0.074
R16302 D.n10998 D.n10988 0.074
R16303 D.n10978 D.n10968 0.074
R16304 D.n10958 D.n10948 0.074
R16305 D.n10938 D.n10928 0.074
R16306 D.n10918 D.n10908 0.074
R16307 D.n10898 D.n10888 0.074
R16308 D.n10878 D.n10868 0.074
R16309 D.n10858 D.n10848 0.074
R16310 D.n10838 D.n10828 0.074
R16311 D.n10818 D.n10808 0.074
R16312 D.n10395 D.n10385 0.074
R16313 D.n10375 D.n10365 0.074
R16314 D.n10355 D.n10345 0.074
R16315 D.n10335 D.n10325 0.074
R16316 D.n10315 D.n10305 0.074
R16317 D.n10295 D.n10285 0.074
R16318 D.n10275 D.n10265 0.074
R16319 D.n10255 D.n10245 0.074
R16320 D.n10235 D.n10225 0.074
R16321 D.n10215 D.n10205 0.074
R16322 D.n10195 D.n10185 0.074
R16323 D.n10175 D.n10165 0.074
R16324 D.n9792 D.n9782 0.074
R16325 D.n9772 D.n9762 0.074
R16326 D.n9752 D.n9742 0.074
R16327 D.n9732 D.n9722 0.074
R16328 D.n9712 D.n9702 0.074
R16329 D.n9692 D.n9682 0.074
R16330 D.n9672 D.n9662 0.074
R16331 D.n9652 D.n9642 0.074
R16332 D.n9632 D.n9622 0.074
R16333 D.n9612 D.n9602 0.074
R16334 D.n9263 D.n9253 0.074
R16335 D.n9243 D.n9233 0.074
R16336 D.n9223 D.n9213 0.074
R16337 D.n9203 D.n9193 0.074
R16338 D.n9183 D.n9173 0.074
R16339 D.n9163 D.n9153 0.074
R16340 D.n9143 D.n9133 0.074
R16341 D.n9123 D.n9113 0.074
R16342 D.n8820 D.n8810 0.074
R16343 D.n8800 D.n8790 0.074
R16344 D.n8780 D.n8770 0.074
R16345 D.n8760 D.n8750 0.074
R16346 D.n8740 D.n8730 0.074
R16347 D.n8720 D.n8710 0.074
R16348 D.n8457 D.n8447 0.074
R16349 D.n8437 D.n8427 0.074
R16350 D.n8417 D.n8407 0.074
R16351 D.n8397 D.n8387 0.074
R16352 D.n8168 D.n8158 0.074
R16353 D.n8148 D.n8138 0.074
R16354 D.n7983 D.n7982 0.073
R16355 D.n13654 D.n13653 0.073
R16356 D.n13653 D.n13652 0.073
R16357 D.n13674 D.n13673 0.073
R16358 D.n13673 D.n13672 0.073
R16359 D.n13619 D.n13618 0.073
R16360 D.n13631 D.n13630 0.073
R16361 D.n12731 D.n12730 0.073
R16362 D.n12730 D.n12729 0.073
R16363 D.n12747 D.n12746 0.073
R16364 D.n12746 D.n12745 0.073
R16365 D.n12696 D.n12695 0.073
R16366 D.n12708 D.n12707 0.073
R16367 D.n11882 D.n11881 0.073
R16368 D.n11881 D.n11880 0.073
R16369 D.n11898 D.n11897 0.073
R16370 D.n11897 D.n11896 0.073
R16371 D.n11847 D.n11846 0.073
R16372 D.n11859 D.n11858 0.073
R16373 D.n11119 D.n11118 0.073
R16374 D.n11118 D.n11117 0.073
R16375 D.n11135 D.n11134 0.073
R16376 D.n11134 D.n11133 0.073
R16377 D.n11084 D.n11083 0.073
R16378 D.n11096 D.n11095 0.073
R16379 D.n10436 D.n10435 0.073
R16380 D.n10435 D.n10434 0.073
R16381 D.n10452 D.n10451 0.073
R16382 D.n10451 D.n10450 0.073
R16383 D.n10401 D.n10400 0.073
R16384 D.n10413 D.n10412 0.073
R16385 D.n9833 D.n9832 0.073
R16386 D.n9832 D.n9831 0.073
R16387 D.n9849 D.n9848 0.073
R16388 D.n9848 D.n9847 0.073
R16389 D.n9798 D.n9797 0.073
R16390 D.n9810 D.n9809 0.073
R16391 D.n9304 D.n9303 0.073
R16392 D.n9303 D.n9302 0.073
R16393 D.n9320 D.n9319 0.073
R16394 D.n9319 D.n9318 0.073
R16395 D.n9269 D.n9268 0.073
R16396 D.n9281 D.n9280 0.073
R16397 D.n8861 D.n8860 0.073
R16398 D.n8860 D.n8859 0.073
R16399 D.n8877 D.n8876 0.073
R16400 D.n8876 D.n8875 0.073
R16401 D.n8826 D.n8825 0.073
R16402 D.n8838 D.n8837 0.073
R16403 D.n8498 D.n8497 0.073
R16404 D.n8497 D.n8496 0.073
R16405 D.n8514 D.n8513 0.073
R16406 D.n8513 D.n8512 0.073
R16407 D.n8463 D.n8462 0.073
R16408 D.n8475 D.n8474 0.073
R16409 D.n8209 D.n8208 0.073
R16410 D.n8208 D.n8207 0.073
R16411 D.n8225 D.n8224 0.073
R16412 D.n8224 D.n8223 0.073
R16413 D.n8174 D.n8173 0.073
R16414 D.n8186 D.n8185 0.073
R16415 D.n8006 D.n8005 0.073
R16416 D.n8005 D.n8004 0.073
R16417 D.n8022 D.n8021 0.073
R16418 D.n8021 D.n8020 0.073
R16419 D.n7969 D.n7968 0.073
R16420 D.n13213 D.n13203 0.073
R16421 D.n12330 D.n12320 0.073
R16422 D.n11521 D.n11511 0.073
R16423 D.n10798 D.n10788 0.073
R16424 D.n10155 D.n10145 0.073
R16425 D.n9592 D.n9582 0.073
R16426 D.n9103 D.n9093 0.073
R16427 D.n8700 D.n8690 0.073
R16428 D.n8377 D.n8367 0.073
R16429 D.n8128 D.n8118 0.073
R16430 D.n13128 D.n13127 0.072
R16431 D.n10086 D.n10085 0.072
R16432 D.n8643 D.n8642 0.072
R16433 D.n42 D.n34 0.072
R16434 D.n7963 D.n7953 0.072
R16435 D.n7843 D.n7833 0.072
R16436 D.n13223 D.n13213 0.072
R16437 D.n13243 D.n13233 0.072
R16438 D.n13263 D.n13253 0.072
R16439 D.n13283 D.n13273 0.072
R16440 D.n13303 D.n13293 0.072
R16441 D.n13323 D.n13313 0.072
R16442 D.n13343 D.n13333 0.072
R16443 D.n13363 D.n13353 0.072
R16444 D.n13383 D.n13373 0.072
R16445 D.n13403 D.n13393 0.072
R16446 D.n13423 D.n13413 0.072
R16447 D.n13443 D.n13433 0.072
R16448 D.n13463 D.n13453 0.072
R16449 D.n13483 D.n13473 0.072
R16450 D.n13503 D.n13493 0.072
R16451 D.n13523 D.n13513 0.072
R16452 D.n13543 D.n13533 0.072
R16453 D.n13563 D.n13553 0.072
R16454 D.n13583 D.n13573 0.072
R16455 D.n13603 D.n13593 0.072
R16456 D.n12340 D.n12330 0.072
R16457 D.n12360 D.n12350 0.072
R16458 D.n12380 D.n12370 0.072
R16459 D.n12400 D.n12390 0.072
R16460 D.n12420 D.n12410 0.072
R16461 D.n12440 D.n12430 0.072
R16462 D.n12460 D.n12450 0.072
R16463 D.n12480 D.n12470 0.072
R16464 D.n12500 D.n12490 0.072
R16465 D.n12520 D.n12510 0.072
R16466 D.n12540 D.n12530 0.072
R16467 D.n12560 D.n12550 0.072
R16468 D.n12580 D.n12570 0.072
R16469 D.n12600 D.n12590 0.072
R16470 D.n12620 D.n12610 0.072
R16471 D.n12640 D.n12630 0.072
R16472 D.n12660 D.n12650 0.072
R16473 D.n12680 D.n12670 0.072
R16474 D.n11531 D.n11521 0.072
R16475 D.n11551 D.n11541 0.072
R16476 D.n11571 D.n11561 0.072
R16477 D.n11591 D.n11581 0.072
R16478 D.n11611 D.n11601 0.072
R16479 D.n11631 D.n11621 0.072
R16480 D.n11651 D.n11641 0.072
R16481 D.n11671 D.n11661 0.072
R16482 D.n11691 D.n11681 0.072
R16483 D.n11711 D.n11701 0.072
R16484 D.n11731 D.n11721 0.072
R16485 D.n11751 D.n11741 0.072
R16486 D.n11771 D.n11761 0.072
R16487 D.n11791 D.n11781 0.072
R16488 D.n11811 D.n11801 0.072
R16489 D.n11831 D.n11821 0.072
R16490 D.n10808 D.n10798 0.072
R16491 D.n10828 D.n10818 0.072
R16492 D.n10848 D.n10838 0.072
R16493 D.n10868 D.n10858 0.072
R16494 D.n10888 D.n10878 0.072
R16495 D.n10908 D.n10898 0.072
R16496 D.n10928 D.n10918 0.072
R16497 D.n10948 D.n10938 0.072
R16498 D.n10968 D.n10958 0.072
R16499 D.n10988 D.n10978 0.072
R16500 D.n11008 D.n10998 0.072
R16501 D.n11028 D.n11018 0.072
R16502 D.n11048 D.n11038 0.072
R16503 D.n11068 D.n11058 0.072
R16504 D.n10165 D.n10155 0.072
R16505 D.n10185 D.n10175 0.072
R16506 D.n10205 D.n10195 0.072
R16507 D.n10225 D.n10215 0.072
R16508 D.n10245 D.n10235 0.072
R16509 D.n10265 D.n10255 0.072
R16510 D.n10285 D.n10275 0.072
R16511 D.n10305 D.n10295 0.072
R16512 D.n10325 D.n10315 0.072
R16513 D.n10345 D.n10335 0.072
R16514 D.n10365 D.n10355 0.072
R16515 D.n10385 D.n10375 0.072
R16516 D.n9602 D.n9592 0.072
R16517 D.n9622 D.n9612 0.072
R16518 D.n9642 D.n9632 0.072
R16519 D.n9662 D.n9652 0.072
R16520 D.n9682 D.n9672 0.072
R16521 D.n9702 D.n9692 0.072
R16522 D.n9722 D.n9712 0.072
R16523 D.n9742 D.n9732 0.072
R16524 D.n9762 D.n9752 0.072
R16525 D.n9782 D.n9772 0.072
R16526 D.n9113 D.n9103 0.072
R16527 D.n9133 D.n9123 0.072
R16528 D.n9153 D.n9143 0.072
R16529 D.n9173 D.n9163 0.072
R16530 D.n9193 D.n9183 0.072
R16531 D.n9213 D.n9203 0.072
R16532 D.n9233 D.n9223 0.072
R16533 D.n9253 D.n9243 0.072
R16534 D.n8710 D.n8700 0.072
R16535 D.n8730 D.n8720 0.072
R16536 D.n8750 D.n8740 0.072
R16537 D.n8770 D.n8760 0.072
R16538 D.n8790 D.n8780 0.072
R16539 D.n8810 D.n8800 0.072
R16540 D.n8387 D.n8377 0.072
R16541 D.n8407 D.n8397 0.072
R16542 D.n8427 D.n8417 0.072
R16543 D.n8447 D.n8437 0.072
R16544 D.n8138 D.n8128 0.072
R16545 D.n8158 D.n8148 0.072
R16546 D.n14097 D.n14096 0.071
R16547 D.n46 D.n45 0.068
R16548 D.n10 D.n3 0.064
R16549 D.n508 D.n12 0.06
R16550 D.n12249 D.n12248 0.059
R16551 D.n11450 D.n11449 0.059
R16552 D.n10731 D.n10730 0.059
R16553 D.n9527 D.n9526 0.059
R16554 D.n9048 D.n9047 0.059
R16555 D.n8324 D.n8323 0.059
R16556 D.n8085 D.n8084 0.059
R16557 D.n14144 D.n14143 0.057
R16558 D.n534 D.n533 0.056
R16559 D.n1161 D.n1160 0.056
R16560 D.n1760 D.n1759 0.056
R16561 D.n2331 D.n2330 0.056
R16562 D.n2874 D.n2873 0.056
R16563 D.n3390 D.n3389 0.056
R16564 D.n3878 D.n3877 0.056
R16565 D.n4338 D.n4337 0.056
R16566 D.n4770 D.n4769 0.056
R16567 D.n5174 D.n5173 0.056
R16568 D.n5550 D.n5549 0.056
R16569 D.n5898 D.n5897 0.056
R16570 D.n6218 D.n6217 0.056
R16571 D.n6510 D.n6509 0.056
R16572 D.n6774 D.n6773 0.056
R16573 D.n7010 D.n7009 0.056
R16574 D.n7218 D.n7217 0.056
R16575 D.n7398 D.n7397 0.056
R16576 D.n7550 D.n7549 0.056
R16577 D.n7674 D.n7673 0.056
R16578 D.n7769 D.n7768 0.056
R16579 D.n12 D.n10 0.055
R16580 D.n517 D.n516 0.055
R16581 D.n7808 D.n7807 0.055
R16582 D.n7900 D.n7899 0.053
R16583 D.n7810 D.n7809 0.053
R16584 D.n49 D.n48 0.053
R16585 D.n7964 D.n7963 0.053
R16586 D.n13688 D.n13687 0.053
R16587 D.n13614 D.n13613 0.053
R16588 D.n12761 D.n12760 0.053
R16589 D.n12691 D.n12690 0.053
R16590 D.n11912 D.n11911 0.053
R16591 D.n11842 D.n11841 0.053
R16592 D.n11149 D.n11148 0.053
R16593 D.n11079 D.n11078 0.053
R16594 D.n10466 D.n10465 0.053
R16595 D.n10396 D.n10395 0.053
R16596 D.n9863 D.n9862 0.053
R16597 D.n9793 D.n9792 0.053
R16598 D.n9334 D.n9333 0.053
R16599 D.n9264 D.n9263 0.053
R16600 D.n8891 D.n8890 0.053
R16601 D.n8821 D.n8820 0.053
R16602 D.n8528 D.n8527 0.053
R16603 D.n8458 D.n8457 0.053
R16604 D.n8239 D.n8238 0.053
R16605 D.n8169 D.n8168 0.053
R16606 D.n8036 D.n8035 0.053
R16607 D.n7840 D.n7839 0.052
R16608 D.n7830 D.n7829 0.052
R16609 D.n451 D.n450 0.052
R16610 D.n442 D.n441 0.052
R16611 D.n33 D.n32 0.052
R16612 D.n7960 D.n7959 0.052
R16613 D.n7945 D.n7944 0.052
R16614 D.n14065 D.n14064 0.052
R16615 D.n14047 D.n14046 0.052
R16616 D.n14029 D.n14028 0.052
R16617 D.n14011 D.n14010 0.052
R16618 D.n13993 D.n13992 0.052
R16619 D.n13975 D.n13974 0.052
R16620 D.n13957 D.n13956 0.052
R16621 D.n13939 D.n13938 0.052
R16622 D.n13921 D.n13920 0.052
R16623 D.n13903 D.n13902 0.052
R16624 D.n13885 D.n13884 0.052
R16625 D.n13867 D.n13866 0.052
R16626 D.n13849 D.n13848 0.052
R16627 D.n13831 D.n13830 0.052
R16628 D.n13813 D.n13812 0.052
R16629 D.n13795 D.n13794 0.052
R16630 D.n13777 D.n13776 0.052
R16631 D.n13759 D.n13758 0.052
R16632 D.n13741 D.n13740 0.052
R16633 D.n13723 D.n13722 0.052
R16634 D.n13705 D.n13704 0.052
R16635 D.n13686 D.n13685 0.052
R16636 D.n13696 D.n13695 0.052
R16637 D.n13714 D.n13713 0.052
R16638 D.n13732 D.n13731 0.052
R16639 D.n13750 D.n13749 0.052
R16640 D.n13768 D.n13767 0.052
R16641 D.n13786 D.n13785 0.052
R16642 D.n13804 D.n13803 0.052
R16643 D.n13822 D.n13821 0.052
R16644 D.n13840 D.n13839 0.052
R16645 D.n13858 D.n13857 0.052
R16646 D.n13876 D.n13875 0.052
R16647 D.n13894 D.n13893 0.052
R16648 D.n13912 D.n13911 0.052
R16649 D.n13930 D.n13929 0.052
R16650 D.n13948 D.n13947 0.052
R16651 D.n13966 D.n13965 0.052
R16652 D.n13984 D.n13983 0.052
R16653 D.n14002 D.n14001 0.052
R16654 D.n14020 D.n14019 0.052
R16655 D.n14038 D.n14037 0.052
R16656 D.n14056 D.n14055 0.052
R16657 D.n14078 D.n14077 0.052
R16658 D.n13211 D.n13210 0.052
R16659 D.n13231 D.n13230 0.052
R16660 D.n13251 D.n13250 0.052
R16661 D.n13271 D.n13270 0.052
R16662 D.n13291 D.n13290 0.052
R16663 D.n13311 D.n13310 0.052
R16664 D.n13331 D.n13330 0.052
R16665 D.n13351 D.n13350 0.052
R16666 D.n13371 D.n13370 0.052
R16667 D.n13391 D.n13390 0.052
R16668 D.n13411 D.n13410 0.052
R16669 D.n13431 D.n13430 0.052
R16670 D.n13451 D.n13450 0.052
R16671 D.n13471 D.n13470 0.052
R16672 D.n13491 D.n13490 0.052
R16673 D.n13511 D.n13510 0.052
R16674 D.n13531 D.n13530 0.052
R16675 D.n13551 D.n13550 0.052
R16676 D.n13571 D.n13570 0.052
R16677 D.n13591 D.n13590 0.052
R16678 D.n13611 D.n13610 0.052
R16679 D.n13600 D.n13599 0.052
R16680 D.n13580 D.n13579 0.052
R16681 D.n13560 D.n13559 0.052
R16682 D.n13540 D.n13539 0.052
R16683 D.n13520 D.n13519 0.052
R16684 D.n13500 D.n13499 0.052
R16685 D.n13480 D.n13479 0.052
R16686 D.n13460 D.n13459 0.052
R16687 D.n13440 D.n13439 0.052
R16688 D.n13420 D.n13419 0.052
R16689 D.n13400 D.n13399 0.052
R16690 D.n13380 D.n13379 0.052
R16691 D.n13360 D.n13359 0.052
R16692 D.n13340 D.n13339 0.052
R16693 D.n13320 D.n13319 0.052
R16694 D.n13300 D.n13299 0.052
R16695 D.n13280 D.n13279 0.052
R16696 D.n13260 D.n13259 0.052
R16697 D.n13240 D.n13239 0.052
R16698 D.n13220 D.n13219 0.052
R16699 D.n13195 D.n13194 0.052
R16700 D.n13102 D.n13101 0.052
R16701 D.n13084 D.n13083 0.052
R16702 D.n13066 D.n13065 0.052
R16703 D.n13048 D.n13047 0.052
R16704 D.n13030 D.n13029 0.052
R16705 D.n13012 D.n13011 0.052
R16706 D.n12994 D.n12993 0.052
R16707 D.n12976 D.n12975 0.052
R16708 D.n12958 D.n12957 0.052
R16709 D.n12940 D.n12939 0.052
R16710 D.n12922 D.n12921 0.052
R16711 D.n12904 D.n12903 0.052
R16712 D.n12886 D.n12885 0.052
R16713 D.n12868 D.n12867 0.052
R16714 D.n12850 D.n12849 0.052
R16715 D.n12832 D.n12831 0.052
R16716 D.n12814 D.n12813 0.052
R16717 D.n12796 D.n12795 0.052
R16718 D.n12778 D.n12777 0.052
R16719 D.n12759 D.n12758 0.052
R16720 D.n12769 D.n12768 0.052
R16721 D.n12787 D.n12786 0.052
R16722 D.n12805 D.n12804 0.052
R16723 D.n12823 D.n12822 0.052
R16724 D.n12841 D.n12840 0.052
R16725 D.n12859 D.n12858 0.052
R16726 D.n12877 D.n12876 0.052
R16727 D.n12895 D.n12894 0.052
R16728 D.n12913 D.n12912 0.052
R16729 D.n12931 D.n12930 0.052
R16730 D.n12949 D.n12948 0.052
R16731 D.n12967 D.n12966 0.052
R16732 D.n12985 D.n12984 0.052
R16733 D.n13003 D.n13002 0.052
R16734 D.n13021 D.n13020 0.052
R16735 D.n13039 D.n13038 0.052
R16736 D.n13057 D.n13056 0.052
R16737 D.n13075 D.n13074 0.052
R16738 D.n13093 D.n13092 0.052
R16739 D.n13114 D.n13113 0.052
R16740 D.n12328 D.n12327 0.052
R16741 D.n12348 D.n12347 0.052
R16742 D.n12368 D.n12367 0.052
R16743 D.n12388 D.n12387 0.052
R16744 D.n12408 D.n12407 0.052
R16745 D.n12428 D.n12427 0.052
R16746 D.n12448 D.n12447 0.052
R16747 D.n12468 D.n12467 0.052
R16748 D.n12488 D.n12487 0.052
R16749 D.n12508 D.n12507 0.052
R16750 D.n12528 D.n12527 0.052
R16751 D.n12548 D.n12547 0.052
R16752 D.n12568 D.n12567 0.052
R16753 D.n12588 D.n12587 0.052
R16754 D.n12608 D.n12607 0.052
R16755 D.n12628 D.n12627 0.052
R16756 D.n12648 D.n12647 0.052
R16757 D.n12668 D.n12667 0.052
R16758 D.n12688 D.n12687 0.052
R16759 D.n12677 D.n12676 0.052
R16760 D.n12657 D.n12656 0.052
R16761 D.n12637 D.n12636 0.052
R16762 D.n12617 D.n12616 0.052
R16763 D.n12597 D.n12596 0.052
R16764 D.n12577 D.n12576 0.052
R16765 D.n12557 D.n12556 0.052
R16766 D.n12537 D.n12536 0.052
R16767 D.n12517 D.n12516 0.052
R16768 D.n12497 D.n12496 0.052
R16769 D.n12477 D.n12476 0.052
R16770 D.n12457 D.n12456 0.052
R16771 D.n12437 D.n12436 0.052
R16772 D.n12417 D.n12416 0.052
R16773 D.n12397 D.n12396 0.052
R16774 D.n12377 D.n12376 0.052
R16775 D.n12357 D.n12356 0.052
R16776 D.n12337 D.n12336 0.052
R16777 D.n12312 D.n12311 0.052
R16778 D.n12217 D.n12216 0.052
R16779 D.n12199 D.n12198 0.052
R16780 D.n12181 D.n12180 0.052
R16781 D.n12163 D.n12162 0.052
R16782 D.n12145 D.n12144 0.052
R16783 D.n12127 D.n12126 0.052
R16784 D.n12109 D.n12108 0.052
R16785 D.n12091 D.n12090 0.052
R16786 D.n12073 D.n12072 0.052
R16787 D.n12055 D.n12054 0.052
R16788 D.n12037 D.n12036 0.052
R16789 D.n12019 D.n12018 0.052
R16790 D.n12001 D.n12000 0.052
R16791 D.n11983 D.n11982 0.052
R16792 D.n11965 D.n11964 0.052
R16793 D.n11947 D.n11946 0.052
R16794 D.n11929 D.n11928 0.052
R16795 D.n11910 D.n11909 0.052
R16796 D.n11920 D.n11919 0.052
R16797 D.n11938 D.n11937 0.052
R16798 D.n11956 D.n11955 0.052
R16799 D.n11974 D.n11973 0.052
R16800 D.n11992 D.n11991 0.052
R16801 D.n12010 D.n12009 0.052
R16802 D.n12028 D.n12027 0.052
R16803 D.n12046 D.n12045 0.052
R16804 D.n12064 D.n12063 0.052
R16805 D.n12082 D.n12081 0.052
R16806 D.n12100 D.n12099 0.052
R16807 D.n12118 D.n12117 0.052
R16808 D.n12136 D.n12135 0.052
R16809 D.n12154 D.n12153 0.052
R16810 D.n12172 D.n12171 0.052
R16811 D.n12190 D.n12189 0.052
R16812 D.n12208 D.n12207 0.052
R16813 D.n12230 D.n12229 0.052
R16814 D.n11519 D.n11518 0.052
R16815 D.n11539 D.n11538 0.052
R16816 D.n11559 D.n11558 0.052
R16817 D.n11579 D.n11578 0.052
R16818 D.n11599 D.n11598 0.052
R16819 D.n11619 D.n11618 0.052
R16820 D.n11639 D.n11638 0.052
R16821 D.n11659 D.n11658 0.052
R16822 D.n11679 D.n11678 0.052
R16823 D.n11699 D.n11698 0.052
R16824 D.n11719 D.n11718 0.052
R16825 D.n11739 D.n11738 0.052
R16826 D.n11759 D.n11758 0.052
R16827 D.n11779 D.n11778 0.052
R16828 D.n11799 D.n11798 0.052
R16829 D.n11819 D.n11818 0.052
R16830 D.n11839 D.n11838 0.052
R16831 D.n11828 D.n11827 0.052
R16832 D.n11808 D.n11807 0.052
R16833 D.n11788 D.n11787 0.052
R16834 D.n11768 D.n11767 0.052
R16835 D.n11748 D.n11747 0.052
R16836 D.n11728 D.n11727 0.052
R16837 D.n11708 D.n11707 0.052
R16838 D.n11688 D.n11687 0.052
R16839 D.n11668 D.n11667 0.052
R16840 D.n11648 D.n11647 0.052
R16841 D.n11628 D.n11627 0.052
R16842 D.n11608 D.n11607 0.052
R16843 D.n11588 D.n11587 0.052
R16844 D.n11568 D.n11567 0.052
R16845 D.n11548 D.n11547 0.052
R16846 D.n11528 D.n11527 0.052
R16847 D.n11505 D.n11504 0.052
R16848 D.n11418 D.n11417 0.052
R16849 D.n11400 D.n11399 0.052
R16850 D.n11382 D.n11381 0.052
R16851 D.n11364 D.n11363 0.052
R16852 D.n11346 D.n11345 0.052
R16853 D.n11328 D.n11327 0.052
R16854 D.n11310 D.n11309 0.052
R16855 D.n11292 D.n11291 0.052
R16856 D.n11274 D.n11273 0.052
R16857 D.n11256 D.n11255 0.052
R16858 D.n11238 D.n11237 0.052
R16859 D.n11220 D.n11219 0.052
R16860 D.n11202 D.n11201 0.052
R16861 D.n11184 D.n11183 0.052
R16862 D.n11166 D.n11165 0.052
R16863 D.n11147 D.n11146 0.052
R16864 D.n11157 D.n11156 0.052
R16865 D.n11175 D.n11174 0.052
R16866 D.n11193 D.n11192 0.052
R16867 D.n11211 D.n11210 0.052
R16868 D.n11229 D.n11228 0.052
R16869 D.n11247 D.n11246 0.052
R16870 D.n11265 D.n11264 0.052
R16871 D.n11283 D.n11282 0.052
R16872 D.n11301 D.n11300 0.052
R16873 D.n11319 D.n11318 0.052
R16874 D.n11337 D.n11336 0.052
R16875 D.n11355 D.n11354 0.052
R16876 D.n11373 D.n11372 0.052
R16877 D.n11391 D.n11390 0.052
R16878 D.n11409 D.n11408 0.052
R16879 D.n11431 D.n11430 0.052
R16880 D.n10796 D.n10795 0.052
R16881 D.n10816 D.n10815 0.052
R16882 D.n10836 D.n10835 0.052
R16883 D.n10856 D.n10855 0.052
R16884 D.n10876 D.n10875 0.052
R16885 D.n10896 D.n10895 0.052
R16886 D.n10916 D.n10915 0.052
R16887 D.n10936 D.n10935 0.052
R16888 D.n10956 D.n10955 0.052
R16889 D.n10976 D.n10975 0.052
R16890 D.n10996 D.n10995 0.052
R16891 D.n11016 D.n11015 0.052
R16892 D.n11036 D.n11035 0.052
R16893 D.n11056 D.n11055 0.052
R16894 D.n11076 D.n11075 0.052
R16895 D.n11065 D.n11064 0.052
R16896 D.n11045 D.n11044 0.052
R16897 D.n11025 D.n11024 0.052
R16898 D.n11005 D.n11004 0.052
R16899 D.n10985 D.n10984 0.052
R16900 D.n10965 D.n10964 0.052
R16901 D.n10945 D.n10944 0.052
R16902 D.n10925 D.n10924 0.052
R16903 D.n10905 D.n10904 0.052
R16904 D.n10885 D.n10884 0.052
R16905 D.n10865 D.n10864 0.052
R16906 D.n10845 D.n10844 0.052
R16907 D.n10825 D.n10824 0.052
R16908 D.n10805 D.n10804 0.052
R16909 D.n10782 D.n10781 0.052
R16910 D.n10699 D.n10698 0.052
R16911 D.n10681 D.n10680 0.052
R16912 D.n10663 D.n10662 0.052
R16913 D.n10645 D.n10644 0.052
R16914 D.n10627 D.n10626 0.052
R16915 D.n10609 D.n10608 0.052
R16916 D.n10591 D.n10590 0.052
R16917 D.n10573 D.n10572 0.052
R16918 D.n10555 D.n10554 0.052
R16919 D.n10537 D.n10536 0.052
R16920 D.n10519 D.n10518 0.052
R16921 D.n10501 D.n10500 0.052
R16922 D.n10483 D.n10482 0.052
R16923 D.n10464 D.n10463 0.052
R16924 D.n10474 D.n10473 0.052
R16925 D.n10492 D.n10491 0.052
R16926 D.n10510 D.n10509 0.052
R16927 D.n10528 D.n10527 0.052
R16928 D.n10546 D.n10545 0.052
R16929 D.n10564 D.n10563 0.052
R16930 D.n10582 D.n10581 0.052
R16931 D.n10600 D.n10599 0.052
R16932 D.n10618 D.n10617 0.052
R16933 D.n10636 D.n10635 0.052
R16934 D.n10654 D.n10653 0.052
R16935 D.n10672 D.n10671 0.052
R16936 D.n10690 D.n10689 0.052
R16937 D.n10712 D.n10711 0.052
R16938 D.n10153 D.n10152 0.052
R16939 D.n10173 D.n10172 0.052
R16940 D.n10193 D.n10192 0.052
R16941 D.n10213 D.n10212 0.052
R16942 D.n10233 D.n10232 0.052
R16943 D.n10253 D.n10252 0.052
R16944 D.n10273 D.n10272 0.052
R16945 D.n10293 D.n10292 0.052
R16946 D.n10313 D.n10312 0.052
R16947 D.n10333 D.n10332 0.052
R16948 D.n10353 D.n10352 0.052
R16949 D.n10373 D.n10372 0.052
R16950 D.n10393 D.n10392 0.052
R16951 D.n10382 D.n10381 0.052
R16952 D.n10362 D.n10361 0.052
R16953 D.n10342 D.n10341 0.052
R16954 D.n10322 D.n10321 0.052
R16955 D.n10302 D.n10301 0.052
R16956 D.n10282 D.n10281 0.052
R16957 D.n10262 D.n10261 0.052
R16958 D.n10242 D.n10241 0.052
R16959 D.n10222 D.n10221 0.052
R16960 D.n10202 D.n10201 0.052
R16961 D.n10182 D.n10181 0.052
R16962 D.n10162 D.n10161 0.052
R16963 D.n10137 D.n10136 0.052
R16964 D.n10060 D.n10059 0.052
R16965 D.n10042 D.n10041 0.052
R16966 D.n10024 D.n10023 0.052
R16967 D.n10006 D.n10005 0.052
R16968 D.n9988 D.n9987 0.052
R16969 D.n9970 D.n9969 0.052
R16970 D.n9952 D.n9951 0.052
R16971 D.n9934 D.n9933 0.052
R16972 D.n9916 D.n9915 0.052
R16973 D.n9898 D.n9897 0.052
R16974 D.n9880 D.n9879 0.052
R16975 D.n9861 D.n9860 0.052
R16976 D.n9871 D.n9870 0.052
R16977 D.n9889 D.n9888 0.052
R16978 D.n9907 D.n9906 0.052
R16979 D.n9925 D.n9924 0.052
R16980 D.n9943 D.n9942 0.052
R16981 D.n9961 D.n9960 0.052
R16982 D.n9979 D.n9978 0.052
R16983 D.n9997 D.n9996 0.052
R16984 D.n10015 D.n10014 0.052
R16985 D.n10033 D.n10032 0.052
R16986 D.n10051 D.n10050 0.052
R16987 D.n10072 D.n10071 0.052
R16988 D.n9590 D.n9589 0.052
R16989 D.n9610 D.n9609 0.052
R16990 D.n9630 D.n9629 0.052
R16991 D.n9650 D.n9649 0.052
R16992 D.n9670 D.n9669 0.052
R16993 D.n9690 D.n9689 0.052
R16994 D.n9710 D.n9709 0.052
R16995 D.n9730 D.n9729 0.052
R16996 D.n9750 D.n9749 0.052
R16997 D.n9770 D.n9769 0.052
R16998 D.n9790 D.n9789 0.052
R16999 D.n9779 D.n9778 0.052
R17000 D.n9759 D.n9758 0.052
R17001 D.n9739 D.n9738 0.052
R17002 D.n9719 D.n9718 0.052
R17003 D.n9699 D.n9698 0.052
R17004 D.n9679 D.n9678 0.052
R17005 D.n9659 D.n9658 0.052
R17006 D.n9639 D.n9638 0.052
R17007 D.n9619 D.n9618 0.052
R17008 D.n9599 D.n9598 0.052
R17009 D.n9574 D.n9573 0.052
R17010 D.n9495 D.n9494 0.052
R17011 D.n9477 D.n9476 0.052
R17012 D.n9459 D.n9458 0.052
R17013 D.n9441 D.n9440 0.052
R17014 D.n9423 D.n9422 0.052
R17015 D.n9405 D.n9404 0.052
R17016 D.n9387 D.n9386 0.052
R17017 D.n9369 D.n9368 0.052
R17018 D.n9351 D.n9350 0.052
R17019 D.n9332 D.n9331 0.052
R17020 D.n9342 D.n9341 0.052
R17021 D.n9360 D.n9359 0.052
R17022 D.n9378 D.n9377 0.052
R17023 D.n9396 D.n9395 0.052
R17024 D.n9414 D.n9413 0.052
R17025 D.n9432 D.n9431 0.052
R17026 D.n9450 D.n9449 0.052
R17027 D.n9468 D.n9467 0.052
R17028 D.n9486 D.n9485 0.052
R17029 D.n9508 D.n9507 0.052
R17030 D.n9101 D.n9100 0.052
R17031 D.n9121 D.n9120 0.052
R17032 D.n9141 D.n9140 0.052
R17033 D.n9161 D.n9160 0.052
R17034 D.n9181 D.n9180 0.052
R17035 D.n9201 D.n9200 0.052
R17036 D.n9221 D.n9220 0.052
R17037 D.n9241 D.n9240 0.052
R17038 D.n9261 D.n9260 0.052
R17039 D.n9250 D.n9249 0.052
R17040 D.n9230 D.n9229 0.052
R17041 D.n9210 D.n9209 0.052
R17042 D.n9190 D.n9189 0.052
R17043 D.n9170 D.n9169 0.052
R17044 D.n9150 D.n9149 0.052
R17045 D.n9130 D.n9129 0.052
R17046 D.n9110 D.n9109 0.052
R17047 D.n9087 D.n9086 0.052
R17048 D.n9016 D.n9015 0.052
R17049 D.n8998 D.n8997 0.052
R17050 D.n8980 D.n8979 0.052
R17051 D.n8962 D.n8961 0.052
R17052 D.n8944 D.n8943 0.052
R17053 D.n8926 D.n8925 0.052
R17054 D.n8908 D.n8907 0.052
R17055 D.n8889 D.n8888 0.052
R17056 D.n8899 D.n8898 0.052
R17057 D.n8917 D.n8916 0.052
R17058 D.n8935 D.n8934 0.052
R17059 D.n8953 D.n8952 0.052
R17060 D.n8971 D.n8970 0.052
R17061 D.n8989 D.n8988 0.052
R17062 D.n9007 D.n9006 0.052
R17063 D.n9029 D.n9028 0.052
R17064 D.n8698 D.n8697 0.052
R17065 D.n8718 D.n8717 0.052
R17066 D.n8738 D.n8737 0.052
R17067 D.n8758 D.n8757 0.052
R17068 D.n8778 D.n8777 0.052
R17069 D.n8798 D.n8797 0.052
R17070 D.n8818 D.n8817 0.052
R17071 D.n8807 D.n8806 0.052
R17072 D.n8787 D.n8786 0.052
R17073 D.n8767 D.n8766 0.052
R17074 D.n8747 D.n8746 0.052
R17075 D.n8727 D.n8726 0.052
R17076 D.n8707 D.n8706 0.052
R17077 D.n8682 D.n8681 0.052
R17078 D.n8617 D.n8616 0.052
R17079 D.n8599 D.n8598 0.052
R17080 D.n8581 D.n8580 0.052
R17081 D.n8563 D.n8562 0.052
R17082 D.n8545 D.n8544 0.052
R17083 D.n8526 D.n8525 0.052
R17084 D.n8536 D.n8535 0.052
R17085 D.n8554 D.n8553 0.052
R17086 D.n8572 D.n8571 0.052
R17087 D.n8590 D.n8589 0.052
R17088 D.n8608 D.n8607 0.052
R17089 D.n8629 D.n8628 0.052
R17090 D.n8375 D.n8374 0.052
R17091 D.n8395 D.n8394 0.052
R17092 D.n8415 D.n8414 0.052
R17093 D.n8435 D.n8434 0.052
R17094 D.n8455 D.n8454 0.052
R17095 D.n8444 D.n8443 0.052
R17096 D.n8424 D.n8423 0.052
R17097 D.n8404 D.n8403 0.052
R17098 D.n8384 D.n8383 0.052
R17099 D.n8359 D.n8358 0.052
R17100 D.n8292 D.n8291 0.052
R17101 D.n8274 D.n8273 0.052
R17102 D.n8256 D.n8255 0.052
R17103 D.n8237 D.n8236 0.052
R17104 D.n8247 D.n8246 0.052
R17105 D.n8265 D.n8264 0.052
R17106 D.n8283 D.n8282 0.052
R17107 D.n8305 D.n8304 0.052
R17108 D.n8126 D.n8125 0.052
R17109 D.n8146 D.n8145 0.052
R17110 D.n8166 D.n8165 0.052
R17111 D.n8155 D.n8154 0.052
R17112 D.n8135 D.n8134 0.052
R17113 D.n8112 D.n8111 0.052
R17114 D.n8053 D.n8052 0.052
R17115 D.n8034 D.n8033 0.052
R17116 D.n8044 D.n8043 0.052
R17117 D.n8066 D.n8065 0.052
R17118 D.n55 D.n54 0.052
R17119 D.n64 D.n63 0.052
R17120 D.n73 D.n72 0.052
R17121 D.n82 D.n81 0.052
R17122 D.n91 D.n90 0.052
R17123 D.n100 D.n99 0.052
R17124 D.n109 D.n108 0.052
R17125 D.n118 D.n117 0.052
R17126 D.n127 D.n126 0.052
R17127 D.n136 D.n135 0.052
R17128 D.n145 D.n144 0.052
R17129 D.n154 D.n153 0.052
R17130 D.n163 D.n162 0.052
R17131 D.n172 D.n171 0.052
R17132 D.n181 D.n180 0.052
R17133 D.n190 D.n189 0.052
R17134 D.n199 D.n198 0.052
R17135 D.n208 D.n207 0.052
R17136 D.n217 D.n216 0.052
R17137 D.n226 D.n225 0.052
R17138 D.n235 D.n234 0.052
R17139 D.n244 D.n243 0.052
R17140 D.n253 D.n252 0.052
R17141 D.n262 D.n261 0.052
R17142 D.n271 D.n270 0.052
R17143 D.n280 D.n279 0.052
R17144 D.n289 D.n288 0.052
R17145 D.n298 D.n297 0.052
R17146 D.n307 D.n306 0.052
R17147 D.n316 D.n315 0.052
R17148 D.n325 D.n324 0.052
R17149 D.n334 D.n333 0.052
R17150 D.n343 D.n342 0.052
R17151 D.n352 D.n351 0.052
R17152 D.n361 D.n360 0.052
R17153 D.n370 D.n369 0.052
R17154 D.n379 D.n378 0.052
R17155 D.n388 D.n387 0.052
R17156 D.n397 D.n396 0.052
R17157 D.n406 D.n405 0.052
R17158 D.n415 D.n414 0.052
R17159 D.n424 D.n423 0.052
R17160 D.n433 D.n432 0.052
R17161 D.n527 D.n526 0.052
R17162 D.n543 D.n542 0.052
R17163 D.n1131 D.n1130 0.052
R17164 D.n1117 D.n1116 0.052
R17165 D.n1103 D.n1102 0.052
R17166 D.n1089 D.n1088 0.052
R17167 D.n1075 D.n1074 0.052
R17168 D.n1061 D.n1060 0.052
R17169 D.n1047 D.n1046 0.052
R17170 D.n1033 D.n1032 0.052
R17171 D.n1019 D.n1018 0.052
R17172 D.n1005 D.n1004 0.052
R17173 D.n991 D.n990 0.052
R17174 D.n977 D.n976 0.052
R17175 D.n963 D.n962 0.052
R17176 D.n949 D.n948 0.052
R17177 D.n935 D.n934 0.052
R17178 D.n921 D.n920 0.052
R17179 D.n907 D.n906 0.052
R17180 D.n893 D.n892 0.052
R17181 D.n879 D.n878 0.052
R17182 D.n865 D.n864 0.052
R17183 D.n851 D.n850 0.052
R17184 D.n837 D.n836 0.052
R17185 D.n823 D.n822 0.052
R17186 D.n809 D.n808 0.052
R17187 D.n795 D.n794 0.052
R17188 D.n781 D.n780 0.052
R17189 D.n767 D.n766 0.052
R17190 D.n753 D.n752 0.052
R17191 D.n739 D.n738 0.052
R17192 D.n725 D.n724 0.052
R17193 D.n711 D.n710 0.052
R17194 D.n697 D.n696 0.052
R17195 D.n683 D.n682 0.052
R17196 D.n669 D.n668 0.052
R17197 D.n655 D.n654 0.052
R17198 D.n641 D.n640 0.052
R17199 D.n627 D.n626 0.052
R17200 D.n613 D.n612 0.052
R17201 D.n599 D.n598 0.052
R17202 D.n585 D.n584 0.052
R17203 D.n571 D.n570 0.052
R17204 D.n557 D.n556 0.052
R17205 D.n1154 D.n1153 0.052
R17206 D.n1170 D.n1169 0.052
R17207 D.n1730 D.n1729 0.052
R17208 D.n1716 D.n1715 0.052
R17209 D.n1702 D.n1701 0.052
R17210 D.n1688 D.n1687 0.052
R17211 D.n1674 D.n1673 0.052
R17212 D.n1660 D.n1659 0.052
R17213 D.n1646 D.n1645 0.052
R17214 D.n1632 D.n1631 0.052
R17215 D.n1618 D.n1617 0.052
R17216 D.n1604 D.n1603 0.052
R17217 D.n1590 D.n1589 0.052
R17218 D.n1576 D.n1575 0.052
R17219 D.n1562 D.n1561 0.052
R17220 D.n1548 D.n1547 0.052
R17221 D.n1534 D.n1533 0.052
R17222 D.n1520 D.n1519 0.052
R17223 D.n1506 D.n1505 0.052
R17224 D.n1492 D.n1491 0.052
R17225 D.n1478 D.n1477 0.052
R17226 D.n1464 D.n1463 0.052
R17227 D.n1450 D.n1449 0.052
R17228 D.n1436 D.n1435 0.052
R17229 D.n1422 D.n1421 0.052
R17230 D.n1408 D.n1407 0.052
R17231 D.n1394 D.n1393 0.052
R17232 D.n1380 D.n1379 0.052
R17233 D.n1366 D.n1365 0.052
R17234 D.n1352 D.n1351 0.052
R17235 D.n1338 D.n1337 0.052
R17236 D.n1324 D.n1323 0.052
R17237 D.n1310 D.n1309 0.052
R17238 D.n1296 D.n1295 0.052
R17239 D.n1282 D.n1281 0.052
R17240 D.n1268 D.n1267 0.052
R17241 D.n1254 D.n1253 0.052
R17242 D.n1240 D.n1239 0.052
R17243 D.n1226 D.n1225 0.052
R17244 D.n1212 D.n1211 0.052
R17245 D.n1198 D.n1197 0.052
R17246 D.n1184 D.n1183 0.052
R17247 D.n1753 D.n1752 0.052
R17248 D.n1769 D.n1768 0.052
R17249 D.n2301 D.n2300 0.052
R17250 D.n2287 D.n2286 0.052
R17251 D.n2273 D.n2272 0.052
R17252 D.n2259 D.n2258 0.052
R17253 D.n2245 D.n2244 0.052
R17254 D.n2231 D.n2230 0.052
R17255 D.n2217 D.n2216 0.052
R17256 D.n2203 D.n2202 0.052
R17257 D.n2189 D.n2188 0.052
R17258 D.n2175 D.n2174 0.052
R17259 D.n2161 D.n2160 0.052
R17260 D.n2147 D.n2146 0.052
R17261 D.n2133 D.n2132 0.052
R17262 D.n2119 D.n2118 0.052
R17263 D.n2105 D.n2104 0.052
R17264 D.n2091 D.n2090 0.052
R17265 D.n2077 D.n2076 0.052
R17266 D.n2063 D.n2062 0.052
R17267 D.n2049 D.n2048 0.052
R17268 D.n2035 D.n2034 0.052
R17269 D.n2021 D.n2020 0.052
R17270 D.n2007 D.n2006 0.052
R17271 D.n1993 D.n1992 0.052
R17272 D.n1979 D.n1978 0.052
R17273 D.n1965 D.n1964 0.052
R17274 D.n1951 D.n1950 0.052
R17275 D.n1937 D.n1936 0.052
R17276 D.n1923 D.n1922 0.052
R17277 D.n1909 D.n1908 0.052
R17278 D.n1895 D.n1894 0.052
R17279 D.n1881 D.n1880 0.052
R17280 D.n1867 D.n1866 0.052
R17281 D.n1853 D.n1852 0.052
R17282 D.n1839 D.n1838 0.052
R17283 D.n1825 D.n1824 0.052
R17284 D.n1811 D.n1810 0.052
R17285 D.n1797 D.n1796 0.052
R17286 D.n1783 D.n1782 0.052
R17287 D.n2324 D.n2323 0.052
R17288 D.n2340 D.n2339 0.052
R17289 D.n2844 D.n2843 0.052
R17290 D.n2830 D.n2829 0.052
R17291 D.n2816 D.n2815 0.052
R17292 D.n2802 D.n2801 0.052
R17293 D.n2788 D.n2787 0.052
R17294 D.n2774 D.n2773 0.052
R17295 D.n2760 D.n2759 0.052
R17296 D.n2746 D.n2745 0.052
R17297 D.n2732 D.n2731 0.052
R17298 D.n2718 D.n2717 0.052
R17299 D.n2704 D.n2703 0.052
R17300 D.n2690 D.n2689 0.052
R17301 D.n2676 D.n2675 0.052
R17302 D.n2662 D.n2661 0.052
R17303 D.n2648 D.n2647 0.052
R17304 D.n2634 D.n2633 0.052
R17305 D.n2620 D.n2619 0.052
R17306 D.n2606 D.n2605 0.052
R17307 D.n2592 D.n2591 0.052
R17308 D.n2578 D.n2577 0.052
R17309 D.n2564 D.n2563 0.052
R17310 D.n2550 D.n2549 0.052
R17311 D.n2536 D.n2535 0.052
R17312 D.n2522 D.n2521 0.052
R17313 D.n2508 D.n2507 0.052
R17314 D.n2494 D.n2493 0.052
R17315 D.n2480 D.n2479 0.052
R17316 D.n2466 D.n2465 0.052
R17317 D.n2452 D.n2451 0.052
R17318 D.n2438 D.n2437 0.052
R17319 D.n2424 D.n2423 0.052
R17320 D.n2410 D.n2409 0.052
R17321 D.n2396 D.n2395 0.052
R17322 D.n2382 D.n2381 0.052
R17323 D.n2368 D.n2367 0.052
R17324 D.n2354 D.n2353 0.052
R17325 D.n2867 D.n2866 0.052
R17326 D.n2883 D.n2882 0.052
R17327 D.n3359 D.n3358 0.052
R17328 D.n3345 D.n3344 0.052
R17329 D.n3331 D.n3330 0.052
R17330 D.n3317 D.n3316 0.052
R17331 D.n3303 D.n3302 0.052
R17332 D.n3289 D.n3288 0.052
R17333 D.n3275 D.n3274 0.052
R17334 D.n3261 D.n3260 0.052
R17335 D.n3247 D.n3246 0.052
R17336 D.n3233 D.n3232 0.052
R17337 D.n3219 D.n3218 0.052
R17338 D.n3205 D.n3204 0.052
R17339 D.n3191 D.n3190 0.052
R17340 D.n3177 D.n3176 0.052
R17341 D.n3163 D.n3162 0.052
R17342 D.n3149 D.n3148 0.052
R17343 D.n3135 D.n3134 0.052
R17344 D.n3121 D.n3120 0.052
R17345 D.n3107 D.n3106 0.052
R17346 D.n3093 D.n3092 0.052
R17347 D.n3079 D.n3078 0.052
R17348 D.n3065 D.n3064 0.052
R17349 D.n3051 D.n3050 0.052
R17350 D.n3037 D.n3036 0.052
R17351 D.n3023 D.n3022 0.052
R17352 D.n3009 D.n3008 0.052
R17353 D.n2995 D.n2994 0.052
R17354 D.n2981 D.n2980 0.052
R17355 D.n2967 D.n2966 0.052
R17356 D.n2953 D.n2952 0.052
R17357 D.n2939 D.n2938 0.052
R17358 D.n2925 D.n2924 0.052
R17359 D.n2911 D.n2910 0.052
R17360 D.n2897 D.n2896 0.052
R17361 D.n3383 D.n3382 0.052
R17362 D.n3399 D.n3398 0.052
R17363 D.n3847 D.n3846 0.052
R17364 D.n3833 D.n3832 0.052
R17365 D.n3819 D.n3818 0.052
R17366 D.n3805 D.n3804 0.052
R17367 D.n3791 D.n3790 0.052
R17368 D.n3777 D.n3776 0.052
R17369 D.n3763 D.n3762 0.052
R17370 D.n3749 D.n3748 0.052
R17371 D.n3735 D.n3734 0.052
R17372 D.n3721 D.n3720 0.052
R17373 D.n3707 D.n3706 0.052
R17374 D.n3693 D.n3692 0.052
R17375 D.n3679 D.n3678 0.052
R17376 D.n3665 D.n3664 0.052
R17377 D.n3651 D.n3650 0.052
R17378 D.n3637 D.n3636 0.052
R17379 D.n3623 D.n3622 0.052
R17380 D.n3609 D.n3608 0.052
R17381 D.n3595 D.n3594 0.052
R17382 D.n3581 D.n3580 0.052
R17383 D.n3567 D.n3566 0.052
R17384 D.n3553 D.n3552 0.052
R17385 D.n3539 D.n3538 0.052
R17386 D.n3525 D.n3524 0.052
R17387 D.n3511 D.n3510 0.052
R17388 D.n3497 D.n3496 0.052
R17389 D.n3483 D.n3482 0.052
R17390 D.n3469 D.n3468 0.052
R17391 D.n3455 D.n3454 0.052
R17392 D.n3441 D.n3440 0.052
R17393 D.n3427 D.n3426 0.052
R17394 D.n3413 D.n3412 0.052
R17395 D.n3871 D.n3870 0.052
R17396 D.n3887 D.n3886 0.052
R17397 D.n4307 D.n4306 0.052
R17398 D.n4293 D.n4292 0.052
R17399 D.n4279 D.n4278 0.052
R17400 D.n4265 D.n4264 0.052
R17401 D.n4251 D.n4250 0.052
R17402 D.n4237 D.n4236 0.052
R17403 D.n4223 D.n4222 0.052
R17404 D.n4209 D.n4208 0.052
R17405 D.n4195 D.n4194 0.052
R17406 D.n4181 D.n4180 0.052
R17407 D.n4167 D.n4166 0.052
R17408 D.n4153 D.n4152 0.052
R17409 D.n4139 D.n4138 0.052
R17410 D.n4125 D.n4124 0.052
R17411 D.n4111 D.n4110 0.052
R17412 D.n4097 D.n4096 0.052
R17413 D.n4083 D.n4082 0.052
R17414 D.n4069 D.n4068 0.052
R17415 D.n4055 D.n4054 0.052
R17416 D.n4041 D.n4040 0.052
R17417 D.n4027 D.n4026 0.052
R17418 D.n4013 D.n4012 0.052
R17419 D.n3999 D.n3998 0.052
R17420 D.n3985 D.n3984 0.052
R17421 D.n3971 D.n3970 0.052
R17422 D.n3957 D.n3956 0.052
R17423 D.n3943 D.n3942 0.052
R17424 D.n3929 D.n3928 0.052
R17425 D.n3915 D.n3914 0.052
R17426 D.n3901 D.n3900 0.052
R17427 D.n4331 D.n4330 0.052
R17428 D.n4347 D.n4346 0.052
R17429 D.n4739 D.n4738 0.052
R17430 D.n4725 D.n4724 0.052
R17431 D.n4711 D.n4710 0.052
R17432 D.n4697 D.n4696 0.052
R17433 D.n4683 D.n4682 0.052
R17434 D.n4669 D.n4668 0.052
R17435 D.n4655 D.n4654 0.052
R17436 D.n4641 D.n4640 0.052
R17437 D.n4627 D.n4626 0.052
R17438 D.n4613 D.n4612 0.052
R17439 D.n4599 D.n4598 0.052
R17440 D.n4585 D.n4584 0.052
R17441 D.n4571 D.n4570 0.052
R17442 D.n4557 D.n4556 0.052
R17443 D.n4543 D.n4542 0.052
R17444 D.n4529 D.n4528 0.052
R17445 D.n4515 D.n4514 0.052
R17446 D.n4501 D.n4500 0.052
R17447 D.n4487 D.n4486 0.052
R17448 D.n4473 D.n4472 0.052
R17449 D.n4459 D.n4458 0.052
R17450 D.n4445 D.n4444 0.052
R17451 D.n4431 D.n4430 0.052
R17452 D.n4417 D.n4416 0.052
R17453 D.n4403 D.n4402 0.052
R17454 D.n4389 D.n4388 0.052
R17455 D.n4375 D.n4374 0.052
R17456 D.n4361 D.n4360 0.052
R17457 D.n4763 D.n4762 0.052
R17458 D.n4779 D.n4778 0.052
R17459 D.n5143 D.n5142 0.052
R17460 D.n5129 D.n5128 0.052
R17461 D.n5115 D.n5114 0.052
R17462 D.n5101 D.n5100 0.052
R17463 D.n5087 D.n5086 0.052
R17464 D.n5073 D.n5072 0.052
R17465 D.n5059 D.n5058 0.052
R17466 D.n5045 D.n5044 0.052
R17467 D.n5031 D.n5030 0.052
R17468 D.n5017 D.n5016 0.052
R17469 D.n5003 D.n5002 0.052
R17470 D.n4989 D.n4988 0.052
R17471 D.n4975 D.n4974 0.052
R17472 D.n4961 D.n4960 0.052
R17473 D.n4947 D.n4946 0.052
R17474 D.n4933 D.n4932 0.052
R17475 D.n4919 D.n4918 0.052
R17476 D.n4905 D.n4904 0.052
R17477 D.n4891 D.n4890 0.052
R17478 D.n4877 D.n4876 0.052
R17479 D.n4863 D.n4862 0.052
R17480 D.n4849 D.n4848 0.052
R17481 D.n4835 D.n4834 0.052
R17482 D.n4821 D.n4820 0.052
R17483 D.n4807 D.n4806 0.052
R17484 D.n4793 D.n4792 0.052
R17485 D.n5167 D.n5166 0.052
R17486 D.n5183 D.n5182 0.052
R17487 D.n5519 D.n5518 0.052
R17488 D.n5505 D.n5504 0.052
R17489 D.n5491 D.n5490 0.052
R17490 D.n5477 D.n5476 0.052
R17491 D.n5463 D.n5462 0.052
R17492 D.n5449 D.n5448 0.052
R17493 D.n5435 D.n5434 0.052
R17494 D.n5421 D.n5420 0.052
R17495 D.n5407 D.n5406 0.052
R17496 D.n5393 D.n5392 0.052
R17497 D.n5379 D.n5378 0.052
R17498 D.n5365 D.n5364 0.052
R17499 D.n5351 D.n5350 0.052
R17500 D.n5337 D.n5336 0.052
R17501 D.n5323 D.n5322 0.052
R17502 D.n5309 D.n5308 0.052
R17503 D.n5295 D.n5294 0.052
R17504 D.n5281 D.n5280 0.052
R17505 D.n5267 D.n5266 0.052
R17506 D.n5253 D.n5252 0.052
R17507 D.n5239 D.n5238 0.052
R17508 D.n5225 D.n5224 0.052
R17509 D.n5211 D.n5210 0.052
R17510 D.n5197 D.n5196 0.052
R17511 D.n5543 D.n5542 0.052
R17512 D.n5559 D.n5558 0.052
R17513 D.n5867 D.n5866 0.052
R17514 D.n5853 D.n5852 0.052
R17515 D.n5839 D.n5838 0.052
R17516 D.n5825 D.n5824 0.052
R17517 D.n5811 D.n5810 0.052
R17518 D.n5797 D.n5796 0.052
R17519 D.n5783 D.n5782 0.052
R17520 D.n5769 D.n5768 0.052
R17521 D.n5755 D.n5754 0.052
R17522 D.n5741 D.n5740 0.052
R17523 D.n5727 D.n5726 0.052
R17524 D.n5713 D.n5712 0.052
R17525 D.n5699 D.n5698 0.052
R17526 D.n5685 D.n5684 0.052
R17527 D.n5671 D.n5670 0.052
R17528 D.n5657 D.n5656 0.052
R17529 D.n5643 D.n5642 0.052
R17530 D.n5629 D.n5628 0.052
R17531 D.n5615 D.n5614 0.052
R17532 D.n5601 D.n5600 0.052
R17533 D.n5587 D.n5586 0.052
R17534 D.n5573 D.n5572 0.052
R17535 D.n5891 D.n5890 0.052
R17536 D.n5907 D.n5906 0.052
R17537 D.n6187 D.n6186 0.052
R17538 D.n6173 D.n6172 0.052
R17539 D.n6159 D.n6158 0.052
R17540 D.n6145 D.n6144 0.052
R17541 D.n6131 D.n6130 0.052
R17542 D.n6117 D.n6116 0.052
R17543 D.n6103 D.n6102 0.052
R17544 D.n6089 D.n6088 0.052
R17545 D.n6075 D.n6074 0.052
R17546 D.n6061 D.n6060 0.052
R17547 D.n6047 D.n6046 0.052
R17548 D.n6033 D.n6032 0.052
R17549 D.n6019 D.n6018 0.052
R17550 D.n6005 D.n6004 0.052
R17551 D.n5991 D.n5990 0.052
R17552 D.n5977 D.n5976 0.052
R17553 D.n5963 D.n5962 0.052
R17554 D.n5949 D.n5948 0.052
R17555 D.n5935 D.n5934 0.052
R17556 D.n5921 D.n5920 0.052
R17557 D.n6211 D.n6210 0.052
R17558 D.n6227 D.n6226 0.052
R17559 D.n6479 D.n6478 0.052
R17560 D.n6465 D.n6464 0.052
R17561 D.n6451 D.n6450 0.052
R17562 D.n6437 D.n6436 0.052
R17563 D.n6423 D.n6422 0.052
R17564 D.n6409 D.n6408 0.052
R17565 D.n6395 D.n6394 0.052
R17566 D.n6381 D.n6380 0.052
R17567 D.n6367 D.n6366 0.052
R17568 D.n6353 D.n6352 0.052
R17569 D.n6339 D.n6338 0.052
R17570 D.n6325 D.n6324 0.052
R17571 D.n6311 D.n6310 0.052
R17572 D.n6297 D.n6296 0.052
R17573 D.n6283 D.n6282 0.052
R17574 D.n6269 D.n6268 0.052
R17575 D.n6255 D.n6254 0.052
R17576 D.n6241 D.n6240 0.052
R17577 D.n6503 D.n6502 0.052
R17578 D.n6519 D.n6518 0.052
R17579 D.n6743 D.n6742 0.052
R17580 D.n6729 D.n6728 0.052
R17581 D.n6715 D.n6714 0.052
R17582 D.n6701 D.n6700 0.052
R17583 D.n6687 D.n6686 0.052
R17584 D.n6673 D.n6672 0.052
R17585 D.n6659 D.n6658 0.052
R17586 D.n6645 D.n6644 0.052
R17587 D.n6631 D.n6630 0.052
R17588 D.n6617 D.n6616 0.052
R17589 D.n6603 D.n6602 0.052
R17590 D.n6589 D.n6588 0.052
R17591 D.n6575 D.n6574 0.052
R17592 D.n6561 D.n6560 0.052
R17593 D.n6547 D.n6546 0.052
R17594 D.n6533 D.n6532 0.052
R17595 D.n6767 D.n6766 0.052
R17596 D.n6783 D.n6782 0.052
R17597 D.n6979 D.n6978 0.052
R17598 D.n6965 D.n6964 0.052
R17599 D.n6951 D.n6950 0.052
R17600 D.n6937 D.n6936 0.052
R17601 D.n6923 D.n6922 0.052
R17602 D.n6909 D.n6908 0.052
R17603 D.n6895 D.n6894 0.052
R17604 D.n6881 D.n6880 0.052
R17605 D.n6867 D.n6866 0.052
R17606 D.n6853 D.n6852 0.052
R17607 D.n6839 D.n6838 0.052
R17608 D.n6825 D.n6824 0.052
R17609 D.n6811 D.n6810 0.052
R17610 D.n6797 D.n6796 0.052
R17611 D.n7003 D.n7002 0.052
R17612 D.n7019 D.n7018 0.052
R17613 D.n7187 D.n7186 0.052
R17614 D.n7173 D.n7172 0.052
R17615 D.n7159 D.n7158 0.052
R17616 D.n7145 D.n7144 0.052
R17617 D.n7131 D.n7130 0.052
R17618 D.n7117 D.n7116 0.052
R17619 D.n7103 D.n7102 0.052
R17620 D.n7089 D.n7088 0.052
R17621 D.n7075 D.n7074 0.052
R17622 D.n7061 D.n7060 0.052
R17623 D.n7047 D.n7046 0.052
R17624 D.n7033 D.n7032 0.052
R17625 D.n7211 D.n7210 0.052
R17626 D.n7227 D.n7226 0.052
R17627 D.n7367 D.n7366 0.052
R17628 D.n7353 D.n7352 0.052
R17629 D.n7339 D.n7338 0.052
R17630 D.n7325 D.n7324 0.052
R17631 D.n7311 D.n7310 0.052
R17632 D.n7297 D.n7296 0.052
R17633 D.n7283 D.n7282 0.052
R17634 D.n7269 D.n7268 0.052
R17635 D.n7255 D.n7254 0.052
R17636 D.n7241 D.n7240 0.052
R17637 D.n7391 D.n7390 0.052
R17638 D.n7407 D.n7406 0.052
R17639 D.n7519 D.n7518 0.052
R17640 D.n7505 D.n7504 0.052
R17641 D.n7491 D.n7490 0.052
R17642 D.n7477 D.n7476 0.052
R17643 D.n7463 D.n7462 0.052
R17644 D.n7449 D.n7448 0.052
R17645 D.n7435 D.n7434 0.052
R17646 D.n7421 D.n7420 0.052
R17647 D.n7543 D.n7542 0.052
R17648 D.n7559 D.n7558 0.052
R17649 D.n7643 D.n7642 0.052
R17650 D.n7629 D.n7628 0.052
R17651 D.n7615 D.n7614 0.052
R17652 D.n7601 D.n7600 0.052
R17653 D.n7587 D.n7586 0.052
R17654 D.n7573 D.n7572 0.052
R17655 D.n7667 D.n7666 0.052
R17656 D.n7683 D.n7682 0.052
R17657 D.n7739 D.n7738 0.052
R17658 D.n7725 D.n7724 0.052
R17659 D.n7711 D.n7710 0.052
R17660 D.n7697 D.n7696 0.052
R17661 D.n7762 D.n7761 0.052
R17662 D.n7778 D.n7777 0.052
R17663 D.n7806 D.n7805 0.052
R17664 D.n7792 D.n7791 0.052
R17665 D.n7845 D.n7844 0.051
R17666 D.n5 D.n4 0.051
R17667 D.n6 D.n5 0.051
R17668 D.n7 D.n6 0.051
R17669 D.n8 D.n7 0.051
R17670 D.n9 D.n8 0.051
R17671 D.n519 D.n518 0.051
R17672 D.n7837 D.n7836 0.051
R17673 D.n7827 D.n7826 0.051
R17674 D.n448 D.n446 0.051
R17675 D.n439 D.n437 0.051
R17676 D.n30 D.n29 0.051
R17677 D.n7957 D.n7956 0.051
R17678 D.n7942 D.n7941 0.051
R17679 D.n14062 D.n14060 0.051
R17680 D.n14044 D.n14042 0.051
R17681 D.n14026 D.n14024 0.051
R17682 D.n14008 D.n14006 0.051
R17683 D.n13990 D.n13988 0.051
R17684 D.n13972 D.n13970 0.051
R17685 D.n13954 D.n13952 0.051
R17686 D.n13936 D.n13934 0.051
R17687 D.n13918 D.n13916 0.051
R17688 D.n13900 D.n13898 0.051
R17689 D.n13882 D.n13880 0.051
R17690 D.n13864 D.n13862 0.051
R17691 D.n13846 D.n13844 0.051
R17692 D.n13828 D.n13826 0.051
R17693 D.n13810 D.n13808 0.051
R17694 D.n13792 D.n13790 0.051
R17695 D.n13774 D.n13772 0.051
R17696 D.n13756 D.n13754 0.051
R17697 D.n13738 D.n13736 0.051
R17698 D.n13720 D.n13718 0.051
R17699 D.n13702 D.n13700 0.051
R17700 D.n13683 D.n13681 0.051
R17701 D.n13693 D.n13692 0.051
R17702 D.n13711 D.n13710 0.051
R17703 D.n13729 D.n13728 0.051
R17704 D.n13747 D.n13746 0.051
R17705 D.n13765 D.n13764 0.051
R17706 D.n13783 D.n13782 0.051
R17707 D.n13801 D.n13800 0.051
R17708 D.n13819 D.n13818 0.051
R17709 D.n13837 D.n13836 0.051
R17710 D.n13855 D.n13854 0.051
R17711 D.n13873 D.n13872 0.051
R17712 D.n13891 D.n13890 0.051
R17713 D.n13909 D.n13908 0.051
R17714 D.n13927 D.n13926 0.051
R17715 D.n13945 D.n13944 0.051
R17716 D.n13963 D.n13962 0.051
R17717 D.n13981 D.n13980 0.051
R17718 D.n13999 D.n13998 0.051
R17719 D.n14017 D.n14016 0.051
R17720 D.n14035 D.n14034 0.051
R17721 D.n14053 D.n14052 0.051
R17722 D.n14075 D.n14074 0.051
R17723 D.n13208 D.n13206 0.051
R17724 D.n13228 D.n13226 0.051
R17725 D.n13248 D.n13246 0.051
R17726 D.n13268 D.n13266 0.051
R17727 D.n13288 D.n13286 0.051
R17728 D.n13308 D.n13306 0.051
R17729 D.n13328 D.n13326 0.051
R17730 D.n13348 D.n13346 0.051
R17731 D.n13368 D.n13366 0.051
R17732 D.n13388 D.n13386 0.051
R17733 D.n13408 D.n13406 0.051
R17734 D.n13428 D.n13426 0.051
R17735 D.n13448 D.n13446 0.051
R17736 D.n13468 D.n13466 0.051
R17737 D.n13488 D.n13486 0.051
R17738 D.n13508 D.n13506 0.051
R17739 D.n13528 D.n13526 0.051
R17740 D.n13548 D.n13546 0.051
R17741 D.n13568 D.n13566 0.051
R17742 D.n13588 D.n13586 0.051
R17743 D.n13608 D.n13606 0.051
R17744 D.n13597 D.n13596 0.051
R17745 D.n13577 D.n13576 0.051
R17746 D.n13557 D.n13556 0.051
R17747 D.n13537 D.n13536 0.051
R17748 D.n13517 D.n13516 0.051
R17749 D.n13497 D.n13496 0.051
R17750 D.n13477 D.n13476 0.051
R17751 D.n13457 D.n13456 0.051
R17752 D.n13437 D.n13436 0.051
R17753 D.n13417 D.n13416 0.051
R17754 D.n13397 D.n13396 0.051
R17755 D.n13377 D.n13376 0.051
R17756 D.n13357 D.n13356 0.051
R17757 D.n13337 D.n13336 0.051
R17758 D.n13317 D.n13316 0.051
R17759 D.n13297 D.n13296 0.051
R17760 D.n13277 D.n13276 0.051
R17761 D.n13257 D.n13256 0.051
R17762 D.n13237 D.n13236 0.051
R17763 D.n13217 D.n13216 0.051
R17764 D.n13192 D.n13191 0.051
R17765 D.n13099 D.n13097 0.051
R17766 D.n13081 D.n13079 0.051
R17767 D.n13063 D.n13061 0.051
R17768 D.n13045 D.n13043 0.051
R17769 D.n13027 D.n13025 0.051
R17770 D.n13009 D.n13007 0.051
R17771 D.n12991 D.n12989 0.051
R17772 D.n12973 D.n12971 0.051
R17773 D.n12955 D.n12953 0.051
R17774 D.n12937 D.n12935 0.051
R17775 D.n12919 D.n12917 0.051
R17776 D.n12901 D.n12899 0.051
R17777 D.n12883 D.n12881 0.051
R17778 D.n12865 D.n12863 0.051
R17779 D.n12847 D.n12845 0.051
R17780 D.n12829 D.n12827 0.051
R17781 D.n12811 D.n12809 0.051
R17782 D.n12793 D.n12791 0.051
R17783 D.n12775 D.n12773 0.051
R17784 D.n12756 D.n12754 0.051
R17785 D.n12766 D.n12765 0.051
R17786 D.n12784 D.n12783 0.051
R17787 D.n12802 D.n12801 0.051
R17788 D.n12820 D.n12819 0.051
R17789 D.n12838 D.n12837 0.051
R17790 D.n12856 D.n12855 0.051
R17791 D.n12874 D.n12873 0.051
R17792 D.n12892 D.n12891 0.051
R17793 D.n12910 D.n12909 0.051
R17794 D.n12928 D.n12927 0.051
R17795 D.n12946 D.n12945 0.051
R17796 D.n12964 D.n12963 0.051
R17797 D.n12982 D.n12981 0.051
R17798 D.n13000 D.n12999 0.051
R17799 D.n13018 D.n13017 0.051
R17800 D.n13036 D.n13035 0.051
R17801 D.n13054 D.n13053 0.051
R17802 D.n13072 D.n13071 0.051
R17803 D.n13090 D.n13089 0.051
R17804 D.n13111 D.n13110 0.051
R17805 D.n12325 D.n12323 0.051
R17806 D.n12345 D.n12343 0.051
R17807 D.n12365 D.n12363 0.051
R17808 D.n12385 D.n12383 0.051
R17809 D.n12405 D.n12403 0.051
R17810 D.n12425 D.n12423 0.051
R17811 D.n12445 D.n12443 0.051
R17812 D.n12465 D.n12463 0.051
R17813 D.n12485 D.n12483 0.051
R17814 D.n12505 D.n12503 0.051
R17815 D.n12525 D.n12523 0.051
R17816 D.n12545 D.n12543 0.051
R17817 D.n12565 D.n12563 0.051
R17818 D.n12585 D.n12583 0.051
R17819 D.n12605 D.n12603 0.051
R17820 D.n12625 D.n12623 0.051
R17821 D.n12645 D.n12643 0.051
R17822 D.n12665 D.n12663 0.051
R17823 D.n12685 D.n12683 0.051
R17824 D.n12674 D.n12673 0.051
R17825 D.n12654 D.n12653 0.051
R17826 D.n12634 D.n12633 0.051
R17827 D.n12614 D.n12613 0.051
R17828 D.n12594 D.n12593 0.051
R17829 D.n12574 D.n12573 0.051
R17830 D.n12554 D.n12553 0.051
R17831 D.n12534 D.n12533 0.051
R17832 D.n12514 D.n12513 0.051
R17833 D.n12494 D.n12493 0.051
R17834 D.n12474 D.n12473 0.051
R17835 D.n12454 D.n12453 0.051
R17836 D.n12434 D.n12433 0.051
R17837 D.n12414 D.n12413 0.051
R17838 D.n12394 D.n12393 0.051
R17839 D.n12374 D.n12373 0.051
R17840 D.n12354 D.n12353 0.051
R17841 D.n12334 D.n12333 0.051
R17842 D.n12309 D.n12308 0.051
R17843 D.n12214 D.n12212 0.051
R17844 D.n12196 D.n12194 0.051
R17845 D.n12178 D.n12176 0.051
R17846 D.n12160 D.n12158 0.051
R17847 D.n12142 D.n12140 0.051
R17848 D.n12124 D.n12122 0.051
R17849 D.n12106 D.n12104 0.051
R17850 D.n12088 D.n12086 0.051
R17851 D.n12070 D.n12068 0.051
R17852 D.n12052 D.n12050 0.051
R17853 D.n12034 D.n12032 0.051
R17854 D.n12016 D.n12014 0.051
R17855 D.n11998 D.n11996 0.051
R17856 D.n11980 D.n11978 0.051
R17857 D.n11962 D.n11960 0.051
R17858 D.n11944 D.n11942 0.051
R17859 D.n11926 D.n11924 0.051
R17860 D.n11907 D.n11905 0.051
R17861 D.n11917 D.n11916 0.051
R17862 D.n11935 D.n11934 0.051
R17863 D.n11953 D.n11952 0.051
R17864 D.n11971 D.n11970 0.051
R17865 D.n11989 D.n11988 0.051
R17866 D.n12007 D.n12006 0.051
R17867 D.n12025 D.n12024 0.051
R17868 D.n12043 D.n12042 0.051
R17869 D.n12061 D.n12060 0.051
R17870 D.n12079 D.n12078 0.051
R17871 D.n12097 D.n12096 0.051
R17872 D.n12115 D.n12114 0.051
R17873 D.n12133 D.n12132 0.051
R17874 D.n12151 D.n12150 0.051
R17875 D.n12169 D.n12168 0.051
R17876 D.n12187 D.n12186 0.051
R17877 D.n12205 D.n12204 0.051
R17878 D.n12227 D.n12226 0.051
R17879 D.n11516 D.n11514 0.051
R17880 D.n11536 D.n11534 0.051
R17881 D.n11556 D.n11554 0.051
R17882 D.n11576 D.n11574 0.051
R17883 D.n11596 D.n11594 0.051
R17884 D.n11616 D.n11614 0.051
R17885 D.n11636 D.n11634 0.051
R17886 D.n11656 D.n11654 0.051
R17887 D.n11676 D.n11674 0.051
R17888 D.n11696 D.n11694 0.051
R17889 D.n11716 D.n11714 0.051
R17890 D.n11736 D.n11734 0.051
R17891 D.n11756 D.n11754 0.051
R17892 D.n11776 D.n11774 0.051
R17893 D.n11796 D.n11794 0.051
R17894 D.n11816 D.n11814 0.051
R17895 D.n11836 D.n11834 0.051
R17896 D.n11825 D.n11824 0.051
R17897 D.n11805 D.n11804 0.051
R17898 D.n11785 D.n11784 0.051
R17899 D.n11765 D.n11764 0.051
R17900 D.n11745 D.n11744 0.051
R17901 D.n11725 D.n11724 0.051
R17902 D.n11705 D.n11704 0.051
R17903 D.n11685 D.n11684 0.051
R17904 D.n11665 D.n11664 0.051
R17905 D.n11645 D.n11644 0.051
R17906 D.n11625 D.n11624 0.051
R17907 D.n11605 D.n11604 0.051
R17908 D.n11585 D.n11584 0.051
R17909 D.n11565 D.n11564 0.051
R17910 D.n11545 D.n11544 0.051
R17911 D.n11525 D.n11524 0.051
R17912 D.n11502 D.n11501 0.051
R17913 D.n11415 D.n11413 0.051
R17914 D.n11397 D.n11395 0.051
R17915 D.n11379 D.n11377 0.051
R17916 D.n11361 D.n11359 0.051
R17917 D.n11343 D.n11341 0.051
R17918 D.n11325 D.n11323 0.051
R17919 D.n11307 D.n11305 0.051
R17920 D.n11289 D.n11287 0.051
R17921 D.n11271 D.n11269 0.051
R17922 D.n11253 D.n11251 0.051
R17923 D.n11235 D.n11233 0.051
R17924 D.n11217 D.n11215 0.051
R17925 D.n11199 D.n11197 0.051
R17926 D.n11181 D.n11179 0.051
R17927 D.n11163 D.n11161 0.051
R17928 D.n11144 D.n11142 0.051
R17929 D.n11154 D.n11153 0.051
R17930 D.n11172 D.n11171 0.051
R17931 D.n11190 D.n11189 0.051
R17932 D.n11208 D.n11207 0.051
R17933 D.n11226 D.n11225 0.051
R17934 D.n11244 D.n11243 0.051
R17935 D.n11262 D.n11261 0.051
R17936 D.n11280 D.n11279 0.051
R17937 D.n11298 D.n11297 0.051
R17938 D.n11316 D.n11315 0.051
R17939 D.n11334 D.n11333 0.051
R17940 D.n11352 D.n11351 0.051
R17941 D.n11370 D.n11369 0.051
R17942 D.n11388 D.n11387 0.051
R17943 D.n11406 D.n11405 0.051
R17944 D.n11428 D.n11427 0.051
R17945 D.n10793 D.n10791 0.051
R17946 D.n10813 D.n10811 0.051
R17947 D.n10833 D.n10831 0.051
R17948 D.n10853 D.n10851 0.051
R17949 D.n10873 D.n10871 0.051
R17950 D.n10893 D.n10891 0.051
R17951 D.n10913 D.n10911 0.051
R17952 D.n10933 D.n10931 0.051
R17953 D.n10953 D.n10951 0.051
R17954 D.n10973 D.n10971 0.051
R17955 D.n10993 D.n10991 0.051
R17956 D.n11013 D.n11011 0.051
R17957 D.n11033 D.n11031 0.051
R17958 D.n11053 D.n11051 0.051
R17959 D.n11073 D.n11071 0.051
R17960 D.n11062 D.n11061 0.051
R17961 D.n11042 D.n11041 0.051
R17962 D.n11022 D.n11021 0.051
R17963 D.n11002 D.n11001 0.051
R17964 D.n10982 D.n10981 0.051
R17965 D.n10962 D.n10961 0.051
R17966 D.n10942 D.n10941 0.051
R17967 D.n10922 D.n10921 0.051
R17968 D.n10902 D.n10901 0.051
R17969 D.n10882 D.n10881 0.051
R17970 D.n10862 D.n10861 0.051
R17971 D.n10842 D.n10841 0.051
R17972 D.n10822 D.n10821 0.051
R17973 D.n10802 D.n10801 0.051
R17974 D.n10779 D.n10778 0.051
R17975 D.n10696 D.n10694 0.051
R17976 D.n10678 D.n10676 0.051
R17977 D.n10660 D.n10658 0.051
R17978 D.n10642 D.n10640 0.051
R17979 D.n10624 D.n10622 0.051
R17980 D.n10606 D.n10604 0.051
R17981 D.n10588 D.n10586 0.051
R17982 D.n10570 D.n10568 0.051
R17983 D.n10552 D.n10550 0.051
R17984 D.n10534 D.n10532 0.051
R17985 D.n10516 D.n10514 0.051
R17986 D.n10498 D.n10496 0.051
R17987 D.n10480 D.n10478 0.051
R17988 D.n10461 D.n10459 0.051
R17989 D.n10471 D.n10470 0.051
R17990 D.n10489 D.n10488 0.051
R17991 D.n10507 D.n10506 0.051
R17992 D.n10525 D.n10524 0.051
R17993 D.n10543 D.n10542 0.051
R17994 D.n10561 D.n10560 0.051
R17995 D.n10579 D.n10578 0.051
R17996 D.n10597 D.n10596 0.051
R17997 D.n10615 D.n10614 0.051
R17998 D.n10633 D.n10632 0.051
R17999 D.n10651 D.n10650 0.051
R18000 D.n10669 D.n10668 0.051
R18001 D.n10687 D.n10686 0.051
R18002 D.n10709 D.n10708 0.051
R18003 D.n10150 D.n10148 0.051
R18004 D.n10170 D.n10168 0.051
R18005 D.n10190 D.n10188 0.051
R18006 D.n10210 D.n10208 0.051
R18007 D.n10230 D.n10228 0.051
R18008 D.n10250 D.n10248 0.051
R18009 D.n10270 D.n10268 0.051
R18010 D.n10290 D.n10288 0.051
R18011 D.n10310 D.n10308 0.051
R18012 D.n10330 D.n10328 0.051
R18013 D.n10350 D.n10348 0.051
R18014 D.n10370 D.n10368 0.051
R18015 D.n10390 D.n10388 0.051
R18016 D.n10379 D.n10378 0.051
R18017 D.n10359 D.n10358 0.051
R18018 D.n10339 D.n10338 0.051
R18019 D.n10319 D.n10318 0.051
R18020 D.n10299 D.n10298 0.051
R18021 D.n10279 D.n10278 0.051
R18022 D.n10259 D.n10258 0.051
R18023 D.n10239 D.n10238 0.051
R18024 D.n10219 D.n10218 0.051
R18025 D.n10199 D.n10198 0.051
R18026 D.n10179 D.n10178 0.051
R18027 D.n10159 D.n10158 0.051
R18028 D.n10134 D.n10133 0.051
R18029 D.n10057 D.n10055 0.051
R18030 D.n10039 D.n10037 0.051
R18031 D.n10021 D.n10019 0.051
R18032 D.n10003 D.n10001 0.051
R18033 D.n9985 D.n9983 0.051
R18034 D.n9967 D.n9965 0.051
R18035 D.n9949 D.n9947 0.051
R18036 D.n9931 D.n9929 0.051
R18037 D.n9913 D.n9911 0.051
R18038 D.n9895 D.n9893 0.051
R18039 D.n9877 D.n9875 0.051
R18040 D.n9858 D.n9856 0.051
R18041 D.n9868 D.n9867 0.051
R18042 D.n9886 D.n9885 0.051
R18043 D.n9904 D.n9903 0.051
R18044 D.n9922 D.n9921 0.051
R18045 D.n9940 D.n9939 0.051
R18046 D.n9958 D.n9957 0.051
R18047 D.n9976 D.n9975 0.051
R18048 D.n9994 D.n9993 0.051
R18049 D.n10012 D.n10011 0.051
R18050 D.n10030 D.n10029 0.051
R18051 D.n10048 D.n10047 0.051
R18052 D.n10069 D.n10068 0.051
R18053 D.n9587 D.n9585 0.051
R18054 D.n9607 D.n9605 0.051
R18055 D.n9627 D.n9625 0.051
R18056 D.n9647 D.n9645 0.051
R18057 D.n9667 D.n9665 0.051
R18058 D.n9687 D.n9685 0.051
R18059 D.n9707 D.n9705 0.051
R18060 D.n9727 D.n9725 0.051
R18061 D.n9747 D.n9745 0.051
R18062 D.n9767 D.n9765 0.051
R18063 D.n9787 D.n9785 0.051
R18064 D.n9776 D.n9775 0.051
R18065 D.n9756 D.n9755 0.051
R18066 D.n9736 D.n9735 0.051
R18067 D.n9716 D.n9715 0.051
R18068 D.n9696 D.n9695 0.051
R18069 D.n9676 D.n9675 0.051
R18070 D.n9656 D.n9655 0.051
R18071 D.n9636 D.n9635 0.051
R18072 D.n9616 D.n9615 0.051
R18073 D.n9596 D.n9595 0.051
R18074 D.n9571 D.n9570 0.051
R18075 D.n9492 D.n9490 0.051
R18076 D.n9474 D.n9472 0.051
R18077 D.n9456 D.n9454 0.051
R18078 D.n9438 D.n9436 0.051
R18079 D.n9420 D.n9418 0.051
R18080 D.n9402 D.n9400 0.051
R18081 D.n9384 D.n9382 0.051
R18082 D.n9366 D.n9364 0.051
R18083 D.n9348 D.n9346 0.051
R18084 D.n9329 D.n9327 0.051
R18085 D.n9339 D.n9338 0.051
R18086 D.n9357 D.n9356 0.051
R18087 D.n9375 D.n9374 0.051
R18088 D.n9393 D.n9392 0.051
R18089 D.n9411 D.n9410 0.051
R18090 D.n9429 D.n9428 0.051
R18091 D.n9447 D.n9446 0.051
R18092 D.n9465 D.n9464 0.051
R18093 D.n9483 D.n9482 0.051
R18094 D.n9505 D.n9504 0.051
R18095 D.n9098 D.n9096 0.051
R18096 D.n9118 D.n9116 0.051
R18097 D.n9138 D.n9136 0.051
R18098 D.n9158 D.n9156 0.051
R18099 D.n9178 D.n9176 0.051
R18100 D.n9198 D.n9196 0.051
R18101 D.n9218 D.n9216 0.051
R18102 D.n9238 D.n9236 0.051
R18103 D.n9258 D.n9256 0.051
R18104 D.n9247 D.n9246 0.051
R18105 D.n9227 D.n9226 0.051
R18106 D.n9207 D.n9206 0.051
R18107 D.n9187 D.n9186 0.051
R18108 D.n9167 D.n9166 0.051
R18109 D.n9147 D.n9146 0.051
R18110 D.n9127 D.n9126 0.051
R18111 D.n9107 D.n9106 0.051
R18112 D.n9084 D.n9083 0.051
R18113 D.n9013 D.n9011 0.051
R18114 D.n8995 D.n8993 0.051
R18115 D.n8977 D.n8975 0.051
R18116 D.n8959 D.n8957 0.051
R18117 D.n8941 D.n8939 0.051
R18118 D.n8923 D.n8921 0.051
R18119 D.n8905 D.n8903 0.051
R18120 D.n8886 D.n8884 0.051
R18121 D.n8896 D.n8895 0.051
R18122 D.n8914 D.n8913 0.051
R18123 D.n8932 D.n8931 0.051
R18124 D.n8950 D.n8949 0.051
R18125 D.n8968 D.n8967 0.051
R18126 D.n8986 D.n8985 0.051
R18127 D.n9004 D.n9003 0.051
R18128 D.n9026 D.n9025 0.051
R18129 D.n8695 D.n8693 0.051
R18130 D.n8715 D.n8713 0.051
R18131 D.n8735 D.n8733 0.051
R18132 D.n8755 D.n8753 0.051
R18133 D.n8775 D.n8773 0.051
R18134 D.n8795 D.n8793 0.051
R18135 D.n8815 D.n8813 0.051
R18136 D.n8804 D.n8803 0.051
R18137 D.n8784 D.n8783 0.051
R18138 D.n8764 D.n8763 0.051
R18139 D.n8744 D.n8743 0.051
R18140 D.n8724 D.n8723 0.051
R18141 D.n8704 D.n8703 0.051
R18142 D.n8679 D.n8678 0.051
R18143 D.n8614 D.n8612 0.051
R18144 D.n8596 D.n8594 0.051
R18145 D.n8578 D.n8576 0.051
R18146 D.n8560 D.n8558 0.051
R18147 D.n8542 D.n8540 0.051
R18148 D.n8523 D.n8521 0.051
R18149 D.n8533 D.n8532 0.051
R18150 D.n8551 D.n8550 0.051
R18151 D.n8569 D.n8568 0.051
R18152 D.n8587 D.n8586 0.051
R18153 D.n8605 D.n8604 0.051
R18154 D.n8626 D.n8625 0.051
R18155 D.n8372 D.n8370 0.051
R18156 D.n8392 D.n8390 0.051
R18157 D.n8412 D.n8410 0.051
R18158 D.n8432 D.n8430 0.051
R18159 D.n8452 D.n8450 0.051
R18160 D.n8441 D.n8440 0.051
R18161 D.n8421 D.n8420 0.051
R18162 D.n8401 D.n8400 0.051
R18163 D.n8381 D.n8380 0.051
R18164 D.n8356 D.n8355 0.051
R18165 D.n8289 D.n8287 0.051
R18166 D.n8271 D.n8269 0.051
R18167 D.n8253 D.n8251 0.051
R18168 D.n8234 D.n8232 0.051
R18169 D.n8244 D.n8243 0.051
R18170 D.n8262 D.n8261 0.051
R18171 D.n8280 D.n8279 0.051
R18172 D.n8302 D.n8301 0.051
R18173 D.n8123 D.n8121 0.051
R18174 D.n8143 D.n8141 0.051
R18175 D.n8163 D.n8161 0.051
R18176 D.n8152 D.n8151 0.051
R18177 D.n8132 D.n8131 0.051
R18178 D.n8109 D.n8108 0.051
R18179 D.n8050 D.n8048 0.051
R18180 D.n8031 D.n8029 0.051
R18181 D.n8041 D.n8040 0.051
R18182 D.n8063 D.n8062 0.051
R18183 D.n52 D.n51 0.051
R18184 D.n61 D.n60 0.051
R18185 D.n70 D.n69 0.051
R18186 D.n79 D.n78 0.051
R18187 D.n88 D.n87 0.051
R18188 D.n97 D.n96 0.051
R18189 D.n106 D.n105 0.051
R18190 D.n115 D.n114 0.051
R18191 D.n124 D.n123 0.051
R18192 D.n133 D.n132 0.051
R18193 D.n142 D.n141 0.051
R18194 D.n151 D.n150 0.051
R18195 D.n160 D.n159 0.051
R18196 D.n169 D.n168 0.051
R18197 D.n178 D.n177 0.051
R18198 D.n187 D.n186 0.051
R18199 D.n196 D.n195 0.051
R18200 D.n205 D.n204 0.051
R18201 D.n214 D.n213 0.051
R18202 D.n223 D.n222 0.051
R18203 D.n232 D.n231 0.051
R18204 D.n241 D.n240 0.051
R18205 D.n250 D.n249 0.051
R18206 D.n259 D.n258 0.051
R18207 D.n268 D.n267 0.051
R18208 D.n277 D.n276 0.051
R18209 D.n286 D.n285 0.051
R18210 D.n295 D.n294 0.051
R18211 D.n304 D.n303 0.051
R18212 D.n313 D.n312 0.051
R18213 D.n322 D.n321 0.051
R18214 D.n331 D.n330 0.051
R18215 D.n340 D.n339 0.051
R18216 D.n349 D.n348 0.051
R18217 D.n358 D.n357 0.051
R18218 D.n367 D.n366 0.051
R18219 D.n376 D.n375 0.051
R18220 D.n385 D.n384 0.051
R18221 D.n394 D.n393 0.051
R18222 D.n403 D.n402 0.051
R18223 D.n412 D.n411 0.051
R18224 D.n421 D.n420 0.051
R18225 D.n430 D.n429 0.051
R18226 D.n524 D.n522 0.051
R18227 D.n540 D.n538 0.051
R18228 D.n1128 D.n1126 0.051
R18229 D.n1114 D.n1112 0.051
R18230 D.n1100 D.n1098 0.051
R18231 D.n1086 D.n1084 0.051
R18232 D.n1072 D.n1070 0.051
R18233 D.n1058 D.n1056 0.051
R18234 D.n1044 D.n1042 0.051
R18235 D.n1030 D.n1028 0.051
R18236 D.n1016 D.n1014 0.051
R18237 D.n1002 D.n1000 0.051
R18238 D.n988 D.n986 0.051
R18239 D.n974 D.n972 0.051
R18240 D.n960 D.n958 0.051
R18241 D.n946 D.n944 0.051
R18242 D.n932 D.n930 0.051
R18243 D.n918 D.n916 0.051
R18244 D.n904 D.n902 0.051
R18245 D.n890 D.n888 0.051
R18246 D.n876 D.n874 0.051
R18247 D.n862 D.n860 0.051
R18248 D.n848 D.n846 0.051
R18249 D.n834 D.n832 0.051
R18250 D.n820 D.n818 0.051
R18251 D.n806 D.n804 0.051
R18252 D.n792 D.n790 0.051
R18253 D.n778 D.n776 0.051
R18254 D.n764 D.n762 0.051
R18255 D.n750 D.n748 0.051
R18256 D.n736 D.n734 0.051
R18257 D.n722 D.n720 0.051
R18258 D.n708 D.n706 0.051
R18259 D.n694 D.n692 0.051
R18260 D.n680 D.n678 0.051
R18261 D.n666 D.n664 0.051
R18262 D.n652 D.n650 0.051
R18263 D.n638 D.n636 0.051
R18264 D.n624 D.n622 0.051
R18265 D.n610 D.n608 0.051
R18266 D.n596 D.n594 0.051
R18267 D.n582 D.n580 0.051
R18268 D.n568 D.n566 0.051
R18269 D.n554 D.n552 0.051
R18270 D.n1151 D.n1149 0.051
R18271 D.n1167 D.n1165 0.051
R18272 D.n1727 D.n1725 0.051
R18273 D.n1713 D.n1711 0.051
R18274 D.n1699 D.n1697 0.051
R18275 D.n1685 D.n1683 0.051
R18276 D.n1671 D.n1669 0.051
R18277 D.n1657 D.n1655 0.051
R18278 D.n1643 D.n1641 0.051
R18279 D.n1629 D.n1627 0.051
R18280 D.n1615 D.n1613 0.051
R18281 D.n1601 D.n1599 0.051
R18282 D.n1587 D.n1585 0.051
R18283 D.n1573 D.n1571 0.051
R18284 D.n1559 D.n1557 0.051
R18285 D.n1545 D.n1543 0.051
R18286 D.n1531 D.n1529 0.051
R18287 D.n1517 D.n1515 0.051
R18288 D.n1503 D.n1501 0.051
R18289 D.n1489 D.n1487 0.051
R18290 D.n1475 D.n1473 0.051
R18291 D.n1461 D.n1459 0.051
R18292 D.n1447 D.n1445 0.051
R18293 D.n1433 D.n1431 0.051
R18294 D.n1419 D.n1417 0.051
R18295 D.n1405 D.n1403 0.051
R18296 D.n1391 D.n1389 0.051
R18297 D.n1377 D.n1375 0.051
R18298 D.n1363 D.n1361 0.051
R18299 D.n1349 D.n1347 0.051
R18300 D.n1335 D.n1333 0.051
R18301 D.n1321 D.n1319 0.051
R18302 D.n1307 D.n1305 0.051
R18303 D.n1293 D.n1291 0.051
R18304 D.n1279 D.n1277 0.051
R18305 D.n1265 D.n1263 0.051
R18306 D.n1251 D.n1249 0.051
R18307 D.n1237 D.n1235 0.051
R18308 D.n1223 D.n1221 0.051
R18309 D.n1209 D.n1207 0.051
R18310 D.n1195 D.n1193 0.051
R18311 D.n1181 D.n1179 0.051
R18312 D.n1750 D.n1748 0.051
R18313 D.n1766 D.n1764 0.051
R18314 D.n2298 D.n2296 0.051
R18315 D.n2284 D.n2282 0.051
R18316 D.n2270 D.n2268 0.051
R18317 D.n2256 D.n2254 0.051
R18318 D.n2242 D.n2240 0.051
R18319 D.n2228 D.n2226 0.051
R18320 D.n2214 D.n2212 0.051
R18321 D.n2200 D.n2198 0.051
R18322 D.n2186 D.n2184 0.051
R18323 D.n2172 D.n2170 0.051
R18324 D.n2158 D.n2156 0.051
R18325 D.n2144 D.n2142 0.051
R18326 D.n2130 D.n2128 0.051
R18327 D.n2116 D.n2114 0.051
R18328 D.n2102 D.n2100 0.051
R18329 D.n2088 D.n2086 0.051
R18330 D.n2074 D.n2072 0.051
R18331 D.n2060 D.n2058 0.051
R18332 D.n2046 D.n2044 0.051
R18333 D.n2032 D.n2030 0.051
R18334 D.n2018 D.n2016 0.051
R18335 D.n2004 D.n2002 0.051
R18336 D.n1990 D.n1988 0.051
R18337 D.n1976 D.n1974 0.051
R18338 D.n1962 D.n1960 0.051
R18339 D.n1948 D.n1946 0.051
R18340 D.n1934 D.n1932 0.051
R18341 D.n1920 D.n1918 0.051
R18342 D.n1906 D.n1904 0.051
R18343 D.n1892 D.n1890 0.051
R18344 D.n1878 D.n1876 0.051
R18345 D.n1864 D.n1862 0.051
R18346 D.n1850 D.n1848 0.051
R18347 D.n1836 D.n1834 0.051
R18348 D.n1822 D.n1820 0.051
R18349 D.n1808 D.n1806 0.051
R18350 D.n1794 D.n1792 0.051
R18351 D.n1780 D.n1778 0.051
R18352 D.n2321 D.n2319 0.051
R18353 D.n2337 D.n2335 0.051
R18354 D.n2841 D.n2839 0.051
R18355 D.n2827 D.n2825 0.051
R18356 D.n2813 D.n2811 0.051
R18357 D.n2799 D.n2797 0.051
R18358 D.n2785 D.n2783 0.051
R18359 D.n2771 D.n2769 0.051
R18360 D.n2757 D.n2755 0.051
R18361 D.n2743 D.n2741 0.051
R18362 D.n2729 D.n2727 0.051
R18363 D.n2715 D.n2713 0.051
R18364 D.n2701 D.n2699 0.051
R18365 D.n2687 D.n2685 0.051
R18366 D.n2673 D.n2671 0.051
R18367 D.n2659 D.n2657 0.051
R18368 D.n2645 D.n2643 0.051
R18369 D.n2631 D.n2629 0.051
R18370 D.n2617 D.n2615 0.051
R18371 D.n2603 D.n2601 0.051
R18372 D.n2589 D.n2587 0.051
R18373 D.n2575 D.n2573 0.051
R18374 D.n2561 D.n2559 0.051
R18375 D.n2547 D.n2545 0.051
R18376 D.n2533 D.n2531 0.051
R18377 D.n2519 D.n2517 0.051
R18378 D.n2505 D.n2503 0.051
R18379 D.n2491 D.n2489 0.051
R18380 D.n2477 D.n2475 0.051
R18381 D.n2463 D.n2461 0.051
R18382 D.n2449 D.n2447 0.051
R18383 D.n2435 D.n2433 0.051
R18384 D.n2421 D.n2419 0.051
R18385 D.n2407 D.n2405 0.051
R18386 D.n2393 D.n2391 0.051
R18387 D.n2379 D.n2377 0.051
R18388 D.n2365 D.n2363 0.051
R18389 D.n2351 D.n2349 0.051
R18390 D.n2864 D.n2862 0.051
R18391 D.n2880 D.n2878 0.051
R18392 D.n3356 D.n3354 0.051
R18393 D.n3342 D.n3340 0.051
R18394 D.n3328 D.n3326 0.051
R18395 D.n3314 D.n3312 0.051
R18396 D.n3300 D.n3298 0.051
R18397 D.n3286 D.n3284 0.051
R18398 D.n3272 D.n3270 0.051
R18399 D.n3258 D.n3256 0.051
R18400 D.n3244 D.n3242 0.051
R18401 D.n3230 D.n3228 0.051
R18402 D.n3216 D.n3214 0.051
R18403 D.n3202 D.n3200 0.051
R18404 D.n3188 D.n3186 0.051
R18405 D.n3174 D.n3172 0.051
R18406 D.n3160 D.n3158 0.051
R18407 D.n3146 D.n3144 0.051
R18408 D.n3132 D.n3130 0.051
R18409 D.n3118 D.n3116 0.051
R18410 D.n3104 D.n3102 0.051
R18411 D.n3090 D.n3088 0.051
R18412 D.n3076 D.n3074 0.051
R18413 D.n3062 D.n3060 0.051
R18414 D.n3048 D.n3046 0.051
R18415 D.n3034 D.n3032 0.051
R18416 D.n3020 D.n3018 0.051
R18417 D.n3006 D.n3004 0.051
R18418 D.n2992 D.n2990 0.051
R18419 D.n2978 D.n2976 0.051
R18420 D.n2964 D.n2962 0.051
R18421 D.n2950 D.n2948 0.051
R18422 D.n2936 D.n2934 0.051
R18423 D.n2922 D.n2920 0.051
R18424 D.n2908 D.n2906 0.051
R18425 D.n2894 D.n2892 0.051
R18426 D.n3380 D.n3378 0.051
R18427 D.n3396 D.n3394 0.051
R18428 D.n3844 D.n3842 0.051
R18429 D.n3830 D.n3828 0.051
R18430 D.n3816 D.n3814 0.051
R18431 D.n3802 D.n3800 0.051
R18432 D.n3788 D.n3786 0.051
R18433 D.n3774 D.n3772 0.051
R18434 D.n3760 D.n3758 0.051
R18435 D.n3746 D.n3744 0.051
R18436 D.n3732 D.n3730 0.051
R18437 D.n3718 D.n3716 0.051
R18438 D.n3704 D.n3702 0.051
R18439 D.n3690 D.n3688 0.051
R18440 D.n3676 D.n3674 0.051
R18441 D.n3662 D.n3660 0.051
R18442 D.n3648 D.n3646 0.051
R18443 D.n3634 D.n3632 0.051
R18444 D.n3620 D.n3618 0.051
R18445 D.n3606 D.n3604 0.051
R18446 D.n3592 D.n3590 0.051
R18447 D.n3578 D.n3576 0.051
R18448 D.n3564 D.n3562 0.051
R18449 D.n3550 D.n3548 0.051
R18450 D.n3536 D.n3534 0.051
R18451 D.n3522 D.n3520 0.051
R18452 D.n3508 D.n3506 0.051
R18453 D.n3494 D.n3492 0.051
R18454 D.n3480 D.n3478 0.051
R18455 D.n3466 D.n3464 0.051
R18456 D.n3452 D.n3450 0.051
R18457 D.n3438 D.n3436 0.051
R18458 D.n3424 D.n3422 0.051
R18459 D.n3410 D.n3408 0.051
R18460 D.n3868 D.n3866 0.051
R18461 D.n3884 D.n3882 0.051
R18462 D.n4304 D.n4302 0.051
R18463 D.n4290 D.n4288 0.051
R18464 D.n4276 D.n4274 0.051
R18465 D.n4262 D.n4260 0.051
R18466 D.n4248 D.n4246 0.051
R18467 D.n4234 D.n4232 0.051
R18468 D.n4220 D.n4218 0.051
R18469 D.n4206 D.n4204 0.051
R18470 D.n4192 D.n4190 0.051
R18471 D.n4178 D.n4176 0.051
R18472 D.n4164 D.n4162 0.051
R18473 D.n4150 D.n4148 0.051
R18474 D.n4136 D.n4134 0.051
R18475 D.n4122 D.n4120 0.051
R18476 D.n4108 D.n4106 0.051
R18477 D.n4094 D.n4092 0.051
R18478 D.n4080 D.n4078 0.051
R18479 D.n4066 D.n4064 0.051
R18480 D.n4052 D.n4050 0.051
R18481 D.n4038 D.n4036 0.051
R18482 D.n4024 D.n4022 0.051
R18483 D.n4010 D.n4008 0.051
R18484 D.n3996 D.n3994 0.051
R18485 D.n3982 D.n3980 0.051
R18486 D.n3968 D.n3966 0.051
R18487 D.n3954 D.n3952 0.051
R18488 D.n3940 D.n3938 0.051
R18489 D.n3926 D.n3924 0.051
R18490 D.n3912 D.n3910 0.051
R18491 D.n3898 D.n3896 0.051
R18492 D.n4328 D.n4326 0.051
R18493 D.n4344 D.n4342 0.051
R18494 D.n4736 D.n4734 0.051
R18495 D.n4722 D.n4720 0.051
R18496 D.n4708 D.n4706 0.051
R18497 D.n4694 D.n4692 0.051
R18498 D.n4680 D.n4678 0.051
R18499 D.n4666 D.n4664 0.051
R18500 D.n4652 D.n4650 0.051
R18501 D.n4638 D.n4636 0.051
R18502 D.n4624 D.n4622 0.051
R18503 D.n4610 D.n4608 0.051
R18504 D.n4596 D.n4594 0.051
R18505 D.n4582 D.n4580 0.051
R18506 D.n4568 D.n4566 0.051
R18507 D.n4554 D.n4552 0.051
R18508 D.n4540 D.n4538 0.051
R18509 D.n4526 D.n4524 0.051
R18510 D.n4512 D.n4510 0.051
R18511 D.n4498 D.n4496 0.051
R18512 D.n4484 D.n4482 0.051
R18513 D.n4470 D.n4468 0.051
R18514 D.n4456 D.n4454 0.051
R18515 D.n4442 D.n4440 0.051
R18516 D.n4428 D.n4426 0.051
R18517 D.n4414 D.n4412 0.051
R18518 D.n4400 D.n4398 0.051
R18519 D.n4386 D.n4384 0.051
R18520 D.n4372 D.n4370 0.051
R18521 D.n4358 D.n4356 0.051
R18522 D.n4760 D.n4758 0.051
R18523 D.n4776 D.n4774 0.051
R18524 D.n5140 D.n5138 0.051
R18525 D.n5126 D.n5124 0.051
R18526 D.n5112 D.n5110 0.051
R18527 D.n5098 D.n5096 0.051
R18528 D.n5084 D.n5082 0.051
R18529 D.n5070 D.n5068 0.051
R18530 D.n5056 D.n5054 0.051
R18531 D.n5042 D.n5040 0.051
R18532 D.n5028 D.n5026 0.051
R18533 D.n5014 D.n5012 0.051
R18534 D.n5000 D.n4998 0.051
R18535 D.n4986 D.n4984 0.051
R18536 D.n4972 D.n4970 0.051
R18537 D.n4958 D.n4956 0.051
R18538 D.n4944 D.n4942 0.051
R18539 D.n4930 D.n4928 0.051
R18540 D.n4916 D.n4914 0.051
R18541 D.n4902 D.n4900 0.051
R18542 D.n4888 D.n4886 0.051
R18543 D.n4874 D.n4872 0.051
R18544 D.n4860 D.n4858 0.051
R18545 D.n4846 D.n4844 0.051
R18546 D.n4832 D.n4830 0.051
R18547 D.n4818 D.n4816 0.051
R18548 D.n4804 D.n4802 0.051
R18549 D.n4790 D.n4788 0.051
R18550 D.n5164 D.n5162 0.051
R18551 D.n5180 D.n5178 0.051
R18552 D.n5516 D.n5514 0.051
R18553 D.n5502 D.n5500 0.051
R18554 D.n5488 D.n5486 0.051
R18555 D.n5474 D.n5472 0.051
R18556 D.n5460 D.n5458 0.051
R18557 D.n5446 D.n5444 0.051
R18558 D.n5432 D.n5430 0.051
R18559 D.n5418 D.n5416 0.051
R18560 D.n5404 D.n5402 0.051
R18561 D.n5390 D.n5388 0.051
R18562 D.n5376 D.n5374 0.051
R18563 D.n5362 D.n5360 0.051
R18564 D.n5348 D.n5346 0.051
R18565 D.n5334 D.n5332 0.051
R18566 D.n5320 D.n5318 0.051
R18567 D.n5306 D.n5304 0.051
R18568 D.n5292 D.n5290 0.051
R18569 D.n5278 D.n5276 0.051
R18570 D.n5264 D.n5262 0.051
R18571 D.n5250 D.n5248 0.051
R18572 D.n5236 D.n5234 0.051
R18573 D.n5222 D.n5220 0.051
R18574 D.n5208 D.n5206 0.051
R18575 D.n5194 D.n5192 0.051
R18576 D.n5540 D.n5538 0.051
R18577 D.n5556 D.n5554 0.051
R18578 D.n5864 D.n5862 0.051
R18579 D.n5850 D.n5848 0.051
R18580 D.n5836 D.n5834 0.051
R18581 D.n5822 D.n5820 0.051
R18582 D.n5808 D.n5806 0.051
R18583 D.n5794 D.n5792 0.051
R18584 D.n5780 D.n5778 0.051
R18585 D.n5766 D.n5764 0.051
R18586 D.n5752 D.n5750 0.051
R18587 D.n5738 D.n5736 0.051
R18588 D.n5724 D.n5722 0.051
R18589 D.n5710 D.n5708 0.051
R18590 D.n5696 D.n5694 0.051
R18591 D.n5682 D.n5680 0.051
R18592 D.n5668 D.n5666 0.051
R18593 D.n5654 D.n5652 0.051
R18594 D.n5640 D.n5638 0.051
R18595 D.n5626 D.n5624 0.051
R18596 D.n5612 D.n5610 0.051
R18597 D.n5598 D.n5596 0.051
R18598 D.n5584 D.n5582 0.051
R18599 D.n5570 D.n5568 0.051
R18600 D.n5888 D.n5886 0.051
R18601 D.n5904 D.n5902 0.051
R18602 D.n6184 D.n6182 0.051
R18603 D.n6170 D.n6168 0.051
R18604 D.n6156 D.n6154 0.051
R18605 D.n6142 D.n6140 0.051
R18606 D.n6128 D.n6126 0.051
R18607 D.n6114 D.n6112 0.051
R18608 D.n6100 D.n6098 0.051
R18609 D.n6086 D.n6084 0.051
R18610 D.n6072 D.n6070 0.051
R18611 D.n6058 D.n6056 0.051
R18612 D.n6044 D.n6042 0.051
R18613 D.n6030 D.n6028 0.051
R18614 D.n6016 D.n6014 0.051
R18615 D.n6002 D.n6000 0.051
R18616 D.n5988 D.n5986 0.051
R18617 D.n5974 D.n5972 0.051
R18618 D.n5960 D.n5958 0.051
R18619 D.n5946 D.n5944 0.051
R18620 D.n5932 D.n5930 0.051
R18621 D.n5918 D.n5916 0.051
R18622 D.n6208 D.n6206 0.051
R18623 D.n6224 D.n6222 0.051
R18624 D.n6476 D.n6474 0.051
R18625 D.n6462 D.n6460 0.051
R18626 D.n6448 D.n6446 0.051
R18627 D.n6434 D.n6432 0.051
R18628 D.n6420 D.n6418 0.051
R18629 D.n6406 D.n6404 0.051
R18630 D.n6392 D.n6390 0.051
R18631 D.n6378 D.n6376 0.051
R18632 D.n6364 D.n6362 0.051
R18633 D.n6350 D.n6348 0.051
R18634 D.n6336 D.n6334 0.051
R18635 D.n6322 D.n6320 0.051
R18636 D.n6308 D.n6306 0.051
R18637 D.n6294 D.n6292 0.051
R18638 D.n6280 D.n6278 0.051
R18639 D.n6266 D.n6264 0.051
R18640 D.n6252 D.n6250 0.051
R18641 D.n6238 D.n6236 0.051
R18642 D.n6500 D.n6498 0.051
R18643 D.n6516 D.n6514 0.051
R18644 D.n6740 D.n6738 0.051
R18645 D.n6726 D.n6724 0.051
R18646 D.n6712 D.n6710 0.051
R18647 D.n6698 D.n6696 0.051
R18648 D.n6684 D.n6682 0.051
R18649 D.n6670 D.n6668 0.051
R18650 D.n6656 D.n6654 0.051
R18651 D.n6642 D.n6640 0.051
R18652 D.n6628 D.n6626 0.051
R18653 D.n6614 D.n6612 0.051
R18654 D.n6600 D.n6598 0.051
R18655 D.n6586 D.n6584 0.051
R18656 D.n6572 D.n6570 0.051
R18657 D.n6558 D.n6556 0.051
R18658 D.n6544 D.n6542 0.051
R18659 D.n6530 D.n6528 0.051
R18660 D.n6764 D.n6762 0.051
R18661 D.n6780 D.n6778 0.051
R18662 D.n6976 D.n6974 0.051
R18663 D.n6962 D.n6960 0.051
R18664 D.n6948 D.n6946 0.051
R18665 D.n6934 D.n6932 0.051
R18666 D.n6920 D.n6918 0.051
R18667 D.n6906 D.n6904 0.051
R18668 D.n6892 D.n6890 0.051
R18669 D.n6878 D.n6876 0.051
R18670 D.n6864 D.n6862 0.051
R18671 D.n6850 D.n6848 0.051
R18672 D.n6836 D.n6834 0.051
R18673 D.n6822 D.n6820 0.051
R18674 D.n6808 D.n6806 0.051
R18675 D.n6794 D.n6792 0.051
R18676 D.n7000 D.n6998 0.051
R18677 D.n7016 D.n7014 0.051
R18678 D.n7184 D.n7182 0.051
R18679 D.n7170 D.n7168 0.051
R18680 D.n7156 D.n7154 0.051
R18681 D.n7142 D.n7140 0.051
R18682 D.n7128 D.n7126 0.051
R18683 D.n7114 D.n7112 0.051
R18684 D.n7100 D.n7098 0.051
R18685 D.n7086 D.n7084 0.051
R18686 D.n7072 D.n7070 0.051
R18687 D.n7058 D.n7056 0.051
R18688 D.n7044 D.n7042 0.051
R18689 D.n7030 D.n7028 0.051
R18690 D.n7208 D.n7206 0.051
R18691 D.n7224 D.n7222 0.051
R18692 D.n7364 D.n7362 0.051
R18693 D.n7350 D.n7348 0.051
R18694 D.n7336 D.n7334 0.051
R18695 D.n7322 D.n7320 0.051
R18696 D.n7308 D.n7306 0.051
R18697 D.n7294 D.n7292 0.051
R18698 D.n7280 D.n7278 0.051
R18699 D.n7266 D.n7264 0.051
R18700 D.n7252 D.n7250 0.051
R18701 D.n7238 D.n7236 0.051
R18702 D.n7388 D.n7386 0.051
R18703 D.n7404 D.n7402 0.051
R18704 D.n7516 D.n7514 0.051
R18705 D.n7502 D.n7500 0.051
R18706 D.n7488 D.n7486 0.051
R18707 D.n7474 D.n7472 0.051
R18708 D.n7460 D.n7458 0.051
R18709 D.n7446 D.n7444 0.051
R18710 D.n7432 D.n7430 0.051
R18711 D.n7418 D.n7416 0.051
R18712 D.n7540 D.n7538 0.051
R18713 D.n7556 D.n7554 0.051
R18714 D.n7640 D.n7638 0.051
R18715 D.n7626 D.n7624 0.051
R18716 D.n7612 D.n7610 0.051
R18717 D.n7598 D.n7596 0.051
R18718 D.n7584 D.n7582 0.051
R18719 D.n7570 D.n7568 0.051
R18720 D.n7664 D.n7662 0.051
R18721 D.n7680 D.n7678 0.051
R18722 D.n7736 D.n7734 0.051
R18723 D.n7722 D.n7720 0.051
R18724 D.n7708 D.n7706 0.051
R18725 D.n7694 D.n7692 0.051
R18726 D.n7759 D.n7757 0.051
R18727 D.n7775 D.n7773 0.051
R18728 D.n7803 D.n7801 0.051
R18729 D.n7789 D.n7787 0.051
R18730 D.n7890 D.n7889 0.051
R18731 D.n7856 D.n7852 0.05
R18732 D.n7849 D.n7819 0.05
R18733 D.n7933 D.n7929 0.05
R18734 D.n14096 D.n14089 0.05
R18735 D.n13183 D.n13179 0.05
R18736 D.n13127 D.n13122 0.05
R18737 D.n12300 D.n12296 0.05
R18738 D.n12248 D.n12241 0.05
R18739 D.n11495 D.n11492 0.05
R18740 D.n11449 D.n11442 0.05
R18741 D.n10772 D.n10769 0.05
R18742 D.n10730 D.n10723 0.05
R18743 D.n10125 D.n10121 0.05
R18744 D.n10085 D.n10080 0.05
R18745 D.n9562 D.n9558 0.05
R18746 D.n9526 D.n9519 0.05
R18747 D.n9077 D.n9074 0.05
R18748 D.n9047 D.n9040 0.05
R18749 D.n8670 D.n8666 0.05
R18750 D.n8642 D.n8637 0.05
R18751 D.n8347 D.n8343 0.05
R18752 D.n8323 D.n8316 0.05
R18753 D.n8102 D.n8099 0.05
R18754 D.n8084 D.n8077 0.05
R18755 D.n7917 D.n7911 0.05
R18756 D.n1141 D.n515 0.05
R18757 D.n1740 D.n1145 0.05
R18758 D.n2311 D.n1744 0.05
R18759 D.n2854 D.n2315 0.05
R18760 D.n3369 D.n2858 0.05
R18761 D.n3857 D.n3374 0.05
R18762 D.n4317 D.n3862 0.05
R18763 D.n4749 D.n4322 0.05
R18764 D.n5153 D.n4754 0.05
R18765 D.n5529 D.n5158 0.05
R18766 D.n5877 D.n5534 0.05
R18767 D.n6197 D.n5882 0.05
R18768 D.n6489 D.n6202 0.05
R18769 D.n6753 D.n6494 0.05
R18770 D.n6989 D.n6758 0.05
R18771 D.n7197 D.n6994 0.05
R18772 D.n7377 D.n7202 0.05
R18773 D.n7529 D.n7382 0.05
R18774 D.n7653 D.n7534 0.05
R18775 D.n7749 D.n7658 0.05
R18776 D.n7816 D.n7753 0.05
R18777 D.n1138 D.n1124 0.049
R18778 D.n1124 D.n1110 0.049
R18779 D.n1110 D.n1096 0.049
R18780 D.n1096 D.n1082 0.049
R18781 D.n1082 D.n1068 0.049
R18782 D.n1068 D.n1054 0.049
R18783 D.n1054 D.n1040 0.049
R18784 D.n1040 D.n1026 0.049
R18785 D.n1026 D.n1012 0.049
R18786 D.n1012 D.n998 0.049
R18787 D.n998 D.n984 0.049
R18788 D.n984 D.n970 0.049
R18789 D.n970 D.n956 0.049
R18790 D.n956 D.n942 0.049
R18791 D.n942 D.n928 0.049
R18792 D.n928 D.n914 0.049
R18793 D.n914 D.n900 0.049
R18794 D.n900 D.n886 0.049
R18795 D.n886 D.n872 0.049
R18796 D.n872 D.n858 0.049
R18797 D.n858 D.n844 0.049
R18798 D.n844 D.n830 0.049
R18799 D.n830 D.n816 0.049
R18800 D.n816 D.n802 0.049
R18801 D.n802 D.n788 0.049
R18802 D.n788 D.n774 0.049
R18803 D.n774 D.n760 0.049
R18804 D.n760 D.n746 0.049
R18805 D.n746 D.n732 0.049
R18806 D.n732 D.n718 0.049
R18807 D.n718 D.n704 0.049
R18808 D.n704 D.n690 0.049
R18809 D.n690 D.n676 0.049
R18810 D.n676 D.n662 0.049
R18811 D.n662 D.n648 0.049
R18812 D.n648 D.n634 0.049
R18813 D.n634 D.n620 0.049
R18814 D.n620 D.n606 0.049
R18815 D.n606 D.n592 0.049
R18816 D.n592 D.n578 0.049
R18817 D.n578 D.n564 0.049
R18818 D.n564 D.n550 0.049
R18819 D.n550 D.n536 0.049
R18820 D.n1737 D.n1723 0.049
R18821 D.n1723 D.n1709 0.049
R18822 D.n1709 D.n1695 0.049
R18823 D.n1695 D.n1681 0.049
R18824 D.n1681 D.n1667 0.049
R18825 D.n1667 D.n1653 0.049
R18826 D.n1653 D.n1639 0.049
R18827 D.n1639 D.n1625 0.049
R18828 D.n1625 D.n1611 0.049
R18829 D.n1611 D.n1597 0.049
R18830 D.n1597 D.n1583 0.049
R18831 D.n1583 D.n1569 0.049
R18832 D.n1569 D.n1555 0.049
R18833 D.n1555 D.n1541 0.049
R18834 D.n1541 D.n1527 0.049
R18835 D.n1527 D.n1513 0.049
R18836 D.n1513 D.n1499 0.049
R18837 D.n1499 D.n1485 0.049
R18838 D.n1485 D.n1471 0.049
R18839 D.n1471 D.n1457 0.049
R18840 D.n1457 D.n1443 0.049
R18841 D.n1443 D.n1429 0.049
R18842 D.n1429 D.n1415 0.049
R18843 D.n1415 D.n1401 0.049
R18844 D.n1401 D.n1387 0.049
R18845 D.n1387 D.n1373 0.049
R18846 D.n1373 D.n1359 0.049
R18847 D.n1359 D.n1345 0.049
R18848 D.n1345 D.n1331 0.049
R18849 D.n1331 D.n1317 0.049
R18850 D.n1317 D.n1303 0.049
R18851 D.n1303 D.n1289 0.049
R18852 D.n1289 D.n1275 0.049
R18853 D.n1275 D.n1261 0.049
R18854 D.n1261 D.n1247 0.049
R18855 D.n1247 D.n1233 0.049
R18856 D.n1233 D.n1219 0.049
R18857 D.n1219 D.n1205 0.049
R18858 D.n1205 D.n1191 0.049
R18859 D.n1191 D.n1177 0.049
R18860 D.n1177 D.n1163 0.049
R18861 D.n2308 D.n2294 0.049
R18862 D.n2294 D.n2280 0.049
R18863 D.n2280 D.n2266 0.049
R18864 D.n2266 D.n2252 0.049
R18865 D.n2252 D.n2238 0.049
R18866 D.n2238 D.n2224 0.049
R18867 D.n2224 D.n2210 0.049
R18868 D.n2210 D.n2196 0.049
R18869 D.n2196 D.n2182 0.049
R18870 D.n2182 D.n2168 0.049
R18871 D.n2168 D.n2154 0.049
R18872 D.n2154 D.n2140 0.049
R18873 D.n2140 D.n2126 0.049
R18874 D.n2126 D.n2112 0.049
R18875 D.n2112 D.n2098 0.049
R18876 D.n2098 D.n2084 0.049
R18877 D.n2084 D.n2070 0.049
R18878 D.n2070 D.n2056 0.049
R18879 D.n2056 D.n2042 0.049
R18880 D.n2042 D.n2028 0.049
R18881 D.n2028 D.n2014 0.049
R18882 D.n2014 D.n2000 0.049
R18883 D.n2000 D.n1986 0.049
R18884 D.n1986 D.n1972 0.049
R18885 D.n1972 D.n1958 0.049
R18886 D.n1958 D.n1944 0.049
R18887 D.n1944 D.n1930 0.049
R18888 D.n1930 D.n1916 0.049
R18889 D.n1916 D.n1902 0.049
R18890 D.n1902 D.n1888 0.049
R18891 D.n1888 D.n1874 0.049
R18892 D.n1874 D.n1860 0.049
R18893 D.n1860 D.n1846 0.049
R18894 D.n1846 D.n1832 0.049
R18895 D.n1832 D.n1818 0.049
R18896 D.n1818 D.n1804 0.049
R18897 D.n1804 D.n1790 0.049
R18898 D.n1790 D.n1776 0.049
R18899 D.n1776 D.n1762 0.049
R18900 D.n2851 D.n2837 0.049
R18901 D.n2837 D.n2823 0.049
R18902 D.n2823 D.n2809 0.049
R18903 D.n2809 D.n2795 0.049
R18904 D.n2795 D.n2781 0.049
R18905 D.n2781 D.n2767 0.049
R18906 D.n2767 D.n2753 0.049
R18907 D.n2753 D.n2739 0.049
R18908 D.n2739 D.n2725 0.049
R18909 D.n2725 D.n2711 0.049
R18910 D.n2711 D.n2697 0.049
R18911 D.n2697 D.n2683 0.049
R18912 D.n2683 D.n2669 0.049
R18913 D.n2669 D.n2655 0.049
R18914 D.n2655 D.n2641 0.049
R18915 D.n2641 D.n2627 0.049
R18916 D.n2627 D.n2613 0.049
R18917 D.n2613 D.n2599 0.049
R18918 D.n2599 D.n2585 0.049
R18919 D.n2585 D.n2571 0.049
R18920 D.n2571 D.n2557 0.049
R18921 D.n2557 D.n2543 0.049
R18922 D.n2543 D.n2529 0.049
R18923 D.n2529 D.n2515 0.049
R18924 D.n2515 D.n2501 0.049
R18925 D.n2501 D.n2487 0.049
R18926 D.n2487 D.n2473 0.049
R18927 D.n2473 D.n2459 0.049
R18928 D.n2459 D.n2445 0.049
R18929 D.n2445 D.n2431 0.049
R18930 D.n2431 D.n2417 0.049
R18931 D.n2417 D.n2403 0.049
R18932 D.n2403 D.n2389 0.049
R18933 D.n2389 D.n2375 0.049
R18934 D.n2375 D.n2361 0.049
R18935 D.n2361 D.n2347 0.049
R18936 D.n2347 D.n2333 0.049
R18937 D.n3366 D.n3352 0.049
R18938 D.n3352 D.n3338 0.049
R18939 D.n3338 D.n3324 0.049
R18940 D.n3324 D.n3310 0.049
R18941 D.n3310 D.n3296 0.049
R18942 D.n3296 D.n3282 0.049
R18943 D.n3282 D.n3268 0.049
R18944 D.n3268 D.n3254 0.049
R18945 D.n3254 D.n3240 0.049
R18946 D.n3240 D.n3226 0.049
R18947 D.n3226 D.n3212 0.049
R18948 D.n3212 D.n3198 0.049
R18949 D.n3198 D.n3184 0.049
R18950 D.n3184 D.n3170 0.049
R18951 D.n3170 D.n3156 0.049
R18952 D.n3156 D.n3142 0.049
R18953 D.n3142 D.n3128 0.049
R18954 D.n3128 D.n3114 0.049
R18955 D.n3114 D.n3100 0.049
R18956 D.n3100 D.n3086 0.049
R18957 D.n3086 D.n3072 0.049
R18958 D.n3072 D.n3058 0.049
R18959 D.n3058 D.n3044 0.049
R18960 D.n3044 D.n3030 0.049
R18961 D.n3030 D.n3016 0.049
R18962 D.n3016 D.n3002 0.049
R18963 D.n3002 D.n2988 0.049
R18964 D.n2988 D.n2974 0.049
R18965 D.n2974 D.n2960 0.049
R18966 D.n2960 D.n2946 0.049
R18967 D.n2946 D.n2932 0.049
R18968 D.n2932 D.n2918 0.049
R18969 D.n2918 D.n2904 0.049
R18970 D.n2904 D.n2890 0.049
R18971 D.n2890 D.n2876 0.049
R18972 D.n3854 D.n3840 0.049
R18973 D.n3840 D.n3826 0.049
R18974 D.n3826 D.n3812 0.049
R18975 D.n3812 D.n3798 0.049
R18976 D.n3798 D.n3784 0.049
R18977 D.n3784 D.n3770 0.049
R18978 D.n3770 D.n3756 0.049
R18979 D.n3756 D.n3742 0.049
R18980 D.n3742 D.n3728 0.049
R18981 D.n3728 D.n3714 0.049
R18982 D.n3714 D.n3700 0.049
R18983 D.n3700 D.n3686 0.049
R18984 D.n3686 D.n3672 0.049
R18985 D.n3672 D.n3658 0.049
R18986 D.n3658 D.n3644 0.049
R18987 D.n3644 D.n3630 0.049
R18988 D.n3630 D.n3616 0.049
R18989 D.n3616 D.n3602 0.049
R18990 D.n3602 D.n3588 0.049
R18991 D.n3588 D.n3574 0.049
R18992 D.n3574 D.n3560 0.049
R18993 D.n3560 D.n3546 0.049
R18994 D.n3546 D.n3532 0.049
R18995 D.n3532 D.n3518 0.049
R18996 D.n3518 D.n3504 0.049
R18997 D.n3504 D.n3490 0.049
R18998 D.n3490 D.n3476 0.049
R18999 D.n3476 D.n3462 0.049
R19000 D.n3462 D.n3448 0.049
R19001 D.n3448 D.n3434 0.049
R19002 D.n3434 D.n3420 0.049
R19003 D.n3420 D.n3406 0.049
R19004 D.n3406 D.n3392 0.049
R19005 D.n4314 D.n4300 0.049
R19006 D.n4300 D.n4286 0.049
R19007 D.n4286 D.n4272 0.049
R19008 D.n4272 D.n4258 0.049
R19009 D.n4258 D.n4244 0.049
R19010 D.n4244 D.n4230 0.049
R19011 D.n4230 D.n4216 0.049
R19012 D.n4216 D.n4202 0.049
R19013 D.n4202 D.n4188 0.049
R19014 D.n4188 D.n4174 0.049
R19015 D.n4174 D.n4160 0.049
R19016 D.n4160 D.n4146 0.049
R19017 D.n4146 D.n4132 0.049
R19018 D.n4132 D.n4118 0.049
R19019 D.n4118 D.n4104 0.049
R19020 D.n4104 D.n4090 0.049
R19021 D.n4090 D.n4076 0.049
R19022 D.n4076 D.n4062 0.049
R19023 D.n4062 D.n4048 0.049
R19024 D.n4048 D.n4034 0.049
R19025 D.n4034 D.n4020 0.049
R19026 D.n4020 D.n4006 0.049
R19027 D.n4006 D.n3992 0.049
R19028 D.n3992 D.n3978 0.049
R19029 D.n3978 D.n3964 0.049
R19030 D.n3964 D.n3950 0.049
R19031 D.n3950 D.n3936 0.049
R19032 D.n3936 D.n3922 0.049
R19033 D.n3922 D.n3908 0.049
R19034 D.n3908 D.n3894 0.049
R19035 D.n3894 D.n3880 0.049
R19036 D.n4746 D.n4732 0.049
R19037 D.n4732 D.n4718 0.049
R19038 D.n4718 D.n4704 0.049
R19039 D.n4704 D.n4690 0.049
R19040 D.n4690 D.n4676 0.049
R19041 D.n4676 D.n4662 0.049
R19042 D.n4662 D.n4648 0.049
R19043 D.n4648 D.n4634 0.049
R19044 D.n4634 D.n4620 0.049
R19045 D.n4620 D.n4606 0.049
R19046 D.n4606 D.n4592 0.049
R19047 D.n4592 D.n4578 0.049
R19048 D.n4578 D.n4564 0.049
R19049 D.n4564 D.n4550 0.049
R19050 D.n4550 D.n4536 0.049
R19051 D.n4536 D.n4522 0.049
R19052 D.n4522 D.n4508 0.049
R19053 D.n4508 D.n4494 0.049
R19054 D.n4494 D.n4480 0.049
R19055 D.n4480 D.n4466 0.049
R19056 D.n4466 D.n4452 0.049
R19057 D.n4452 D.n4438 0.049
R19058 D.n4438 D.n4424 0.049
R19059 D.n4424 D.n4410 0.049
R19060 D.n4410 D.n4396 0.049
R19061 D.n4396 D.n4382 0.049
R19062 D.n4382 D.n4368 0.049
R19063 D.n4368 D.n4354 0.049
R19064 D.n4354 D.n4340 0.049
R19065 D.n5150 D.n5136 0.049
R19066 D.n5136 D.n5122 0.049
R19067 D.n5122 D.n5108 0.049
R19068 D.n5108 D.n5094 0.049
R19069 D.n5094 D.n5080 0.049
R19070 D.n5080 D.n5066 0.049
R19071 D.n5066 D.n5052 0.049
R19072 D.n5052 D.n5038 0.049
R19073 D.n5038 D.n5024 0.049
R19074 D.n5024 D.n5010 0.049
R19075 D.n5010 D.n4996 0.049
R19076 D.n4996 D.n4982 0.049
R19077 D.n4982 D.n4968 0.049
R19078 D.n4968 D.n4954 0.049
R19079 D.n4954 D.n4940 0.049
R19080 D.n4940 D.n4926 0.049
R19081 D.n4926 D.n4912 0.049
R19082 D.n4912 D.n4898 0.049
R19083 D.n4898 D.n4884 0.049
R19084 D.n4884 D.n4870 0.049
R19085 D.n4870 D.n4856 0.049
R19086 D.n4856 D.n4842 0.049
R19087 D.n4842 D.n4828 0.049
R19088 D.n4828 D.n4814 0.049
R19089 D.n4814 D.n4800 0.049
R19090 D.n4800 D.n4786 0.049
R19091 D.n4786 D.n4772 0.049
R19092 D.n5526 D.n5512 0.049
R19093 D.n5512 D.n5498 0.049
R19094 D.n5498 D.n5484 0.049
R19095 D.n5484 D.n5470 0.049
R19096 D.n5470 D.n5456 0.049
R19097 D.n5456 D.n5442 0.049
R19098 D.n5442 D.n5428 0.049
R19099 D.n5428 D.n5414 0.049
R19100 D.n5414 D.n5400 0.049
R19101 D.n5400 D.n5386 0.049
R19102 D.n5386 D.n5372 0.049
R19103 D.n5372 D.n5358 0.049
R19104 D.n5358 D.n5344 0.049
R19105 D.n5344 D.n5330 0.049
R19106 D.n5330 D.n5316 0.049
R19107 D.n5316 D.n5302 0.049
R19108 D.n5302 D.n5288 0.049
R19109 D.n5288 D.n5274 0.049
R19110 D.n5274 D.n5260 0.049
R19111 D.n5260 D.n5246 0.049
R19112 D.n5246 D.n5232 0.049
R19113 D.n5232 D.n5218 0.049
R19114 D.n5218 D.n5204 0.049
R19115 D.n5204 D.n5190 0.049
R19116 D.n5190 D.n5176 0.049
R19117 D.n5874 D.n5860 0.049
R19118 D.n5860 D.n5846 0.049
R19119 D.n5846 D.n5832 0.049
R19120 D.n5832 D.n5818 0.049
R19121 D.n5818 D.n5804 0.049
R19122 D.n5804 D.n5790 0.049
R19123 D.n5790 D.n5776 0.049
R19124 D.n5776 D.n5762 0.049
R19125 D.n5762 D.n5748 0.049
R19126 D.n5748 D.n5734 0.049
R19127 D.n5734 D.n5720 0.049
R19128 D.n5720 D.n5706 0.049
R19129 D.n5706 D.n5692 0.049
R19130 D.n5692 D.n5678 0.049
R19131 D.n5678 D.n5664 0.049
R19132 D.n5664 D.n5650 0.049
R19133 D.n5650 D.n5636 0.049
R19134 D.n5636 D.n5622 0.049
R19135 D.n5622 D.n5608 0.049
R19136 D.n5608 D.n5594 0.049
R19137 D.n5594 D.n5580 0.049
R19138 D.n5580 D.n5566 0.049
R19139 D.n5566 D.n5552 0.049
R19140 D.n6194 D.n6180 0.049
R19141 D.n6180 D.n6166 0.049
R19142 D.n6166 D.n6152 0.049
R19143 D.n6152 D.n6138 0.049
R19144 D.n6138 D.n6124 0.049
R19145 D.n6124 D.n6110 0.049
R19146 D.n6110 D.n6096 0.049
R19147 D.n6096 D.n6082 0.049
R19148 D.n6082 D.n6068 0.049
R19149 D.n6068 D.n6054 0.049
R19150 D.n6054 D.n6040 0.049
R19151 D.n6040 D.n6026 0.049
R19152 D.n6026 D.n6012 0.049
R19153 D.n6012 D.n5998 0.049
R19154 D.n5998 D.n5984 0.049
R19155 D.n5984 D.n5970 0.049
R19156 D.n5970 D.n5956 0.049
R19157 D.n5956 D.n5942 0.049
R19158 D.n5942 D.n5928 0.049
R19159 D.n5928 D.n5914 0.049
R19160 D.n5914 D.n5900 0.049
R19161 D.n6486 D.n6472 0.049
R19162 D.n6472 D.n6458 0.049
R19163 D.n6458 D.n6444 0.049
R19164 D.n6444 D.n6430 0.049
R19165 D.n6430 D.n6416 0.049
R19166 D.n6416 D.n6402 0.049
R19167 D.n6402 D.n6388 0.049
R19168 D.n6388 D.n6374 0.049
R19169 D.n6374 D.n6360 0.049
R19170 D.n6360 D.n6346 0.049
R19171 D.n6346 D.n6332 0.049
R19172 D.n6332 D.n6318 0.049
R19173 D.n6318 D.n6304 0.049
R19174 D.n6304 D.n6290 0.049
R19175 D.n6290 D.n6276 0.049
R19176 D.n6276 D.n6262 0.049
R19177 D.n6262 D.n6248 0.049
R19178 D.n6248 D.n6234 0.049
R19179 D.n6234 D.n6220 0.049
R19180 D.n6750 D.n6736 0.049
R19181 D.n6736 D.n6722 0.049
R19182 D.n6722 D.n6708 0.049
R19183 D.n6708 D.n6694 0.049
R19184 D.n6694 D.n6680 0.049
R19185 D.n6680 D.n6666 0.049
R19186 D.n6666 D.n6652 0.049
R19187 D.n6652 D.n6638 0.049
R19188 D.n6638 D.n6624 0.049
R19189 D.n6624 D.n6610 0.049
R19190 D.n6610 D.n6596 0.049
R19191 D.n6596 D.n6582 0.049
R19192 D.n6582 D.n6568 0.049
R19193 D.n6568 D.n6554 0.049
R19194 D.n6554 D.n6540 0.049
R19195 D.n6540 D.n6526 0.049
R19196 D.n6526 D.n6512 0.049
R19197 D.n6986 D.n6972 0.049
R19198 D.n6972 D.n6958 0.049
R19199 D.n6958 D.n6944 0.049
R19200 D.n6944 D.n6930 0.049
R19201 D.n6930 D.n6916 0.049
R19202 D.n6916 D.n6902 0.049
R19203 D.n6902 D.n6888 0.049
R19204 D.n6888 D.n6874 0.049
R19205 D.n6874 D.n6860 0.049
R19206 D.n6860 D.n6846 0.049
R19207 D.n6846 D.n6832 0.049
R19208 D.n6832 D.n6818 0.049
R19209 D.n6818 D.n6804 0.049
R19210 D.n6804 D.n6790 0.049
R19211 D.n6790 D.n6776 0.049
R19212 D.n7194 D.n7180 0.049
R19213 D.n7180 D.n7166 0.049
R19214 D.n7166 D.n7152 0.049
R19215 D.n7152 D.n7138 0.049
R19216 D.n7138 D.n7124 0.049
R19217 D.n7124 D.n7110 0.049
R19218 D.n7110 D.n7096 0.049
R19219 D.n7096 D.n7082 0.049
R19220 D.n7082 D.n7068 0.049
R19221 D.n7068 D.n7054 0.049
R19222 D.n7054 D.n7040 0.049
R19223 D.n7040 D.n7026 0.049
R19224 D.n7026 D.n7012 0.049
R19225 D.n7374 D.n7360 0.049
R19226 D.n7360 D.n7346 0.049
R19227 D.n7346 D.n7332 0.049
R19228 D.n7332 D.n7318 0.049
R19229 D.n7318 D.n7304 0.049
R19230 D.n7304 D.n7290 0.049
R19231 D.n7290 D.n7276 0.049
R19232 D.n7276 D.n7262 0.049
R19233 D.n7262 D.n7248 0.049
R19234 D.n7248 D.n7234 0.049
R19235 D.n7234 D.n7220 0.049
R19236 D.n7526 D.n7512 0.049
R19237 D.n7512 D.n7498 0.049
R19238 D.n7498 D.n7484 0.049
R19239 D.n7484 D.n7470 0.049
R19240 D.n7470 D.n7456 0.049
R19241 D.n7456 D.n7442 0.049
R19242 D.n7442 D.n7428 0.049
R19243 D.n7428 D.n7414 0.049
R19244 D.n7414 D.n7400 0.049
R19245 D.n7650 D.n7636 0.049
R19246 D.n7636 D.n7622 0.049
R19247 D.n7622 D.n7608 0.049
R19248 D.n7608 D.n7594 0.049
R19249 D.n7594 D.n7580 0.049
R19250 D.n7580 D.n7566 0.049
R19251 D.n7566 D.n7552 0.049
R19252 D.n7746 D.n7732 0.049
R19253 D.n7732 D.n7718 0.049
R19254 D.n7718 D.n7704 0.049
R19255 D.n7704 D.n7690 0.049
R19256 D.n7690 D.n7676 0.049
R19257 D.n7815 D.n7799 0.049
R19258 D.n7799 D.n7785 0.049
R19259 D.n7785 D.n7771 0.049
R19260 D.n12 D.n11 0.049
R19261 D.n457 D.n456 0.049
R19262 D.n458 D.n457 0.049
R19263 D.n459 D.n458 0.049
R19264 D.n460 D.n459 0.049
R19265 D.n461 D.n460 0.049
R19266 D.n462 D.n461 0.049
R19267 D.n463 D.n462 0.049
R19268 D.n464 D.n463 0.049
R19269 D.n465 D.n464 0.049
R19270 D.n466 D.n465 0.049
R19271 D.n467 D.n466 0.049
R19272 D.n468 D.n467 0.049
R19273 D.n469 D.n468 0.049
R19274 D.n470 D.n469 0.049
R19275 D.n471 D.n470 0.049
R19276 D.n472 D.n471 0.049
R19277 D.n473 D.n472 0.049
R19278 D.n474 D.n473 0.049
R19279 D.n475 D.n474 0.049
R19280 D.n476 D.n475 0.049
R19281 D.n477 D.n476 0.049
R19282 D.n478 D.n477 0.049
R19283 D.n479 D.n478 0.049
R19284 D.n480 D.n479 0.049
R19285 D.n481 D.n480 0.049
R19286 D.n482 D.n481 0.049
R19287 D.n483 D.n482 0.049
R19288 D.n484 D.n483 0.049
R19289 D.n485 D.n484 0.049
R19290 D.n486 D.n485 0.049
R19291 D.n487 D.n486 0.049
R19292 D.n488 D.n487 0.049
R19293 D.n489 D.n488 0.049
R19294 D.n490 D.n489 0.049
R19295 D.n491 D.n490 0.049
R19296 D.n492 D.n491 0.049
R19297 D.n493 D.n492 0.049
R19298 D.n494 D.n493 0.049
R19299 D.n495 D.n494 0.049
R19300 D.n496 D.n495 0.049
R19301 D.n497 D.n496 0.049
R19302 D.n498 D.n497 0.049
R19303 D.n499 D.n498 0.049
R19304 D.n500 D.n499 0.049
R19305 D.n501 D.n500 0.049
R19306 D.n14098 D.n14097 0.049
R19307 D.n14099 D.n14098 0.049
R19308 D.n14100 D.n14099 0.049
R19309 D.n14101 D.n14100 0.049
R19310 D.n14102 D.n14101 0.049
R19311 D.n14103 D.n14102 0.049
R19312 D.n14104 D.n14103 0.049
R19313 D.n14105 D.n14104 0.049
R19314 D.n14106 D.n14105 0.049
R19315 D.n14107 D.n14106 0.049
R19316 D.n14108 D.n14107 0.049
R19317 D.n14109 D.n14108 0.049
R19318 D.n14110 D.n14109 0.049
R19319 D.n14111 D.n14110 0.049
R19320 D.n14112 D.n14111 0.049
R19321 D.n14113 D.n14112 0.049
R19322 D.n14114 D.n14113 0.049
R19323 D.n14115 D.n14114 0.049
R19324 D.n14116 D.n14115 0.049
R19325 D.n14117 D.n14116 0.049
R19326 D.n14118 D.n14117 0.049
R19327 D.n14119 D.n14118 0.049
R19328 D.n14120 D.n14119 0.049
R19329 D.n14121 D.n14120 0.049
R19330 D.n14122 D.n14121 0.049
R19331 D.n14123 D.n14122 0.049
R19332 D.n14124 D.n14123 0.049
R19333 D.n14125 D.n14124 0.049
R19334 D.n14126 D.n14125 0.049
R19335 D.n14127 D.n14126 0.049
R19336 D.n14128 D.n14127 0.049
R19337 D.n14129 D.n14128 0.049
R19338 D.n14130 D.n14129 0.049
R19339 D.n14131 D.n14130 0.049
R19340 D.n14132 D.n14131 0.049
R19341 D.n14133 D.n14132 0.049
R19342 D.n14134 D.n14133 0.049
R19343 D.n14135 D.n14134 0.049
R19344 D.n14136 D.n14135 0.049
R19345 D.n14137 D.n14136 0.049
R19346 D.n14138 D.n14137 0.049
R19347 D.n14139 D.n14138 0.049
R19348 D.n14140 D.n14139 0.049
R19349 D.n13129 D.n13128 0.049
R19350 D.n13130 D.n13129 0.049
R19351 D.n13131 D.n13130 0.049
R19352 D.n13132 D.n13131 0.049
R19353 D.n13133 D.n13132 0.049
R19354 D.n13134 D.n13133 0.049
R19355 D.n13135 D.n13134 0.049
R19356 D.n13136 D.n13135 0.049
R19357 D.n13137 D.n13136 0.049
R19358 D.n13138 D.n13137 0.049
R19359 D.n13139 D.n13138 0.049
R19360 D.n13140 D.n13139 0.049
R19361 D.n13141 D.n13140 0.049
R19362 D.n13142 D.n13141 0.049
R19363 D.n13143 D.n13142 0.049
R19364 D.n13144 D.n13143 0.049
R19365 D.n13145 D.n13144 0.049
R19366 D.n13146 D.n13145 0.049
R19367 D.n13147 D.n13146 0.049
R19368 D.n13148 D.n13147 0.049
R19369 D.n13149 D.n13148 0.049
R19370 D.n13150 D.n13149 0.049
R19371 D.n13151 D.n13150 0.049
R19372 D.n13152 D.n13151 0.049
R19373 D.n13153 D.n13152 0.049
R19374 D.n13154 D.n13153 0.049
R19375 D.n13155 D.n13154 0.049
R19376 D.n13156 D.n13155 0.049
R19377 D.n13157 D.n13156 0.049
R19378 D.n13158 D.n13157 0.049
R19379 D.n13159 D.n13158 0.049
R19380 D.n13160 D.n13159 0.049
R19381 D.n13161 D.n13160 0.049
R19382 D.n13162 D.n13161 0.049
R19383 D.n13163 D.n13162 0.049
R19384 D.n13164 D.n13163 0.049
R19385 D.n13165 D.n13164 0.049
R19386 D.n13166 D.n13165 0.049
R19387 D.n13167 D.n13166 0.049
R19388 D.n12250 D.n12249 0.049
R19389 D.n12251 D.n12250 0.049
R19390 D.n12252 D.n12251 0.049
R19391 D.n12253 D.n12252 0.049
R19392 D.n12254 D.n12253 0.049
R19393 D.n12255 D.n12254 0.049
R19394 D.n12256 D.n12255 0.049
R19395 D.n12257 D.n12256 0.049
R19396 D.n12258 D.n12257 0.049
R19397 D.n12259 D.n12258 0.049
R19398 D.n12260 D.n12259 0.049
R19399 D.n12261 D.n12260 0.049
R19400 D.n12262 D.n12261 0.049
R19401 D.n12263 D.n12262 0.049
R19402 D.n12264 D.n12263 0.049
R19403 D.n12265 D.n12264 0.049
R19404 D.n12266 D.n12265 0.049
R19405 D.n12267 D.n12266 0.049
R19406 D.n12268 D.n12267 0.049
R19407 D.n12269 D.n12268 0.049
R19408 D.n12270 D.n12269 0.049
R19409 D.n12271 D.n12270 0.049
R19410 D.n12272 D.n12271 0.049
R19411 D.n12273 D.n12272 0.049
R19412 D.n12274 D.n12273 0.049
R19413 D.n12275 D.n12274 0.049
R19414 D.n12276 D.n12275 0.049
R19415 D.n12277 D.n12276 0.049
R19416 D.n12278 D.n12277 0.049
R19417 D.n12279 D.n12278 0.049
R19418 D.n12280 D.n12279 0.049
R19419 D.n12281 D.n12280 0.049
R19420 D.n12282 D.n12281 0.049
R19421 D.n12283 D.n12282 0.049
R19422 D.n12284 D.n12283 0.049
R19423 D.n11451 D.n11450 0.049
R19424 D.n11452 D.n11451 0.049
R19425 D.n11453 D.n11452 0.049
R19426 D.n11454 D.n11453 0.049
R19427 D.n11455 D.n11454 0.049
R19428 D.n11456 D.n11455 0.049
R19429 D.n11457 D.n11456 0.049
R19430 D.n11458 D.n11457 0.049
R19431 D.n11459 D.n11458 0.049
R19432 D.n11460 D.n11459 0.049
R19433 D.n11461 D.n11460 0.049
R19434 D.n11462 D.n11461 0.049
R19435 D.n11463 D.n11462 0.049
R19436 D.n11464 D.n11463 0.049
R19437 D.n11465 D.n11464 0.049
R19438 D.n11466 D.n11465 0.049
R19439 D.n11467 D.n11466 0.049
R19440 D.n11468 D.n11467 0.049
R19441 D.n11469 D.n11468 0.049
R19442 D.n11470 D.n11469 0.049
R19443 D.n11471 D.n11470 0.049
R19444 D.n11472 D.n11471 0.049
R19445 D.n11473 D.n11472 0.049
R19446 D.n11474 D.n11473 0.049
R19447 D.n11475 D.n11474 0.049
R19448 D.n11476 D.n11475 0.049
R19449 D.n11477 D.n11476 0.049
R19450 D.n11478 D.n11477 0.049
R19451 D.n11479 D.n11478 0.049
R19452 D.n11480 D.n11479 0.049
R19453 D.n11481 D.n11480 0.049
R19454 D.n10732 D.n10731 0.049
R19455 D.n10733 D.n10732 0.049
R19456 D.n10734 D.n10733 0.049
R19457 D.n10735 D.n10734 0.049
R19458 D.n10736 D.n10735 0.049
R19459 D.n10737 D.n10736 0.049
R19460 D.n10738 D.n10737 0.049
R19461 D.n10739 D.n10738 0.049
R19462 D.n10740 D.n10739 0.049
R19463 D.n10741 D.n10740 0.049
R19464 D.n10742 D.n10741 0.049
R19465 D.n10743 D.n10742 0.049
R19466 D.n10744 D.n10743 0.049
R19467 D.n10745 D.n10744 0.049
R19468 D.n10746 D.n10745 0.049
R19469 D.n10747 D.n10746 0.049
R19470 D.n10748 D.n10747 0.049
R19471 D.n10749 D.n10748 0.049
R19472 D.n10750 D.n10749 0.049
R19473 D.n10751 D.n10750 0.049
R19474 D.n10752 D.n10751 0.049
R19475 D.n10753 D.n10752 0.049
R19476 D.n10754 D.n10753 0.049
R19477 D.n10755 D.n10754 0.049
R19478 D.n10756 D.n10755 0.049
R19479 D.n10757 D.n10756 0.049
R19480 D.n10758 D.n10757 0.049
R19481 D.n10087 D.n10086 0.049
R19482 D.n10088 D.n10087 0.049
R19483 D.n10089 D.n10088 0.049
R19484 D.n10090 D.n10089 0.049
R19485 D.n10091 D.n10090 0.049
R19486 D.n10092 D.n10091 0.049
R19487 D.n10093 D.n10092 0.049
R19488 D.n10094 D.n10093 0.049
R19489 D.n10095 D.n10094 0.049
R19490 D.n10096 D.n10095 0.049
R19491 D.n10097 D.n10096 0.049
R19492 D.n10098 D.n10097 0.049
R19493 D.n10099 D.n10098 0.049
R19494 D.n10100 D.n10099 0.049
R19495 D.n10101 D.n10100 0.049
R19496 D.n10102 D.n10101 0.049
R19497 D.n10103 D.n10102 0.049
R19498 D.n10104 D.n10103 0.049
R19499 D.n10105 D.n10104 0.049
R19500 D.n10106 D.n10105 0.049
R19501 D.n10107 D.n10106 0.049
R19502 D.n10108 D.n10107 0.049
R19503 D.n10109 D.n10108 0.049
R19504 D.n9528 D.n9527 0.049
R19505 D.n9529 D.n9528 0.049
R19506 D.n9530 D.n9529 0.049
R19507 D.n9531 D.n9530 0.049
R19508 D.n9532 D.n9531 0.049
R19509 D.n9533 D.n9532 0.049
R19510 D.n9534 D.n9533 0.049
R19511 D.n9535 D.n9534 0.049
R19512 D.n9536 D.n9535 0.049
R19513 D.n9537 D.n9536 0.049
R19514 D.n9538 D.n9537 0.049
R19515 D.n9539 D.n9538 0.049
R19516 D.n9540 D.n9539 0.049
R19517 D.n9541 D.n9540 0.049
R19518 D.n9542 D.n9541 0.049
R19519 D.n9543 D.n9542 0.049
R19520 D.n9544 D.n9543 0.049
R19521 D.n9545 D.n9544 0.049
R19522 D.n9546 D.n9545 0.049
R19523 D.n9049 D.n9048 0.049
R19524 D.n9050 D.n9049 0.049
R19525 D.n9051 D.n9050 0.049
R19526 D.n9052 D.n9051 0.049
R19527 D.n9053 D.n9052 0.049
R19528 D.n9054 D.n9053 0.049
R19529 D.n9055 D.n9054 0.049
R19530 D.n9056 D.n9055 0.049
R19531 D.n9057 D.n9056 0.049
R19532 D.n9058 D.n9057 0.049
R19533 D.n9059 D.n9058 0.049
R19534 D.n9060 D.n9059 0.049
R19535 D.n9061 D.n9060 0.049
R19536 D.n9062 D.n9061 0.049
R19537 D.n9063 D.n9062 0.049
R19538 D.n8644 D.n8643 0.049
R19539 D.n8645 D.n8644 0.049
R19540 D.n8646 D.n8645 0.049
R19541 D.n8647 D.n8646 0.049
R19542 D.n8648 D.n8647 0.049
R19543 D.n8649 D.n8648 0.049
R19544 D.n8650 D.n8649 0.049
R19545 D.n8651 D.n8650 0.049
R19546 D.n8652 D.n8651 0.049
R19547 D.n8653 D.n8652 0.049
R19548 D.n8654 D.n8653 0.049
R19549 D.n8325 D.n8324 0.049
R19550 D.n8326 D.n8325 0.049
R19551 D.n8327 D.n8326 0.049
R19552 D.n8328 D.n8327 0.049
R19553 D.n8329 D.n8328 0.049
R19554 D.n8330 D.n8329 0.049
R19555 D.n8331 D.n8330 0.049
R19556 D.n8086 D.n8085 0.049
R19557 D.n8087 D.n8086 0.049
R19558 D.n8088 D.n8087 0.049
R19559 D.n14141 D.n14140 0.049
R19560 D.n13168 D.n13167 0.049
R19561 D.n12285 D.n12284 0.049
R19562 D.n11482 D.n11481 0.049
R19563 D.n10759 D.n10758 0.049
R19564 D.n10110 D.n10109 0.049
R19565 D.n9547 D.n9546 0.049
R19566 D.n9064 D.n9063 0.049
R19567 D.n8655 D.n8654 0.049
R19568 D.n8332 D.n8331 0.049
R19569 D.n8089 D.n8088 0.049
R19570 D.n1141 D.n1138 0.047
R19571 D.n1740 D.n1737 0.047
R19572 D.n2311 D.n2308 0.047
R19573 D.n2854 D.n2851 0.047
R19574 D.n3369 D.n3366 0.047
R19575 D.n3857 D.n3854 0.047
R19576 D.n4317 D.n4314 0.047
R19577 D.n4749 D.n4746 0.047
R19578 D.n5153 D.n5150 0.047
R19579 D.n5529 D.n5526 0.047
R19580 D.n5877 D.n5874 0.047
R19581 D.n6197 D.n6194 0.047
R19582 D.n6489 D.n6486 0.047
R19583 D.n6753 D.n6750 0.047
R19584 D.n6989 D.n6986 0.047
R19585 D.n7197 D.n7194 0.047
R19586 D.n7377 D.n7374 0.047
R19587 D.n7529 D.n7526 0.047
R19588 D.n7653 D.n7650 0.047
R19589 D.n7749 D.n7746 0.047
R19590 D.n7816 D.n7815 0.047
R19591 D.n7897 D.n7896 0.045
R19592 D.n7980 D.n7979 0.045
R19593 D.n13647 D.n13646 0.045
R19594 D.n13663 D.n13662 0.045
R19595 D.n13616 D.n13615 0.045
R19596 D.n13628 D.n13627 0.045
R19597 D.n12724 D.n12723 0.045
R19598 D.n12740 D.n12739 0.045
R19599 D.n12693 D.n12692 0.045
R19600 D.n12705 D.n12704 0.045
R19601 D.n11875 D.n11874 0.045
R19602 D.n11891 D.n11890 0.045
R19603 D.n11844 D.n11843 0.045
R19604 D.n11856 D.n11855 0.045
R19605 D.n11112 D.n11111 0.045
R19606 D.n11128 D.n11127 0.045
R19607 D.n11081 D.n11080 0.045
R19608 D.n11093 D.n11092 0.045
R19609 D.n10429 D.n10428 0.045
R19610 D.n10445 D.n10444 0.045
R19611 D.n10398 D.n10397 0.045
R19612 D.n10410 D.n10409 0.045
R19613 D.n9826 D.n9825 0.045
R19614 D.n9842 D.n9841 0.045
R19615 D.n9795 D.n9794 0.045
R19616 D.n9807 D.n9806 0.045
R19617 D.n9297 D.n9296 0.045
R19618 D.n9313 D.n9312 0.045
R19619 D.n9266 D.n9265 0.045
R19620 D.n9278 D.n9277 0.045
R19621 D.n8854 D.n8853 0.045
R19622 D.n8870 D.n8869 0.045
R19623 D.n8823 D.n8822 0.045
R19624 D.n8835 D.n8834 0.045
R19625 D.n8491 D.n8490 0.045
R19626 D.n8507 D.n8506 0.045
R19627 D.n8460 D.n8459 0.045
R19628 D.n8472 D.n8471 0.045
R19629 D.n8202 D.n8201 0.045
R19630 D.n8218 D.n8217 0.045
R19631 D.n8171 D.n8170 0.045
R19632 D.n8183 D.n8182 0.045
R19633 D.n7999 D.n7998 0.045
R19634 D.n8015 D.n8014 0.045
R19635 D.n7966 D.n7965 0.045
R19636 D.n7890 D.n7887 0.044
R19637 D.n502 D.n501 0.044
R19638 D.n7950 D.n7949 0.043
R19639 D.n13200 D.n13199 0.043
R19640 D.n12317 D.n12316 0.043
R19641 D.n12236 D.n12235 0.043
R19642 D.n11508 D.n11507 0.043
R19643 D.n11437 D.n11436 0.043
R19644 D.n10785 D.n10784 0.043
R19645 D.n10718 D.n10717 0.043
R19646 D.n10142 D.n10141 0.043
R19647 D.n9579 D.n9578 0.043
R19648 D.n9514 D.n9513 0.043
R19649 D.n9090 D.n9089 0.043
R19650 D.n9035 D.n9034 0.043
R19651 D.n8687 D.n8686 0.043
R19652 D.n8364 D.n8363 0.043
R19653 D.n8311 D.n8310 0.043
R19654 D.n8115 D.n8114 0.043
R19655 D.n8072 D.n8071 0.043
R19656 D.n14071 D.n14070 0.043
R19657 D.n13188 D.n13187 0.043
R19658 D.n13107 D.n13106 0.043
R19659 D.n12305 D.n12304 0.043
R19660 D.n12223 D.n12222 0.043
R19661 D.n11498 D.n11497 0.043
R19662 D.n11424 D.n11423 0.043
R19663 D.n10775 D.n10774 0.043
R19664 D.n10705 D.n10704 0.043
R19665 D.n10130 D.n10129 0.043
R19666 D.n10065 D.n10064 0.043
R19667 D.n9567 D.n9566 0.043
R19668 D.n9501 D.n9500 0.043
R19669 D.n9080 D.n9079 0.043
R19670 D.n9022 D.n9021 0.043
R19671 D.n8675 D.n8674 0.043
R19672 D.n8622 D.n8621 0.043
R19673 D.n8352 D.n8351 0.043
R19674 D.n8298 D.n8297 0.043
R19675 D.n8105 D.n8104 0.043
R19676 D.n8059 D.n8058 0.043
R19677 D.n7938 D.n7937 0.043
R19678 D.n549 D.n548 0.042
R19679 D.n563 D.n562 0.042
R19680 D.n577 D.n576 0.042
R19681 D.n591 D.n590 0.042
R19682 D.n605 D.n604 0.042
R19683 D.n619 D.n618 0.042
R19684 D.n633 D.n632 0.042
R19685 D.n647 D.n646 0.042
R19686 D.n661 D.n660 0.042
R19687 D.n675 D.n674 0.042
R19688 D.n689 D.n688 0.042
R19689 D.n703 D.n702 0.042
R19690 D.n717 D.n716 0.042
R19691 D.n731 D.n730 0.042
R19692 D.n745 D.n744 0.042
R19693 D.n759 D.n758 0.042
R19694 D.n773 D.n772 0.042
R19695 D.n787 D.n786 0.042
R19696 D.n801 D.n800 0.042
R19697 D.n815 D.n814 0.042
R19698 D.n829 D.n828 0.042
R19699 D.n843 D.n842 0.042
R19700 D.n857 D.n856 0.042
R19701 D.n871 D.n870 0.042
R19702 D.n885 D.n884 0.042
R19703 D.n899 D.n898 0.042
R19704 D.n913 D.n912 0.042
R19705 D.n927 D.n926 0.042
R19706 D.n941 D.n940 0.042
R19707 D.n955 D.n954 0.042
R19708 D.n969 D.n968 0.042
R19709 D.n983 D.n982 0.042
R19710 D.n997 D.n996 0.042
R19711 D.n1011 D.n1010 0.042
R19712 D.n1025 D.n1024 0.042
R19713 D.n1039 D.n1038 0.042
R19714 D.n1053 D.n1052 0.042
R19715 D.n1067 D.n1066 0.042
R19716 D.n1081 D.n1080 0.042
R19717 D.n1095 D.n1094 0.042
R19718 D.n1109 D.n1108 0.042
R19719 D.n1123 D.n1122 0.042
R19720 D.n1137 D.n1136 0.042
R19721 D.n1176 D.n1175 0.042
R19722 D.n1190 D.n1189 0.042
R19723 D.n1204 D.n1203 0.042
R19724 D.n1218 D.n1217 0.042
R19725 D.n1232 D.n1231 0.042
R19726 D.n1246 D.n1245 0.042
R19727 D.n1260 D.n1259 0.042
R19728 D.n1274 D.n1273 0.042
R19729 D.n1288 D.n1287 0.042
R19730 D.n1302 D.n1301 0.042
R19731 D.n1316 D.n1315 0.042
R19732 D.n1330 D.n1329 0.042
R19733 D.n1344 D.n1343 0.042
R19734 D.n1358 D.n1357 0.042
R19735 D.n1372 D.n1371 0.042
R19736 D.n1386 D.n1385 0.042
R19737 D.n1400 D.n1399 0.042
R19738 D.n1414 D.n1413 0.042
R19739 D.n1428 D.n1427 0.042
R19740 D.n1442 D.n1441 0.042
R19741 D.n1456 D.n1455 0.042
R19742 D.n1470 D.n1469 0.042
R19743 D.n1484 D.n1483 0.042
R19744 D.n1498 D.n1497 0.042
R19745 D.n1512 D.n1511 0.042
R19746 D.n1526 D.n1525 0.042
R19747 D.n1540 D.n1539 0.042
R19748 D.n1554 D.n1553 0.042
R19749 D.n1568 D.n1567 0.042
R19750 D.n1582 D.n1581 0.042
R19751 D.n1596 D.n1595 0.042
R19752 D.n1610 D.n1609 0.042
R19753 D.n1624 D.n1623 0.042
R19754 D.n1638 D.n1637 0.042
R19755 D.n1652 D.n1651 0.042
R19756 D.n1666 D.n1665 0.042
R19757 D.n1680 D.n1679 0.042
R19758 D.n1694 D.n1693 0.042
R19759 D.n1708 D.n1707 0.042
R19760 D.n1722 D.n1721 0.042
R19761 D.n1736 D.n1735 0.042
R19762 D.n1775 D.n1774 0.042
R19763 D.n1789 D.n1788 0.042
R19764 D.n1803 D.n1802 0.042
R19765 D.n1817 D.n1816 0.042
R19766 D.n1831 D.n1830 0.042
R19767 D.n1845 D.n1844 0.042
R19768 D.n1859 D.n1858 0.042
R19769 D.n1873 D.n1872 0.042
R19770 D.n1887 D.n1886 0.042
R19771 D.n1901 D.n1900 0.042
R19772 D.n1915 D.n1914 0.042
R19773 D.n1929 D.n1928 0.042
R19774 D.n1943 D.n1942 0.042
R19775 D.n1957 D.n1956 0.042
R19776 D.n1971 D.n1970 0.042
R19777 D.n1985 D.n1984 0.042
R19778 D.n1999 D.n1998 0.042
R19779 D.n2013 D.n2012 0.042
R19780 D.n2027 D.n2026 0.042
R19781 D.n2041 D.n2040 0.042
R19782 D.n2055 D.n2054 0.042
R19783 D.n2069 D.n2068 0.042
R19784 D.n2083 D.n2082 0.042
R19785 D.n2097 D.n2096 0.042
R19786 D.n2111 D.n2110 0.042
R19787 D.n2125 D.n2124 0.042
R19788 D.n2139 D.n2138 0.042
R19789 D.n2153 D.n2152 0.042
R19790 D.n2167 D.n2166 0.042
R19791 D.n2181 D.n2180 0.042
R19792 D.n2195 D.n2194 0.042
R19793 D.n2209 D.n2208 0.042
R19794 D.n2223 D.n2222 0.042
R19795 D.n2237 D.n2236 0.042
R19796 D.n2251 D.n2250 0.042
R19797 D.n2265 D.n2264 0.042
R19798 D.n2279 D.n2278 0.042
R19799 D.n2293 D.n2292 0.042
R19800 D.n2307 D.n2306 0.042
R19801 D.n2346 D.n2345 0.042
R19802 D.n2360 D.n2359 0.042
R19803 D.n2374 D.n2373 0.042
R19804 D.n2388 D.n2387 0.042
R19805 D.n2402 D.n2401 0.042
R19806 D.n2416 D.n2415 0.042
R19807 D.n2430 D.n2429 0.042
R19808 D.n2444 D.n2443 0.042
R19809 D.n2458 D.n2457 0.042
R19810 D.n2472 D.n2471 0.042
R19811 D.n2486 D.n2485 0.042
R19812 D.n2500 D.n2499 0.042
R19813 D.n2514 D.n2513 0.042
R19814 D.n2528 D.n2527 0.042
R19815 D.n2542 D.n2541 0.042
R19816 D.n2556 D.n2555 0.042
R19817 D.n2570 D.n2569 0.042
R19818 D.n2584 D.n2583 0.042
R19819 D.n2598 D.n2597 0.042
R19820 D.n2612 D.n2611 0.042
R19821 D.n2626 D.n2625 0.042
R19822 D.n2640 D.n2639 0.042
R19823 D.n2654 D.n2653 0.042
R19824 D.n2668 D.n2667 0.042
R19825 D.n2682 D.n2681 0.042
R19826 D.n2696 D.n2695 0.042
R19827 D.n2710 D.n2709 0.042
R19828 D.n2724 D.n2723 0.042
R19829 D.n2738 D.n2737 0.042
R19830 D.n2752 D.n2751 0.042
R19831 D.n2766 D.n2765 0.042
R19832 D.n2780 D.n2779 0.042
R19833 D.n2794 D.n2793 0.042
R19834 D.n2808 D.n2807 0.042
R19835 D.n2822 D.n2821 0.042
R19836 D.n2836 D.n2835 0.042
R19837 D.n2850 D.n2849 0.042
R19838 D.n2889 D.n2888 0.042
R19839 D.n2903 D.n2902 0.042
R19840 D.n2917 D.n2916 0.042
R19841 D.n2931 D.n2930 0.042
R19842 D.n2945 D.n2944 0.042
R19843 D.n2959 D.n2958 0.042
R19844 D.n2973 D.n2972 0.042
R19845 D.n2987 D.n2986 0.042
R19846 D.n3001 D.n3000 0.042
R19847 D.n3015 D.n3014 0.042
R19848 D.n3029 D.n3028 0.042
R19849 D.n3043 D.n3042 0.042
R19850 D.n3057 D.n3056 0.042
R19851 D.n3071 D.n3070 0.042
R19852 D.n3085 D.n3084 0.042
R19853 D.n3099 D.n3098 0.042
R19854 D.n3113 D.n3112 0.042
R19855 D.n3127 D.n3126 0.042
R19856 D.n3141 D.n3140 0.042
R19857 D.n3155 D.n3154 0.042
R19858 D.n3169 D.n3168 0.042
R19859 D.n3183 D.n3182 0.042
R19860 D.n3197 D.n3196 0.042
R19861 D.n3211 D.n3210 0.042
R19862 D.n3225 D.n3224 0.042
R19863 D.n3239 D.n3238 0.042
R19864 D.n3253 D.n3252 0.042
R19865 D.n3267 D.n3266 0.042
R19866 D.n3281 D.n3280 0.042
R19867 D.n3295 D.n3294 0.042
R19868 D.n3309 D.n3308 0.042
R19869 D.n3323 D.n3322 0.042
R19870 D.n3337 D.n3336 0.042
R19871 D.n3351 D.n3350 0.042
R19872 D.n3365 D.n3364 0.042
R19873 D.n3405 D.n3404 0.042
R19874 D.n3419 D.n3418 0.042
R19875 D.n3433 D.n3432 0.042
R19876 D.n3447 D.n3446 0.042
R19877 D.n3461 D.n3460 0.042
R19878 D.n3475 D.n3474 0.042
R19879 D.n3489 D.n3488 0.042
R19880 D.n3503 D.n3502 0.042
R19881 D.n3517 D.n3516 0.042
R19882 D.n3531 D.n3530 0.042
R19883 D.n3545 D.n3544 0.042
R19884 D.n3559 D.n3558 0.042
R19885 D.n3573 D.n3572 0.042
R19886 D.n3587 D.n3586 0.042
R19887 D.n3601 D.n3600 0.042
R19888 D.n3615 D.n3614 0.042
R19889 D.n3629 D.n3628 0.042
R19890 D.n3643 D.n3642 0.042
R19891 D.n3657 D.n3656 0.042
R19892 D.n3671 D.n3670 0.042
R19893 D.n3685 D.n3684 0.042
R19894 D.n3699 D.n3698 0.042
R19895 D.n3713 D.n3712 0.042
R19896 D.n3727 D.n3726 0.042
R19897 D.n3741 D.n3740 0.042
R19898 D.n3755 D.n3754 0.042
R19899 D.n3769 D.n3768 0.042
R19900 D.n3783 D.n3782 0.042
R19901 D.n3797 D.n3796 0.042
R19902 D.n3811 D.n3810 0.042
R19903 D.n3825 D.n3824 0.042
R19904 D.n3839 D.n3838 0.042
R19905 D.n3853 D.n3852 0.042
R19906 D.n3893 D.n3892 0.042
R19907 D.n3907 D.n3906 0.042
R19908 D.n3921 D.n3920 0.042
R19909 D.n3935 D.n3934 0.042
R19910 D.n3949 D.n3948 0.042
R19911 D.n3963 D.n3962 0.042
R19912 D.n3977 D.n3976 0.042
R19913 D.n3991 D.n3990 0.042
R19914 D.n4005 D.n4004 0.042
R19915 D.n4019 D.n4018 0.042
R19916 D.n4033 D.n4032 0.042
R19917 D.n4047 D.n4046 0.042
R19918 D.n4061 D.n4060 0.042
R19919 D.n4075 D.n4074 0.042
R19920 D.n4089 D.n4088 0.042
R19921 D.n4103 D.n4102 0.042
R19922 D.n4117 D.n4116 0.042
R19923 D.n4131 D.n4130 0.042
R19924 D.n4145 D.n4144 0.042
R19925 D.n4159 D.n4158 0.042
R19926 D.n4173 D.n4172 0.042
R19927 D.n4187 D.n4186 0.042
R19928 D.n4201 D.n4200 0.042
R19929 D.n4215 D.n4214 0.042
R19930 D.n4229 D.n4228 0.042
R19931 D.n4243 D.n4242 0.042
R19932 D.n4257 D.n4256 0.042
R19933 D.n4271 D.n4270 0.042
R19934 D.n4285 D.n4284 0.042
R19935 D.n4299 D.n4298 0.042
R19936 D.n4313 D.n4312 0.042
R19937 D.n4353 D.n4352 0.042
R19938 D.n4367 D.n4366 0.042
R19939 D.n4381 D.n4380 0.042
R19940 D.n4395 D.n4394 0.042
R19941 D.n4409 D.n4408 0.042
R19942 D.n4423 D.n4422 0.042
R19943 D.n4437 D.n4436 0.042
R19944 D.n4451 D.n4450 0.042
R19945 D.n4465 D.n4464 0.042
R19946 D.n4479 D.n4478 0.042
R19947 D.n4493 D.n4492 0.042
R19948 D.n4507 D.n4506 0.042
R19949 D.n4521 D.n4520 0.042
R19950 D.n4535 D.n4534 0.042
R19951 D.n4549 D.n4548 0.042
R19952 D.n4563 D.n4562 0.042
R19953 D.n4577 D.n4576 0.042
R19954 D.n4591 D.n4590 0.042
R19955 D.n4605 D.n4604 0.042
R19956 D.n4619 D.n4618 0.042
R19957 D.n4633 D.n4632 0.042
R19958 D.n4647 D.n4646 0.042
R19959 D.n4661 D.n4660 0.042
R19960 D.n4675 D.n4674 0.042
R19961 D.n4689 D.n4688 0.042
R19962 D.n4703 D.n4702 0.042
R19963 D.n4717 D.n4716 0.042
R19964 D.n4731 D.n4730 0.042
R19965 D.n4745 D.n4744 0.042
R19966 D.n4785 D.n4784 0.042
R19967 D.n4799 D.n4798 0.042
R19968 D.n4813 D.n4812 0.042
R19969 D.n4827 D.n4826 0.042
R19970 D.n4841 D.n4840 0.042
R19971 D.n4855 D.n4854 0.042
R19972 D.n4869 D.n4868 0.042
R19973 D.n4883 D.n4882 0.042
R19974 D.n4897 D.n4896 0.042
R19975 D.n4911 D.n4910 0.042
R19976 D.n4925 D.n4924 0.042
R19977 D.n4939 D.n4938 0.042
R19978 D.n4953 D.n4952 0.042
R19979 D.n4967 D.n4966 0.042
R19980 D.n4981 D.n4980 0.042
R19981 D.n4995 D.n4994 0.042
R19982 D.n5009 D.n5008 0.042
R19983 D.n5023 D.n5022 0.042
R19984 D.n5037 D.n5036 0.042
R19985 D.n5051 D.n5050 0.042
R19986 D.n5065 D.n5064 0.042
R19987 D.n5079 D.n5078 0.042
R19988 D.n5093 D.n5092 0.042
R19989 D.n5107 D.n5106 0.042
R19990 D.n5121 D.n5120 0.042
R19991 D.n5135 D.n5134 0.042
R19992 D.n5149 D.n5148 0.042
R19993 D.n5189 D.n5188 0.042
R19994 D.n5203 D.n5202 0.042
R19995 D.n5217 D.n5216 0.042
R19996 D.n5231 D.n5230 0.042
R19997 D.n5245 D.n5244 0.042
R19998 D.n5259 D.n5258 0.042
R19999 D.n5273 D.n5272 0.042
R20000 D.n5287 D.n5286 0.042
R20001 D.n5301 D.n5300 0.042
R20002 D.n5315 D.n5314 0.042
R20003 D.n5329 D.n5328 0.042
R20004 D.n5343 D.n5342 0.042
R20005 D.n5357 D.n5356 0.042
R20006 D.n5371 D.n5370 0.042
R20007 D.n5385 D.n5384 0.042
R20008 D.n5399 D.n5398 0.042
R20009 D.n5413 D.n5412 0.042
R20010 D.n5427 D.n5426 0.042
R20011 D.n5441 D.n5440 0.042
R20012 D.n5455 D.n5454 0.042
R20013 D.n5469 D.n5468 0.042
R20014 D.n5483 D.n5482 0.042
R20015 D.n5497 D.n5496 0.042
R20016 D.n5511 D.n5510 0.042
R20017 D.n5525 D.n5524 0.042
R20018 D.n5565 D.n5564 0.042
R20019 D.n5579 D.n5578 0.042
R20020 D.n5593 D.n5592 0.042
R20021 D.n5607 D.n5606 0.042
R20022 D.n5621 D.n5620 0.042
R20023 D.n5635 D.n5634 0.042
R20024 D.n5649 D.n5648 0.042
R20025 D.n5663 D.n5662 0.042
R20026 D.n5677 D.n5676 0.042
R20027 D.n5691 D.n5690 0.042
R20028 D.n5705 D.n5704 0.042
R20029 D.n5719 D.n5718 0.042
R20030 D.n5733 D.n5732 0.042
R20031 D.n5747 D.n5746 0.042
R20032 D.n5761 D.n5760 0.042
R20033 D.n5775 D.n5774 0.042
R20034 D.n5789 D.n5788 0.042
R20035 D.n5803 D.n5802 0.042
R20036 D.n5817 D.n5816 0.042
R20037 D.n5831 D.n5830 0.042
R20038 D.n5845 D.n5844 0.042
R20039 D.n5859 D.n5858 0.042
R20040 D.n5873 D.n5872 0.042
R20041 D.n5913 D.n5912 0.042
R20042 D.n5927 D.n5926 0.042
R20043 D.n5941 D.n5940 0.042
R20044 D.n5955 D.n5954 0.042
R20045 D.n5969 D.n5968 0.042
R20046 D.n5983 D.n5982 0.042
R20047 D.n5997 D.n5996 0.042
R20048 D.n6011 D.n6010 0.042
R20049 D.n6025 D.n6024 0.042
R20050 D.n6039 D.n6038 0.042
R20051 D.n6053 D.n6052 0.042
R20052 D.n6067 D.n6066 0.042
R20053 D.n6081 D.n6080 0.042
R20054 D.n6095 D.n6094 0.042
R20055 D.n6109 D.n6108 0.042
R20056 D.n6123 D.n6122 0.042
R20057 D.n6137 D.n6136 0.042
R20058 D.n6151 D.n6150 0.042
R20059 D.n6165 D.n6164 0.042
R20060 D.n6179 D.n6178 0.042
R20061 D.n6193 D.n6192 0.042
R20062 D.n6233 D.n6232 0.042
R20063 D.n6247 D.n6246 0.042
R20064 D.n6261 D.n6260 0.042
R20065 D.n6275 D.n6274 0.042
R20066 D.n6289 D.n6288 0.042
R20067 D.n6303 D.n6302 0.042
R20068 D.n6317 D.n6316 0.042
R20069 D.n6331 D.n6330 0.042
R20070 D.n6345 D.n6344 0.042
R20071 D.n6359 D.n6358 0.042
R20072 D.n6373 D.n6372 0.042
R20073 D.n6387 D.n6386 0.042
R20074 D.n6401 D.n6400 0.042
R20075 D.n6415 D.n6414 0.042
R20076 D.n6429 D.n6428 0.042
R20077 D.n6443 D.n6442 0.042
R20078 D.n6457 D.n6456 0.042
R20079 D.n6471 D.n6470 0.042
R20080 D.n6485 D.n6484 0.042
R20081 D.n6525 D.n6524 0.042
R20082 D.n6539 D.n6538 0.042
R20083 D.n6553 D.n6552 0.042
R20084 D.n6567 D.n6566 0.042
R20085 D.n6581 D.n6580 0.042
R20086 D.n6595 D.n6594 0.042
R20087 D.n6609 D.n6608 0.042
R20088 D.n6623 D.n6622 0.042
R20089 D.n6637 D.n6636 0.042
R20090 D.n6651 D.n6650 0.042
R20091 D.n6665 D.n6664 0.042
R20092 D.n6679 D.n6678 0.042
R20093 D.n6693 D.n6692 0.042
R20094 D.n6707 D.n6706 0.042
R20095 D.n6721 D.n6720 0.042
R20096 D.n6735 D.n6734 0.042
R20097 D.n6749 D.n6748 0.042
R20098 D.n6789 D.n6788 0.042
R20099 D.n6803 D.n6802 0.042
R20100 D.n6817 D.n6816 0.042
R20101 D.n6831 D.n6830 0.042
R20102 D.n6845 D.n6844 0.042
R20103 D.n6859 D.n6858 0.042
R20104 D.n6873 D.n6872 0.042
R20105 D.n6887 D.n6886 0.042
R20106 D.n6901 D.n6900 0.042
R20107 D.n6915 D.n6914 0.042
R20108 D.n6929 D.n6928 0.042
R20109 D.n6943 D.n6942 0.042
R20110 D.n6957 D.n6956 0.042
R20111 D.n6971 D.n6970 0.042
R20112 D.n6985 D.n6984 0.042
R20113 D.n7025 D.n7024 0.042
R20114 D.n7039 D.n7038 0.042
R20115 D.n7053 D.n7052 0.042
R20116 D.n7067 D.n7066 0.042
R20117 D.n7081 D.n7080 0.042
R20118 D.n7095 D.n7094 0.042
R20119 D.n7109 D.n7108 0.042
R20120 D.n7123 D.n7122 0.042
R20121 D.n7137 D.n7136 0.042
R20122 D.n7151 D.n7150 0.042
R20123 D.n7165 D.n7164 0.042
R20124 D.n7179 D.n7178 0.042
R20125 D.n7193 D.n7192 0.042
R20126 D.n7233 D.n7232 0.042
R20127 D.n7247 D.n7246 0.042
R20128 D.n7261 D.n7260 0.042
R20129 D.n7275 D.n7274 0.042
R20130 D.n7289 D.n7288 0.042
R20131 D.n7303 D.n7302 0.042
R20132 D.n7317 D.n7316 0.042
R20133 D.n7331 D.n7330 0.042
R20134 D.n7345 D.n7344 0.042
R20135 D.n7359 D.n7358 0.042
R20136 D.n7373 D.n7372 0.042
R20137 D.n7413 D.n7412 0.042
R20138 D.n7427 D.n7426 0.042
R20139 D.n7441 D.n7440 0.042
R20140 D.n7455 D.n7454 0.042
R20141 D.n7469 D.n7468 0.042
R20142 D.n7483 D.n7482 0.042
R20143 D.n7497 D.n7496 0.042
R20144 D.n7511 D.n7510 0.042
R20145 D.n7525 D.n7524 0.042
R20146 D.n7565 D.n7564 0.042
R20147 D.n7579 D.n7578 0.042
R20148 D.n7593 D.n7592 0.042
R20149 D.n7607 D.n7606 0.042
R20150 D.n7621 D.n7620 0.042
R20151 D.n7635 D.n7634 0.042
R20152 D.n7649 D.n7648 0.042
R20153 D.n7689 D.n7688 0.042
R20154 D.n7703 D.n7702 0.042
R20155 D.n7717 D.n7716 0.042
R20156 D.n7731 D.n7730 0.042
R20157 D.n7745 D.n7744 0.042
R20158 D.n7784 D.n7783 0.042
R20159 D.n7798 D.n7797 0.042
R20160 D.n7814 D.n7813 0.042
R20161 D.n13652 D.n13651 0.041
R20162 D.n12729 D.n12728 0.041
R20163 D.n11880 D.n11879 0.041
R20164 D.n11117 D.n11116 0.041
R20165 D.n10434 D.n10433 0.041
R20166 D.n9831 D.n9830 0.041
R20167 D.n9302 D.n9301 0.041
R20168 D.n8859 D.n8858 0.041
R20169 D.n8496 D.n8495 0.041
R20170 D.n8207 D.n8206 0.041
R20171 D.n8004 D.n8003 0.041
R20172 D.n13672 D.n13671 0.041
R20173 D.n12745 D.n12744 0.041
R20174 D.n11896 D.n11895 0.041
R20175 D.n11133 D.n11132 0.041
R20176 D.n10450 D.n10449 0.041
R20177 D.n9847 D.n9846 0.041
R20178 D.n9318 D.n9317 0.041
R20179 D.n8875 D.n8874 0.041
R20180 D.n8512 D.n8511 0.041
R20181 D.n8223 D.n8222 0.041
R20182 D.n8020 D.n8019 0.041
R20183 D.n7986 D.n7985 0.039
R20184 D.n7988 D.n7986 0.039
R20185 D.n7947 D.n7946 0.039
R20186 D.n13657 D.n13656 0.039
R20187 D.n13677 D.n13676 0.039
R20188 D.n13679 D.n13677 0.039
R20189 D.n14083 D.n14082 0.039
R20190 D.n13622 D.n13621 0.039
R20191 D.n13634 D.n13633 0.039
R20192 D.n13636 D.n13634 0.039
R20193 D.n13197 D.n13196 0.039
R20194 D.n13175 D.n13174 0.039
R20195 D.n12734 D.n12733 0.039
R20196 D.n12750 D.n12749 0.039
R20197 D.n12752 D.n12750 0.039
R20198 D.n12699 D.n12698 0.039
R20199 D.n12711 D.n12710 0.039
R20200 D.n12713 D.n12711 0.039
R20201 D.n12314 D.n12313 0.039
R20202 D.n12292 D.n12291 0.039
R20203 D.n11885 D.n11884 0.039
R20204 D.n11901 D.n11900 0.039
R20205 D.n11903 D.n11901 0.039
R20206 D.n12234 D.n12233 0.039
R20207 D.n11850 D.n11849 0.039
R20208 D.n11862 D.n11861 0.039
R20209 D.n11864 D.n11862 0.039
R20210 D.n11122 D.n11121 0.039
R20211 D.n11138 D.n11137 0.039
R20212 D.n11140 D.n11138 0.039
R20213 D.n11435 D.n11434 0.039
R20214 D.n11087 D.n11086 0.039
R20215 D.n11099 D.n11098 0.039
R20216 D.n11101 D.n11099 0.039
R20217 D.n10439 D.n10438 0.039
R20218 D.n10455 D.n10454 0.039
R20219 D.n10457 D.n10455 0.039
R20220 D.n10716 D.n10715 0.039
R20221 D.n10404 D.n10403 0.039
R20222 D.n10416 D.n10415 0.039
R20223 D.n10418 D.n10416 0.039
R20224 D.n10139 D.n10138 0.039
R20225 D.n10117 D.n10116 0.039
R20226 D.n9836 D.n9835 0.039
R20227 D.n9852 D.n9851 0.039
R20228 D.n9854 D.n9852 0.039
R20229 D.n9801 D.n9800 0.039
R20230 D.n9813 D.n9812 0.039
R20231 D.n9815 D.n9813 0.039
R20232 D.n9576 D.n9575 0.039
R20233 D.n9554 D.n9553 0.039
R20234 D.n9307 D.n9306 0.039
R20235 D.n9323 D.n9322 0.039
R20236 D.n9325 D.n9323 0.039
R20237 D.n9512 D.n9511 0.039
R20238 D.n9272 D.n9271 0.039
R20239 D.n9284 D.n9283 0.039
R20240 D.n9286 D.n9284 0.039
R20241 D.n8864 D.n8863 0.039
R20242 D.n8880 D.n8879 0.039
R20243 D.n8882 D.n8880 0.039
R20244 D.n9033 D.n9032 0.039
R20245 D.n8829 D.n8828 0.039
R20246 D.n8841 D.n8840 0.039
R20247 D.n8843 D.n8841 0.039
R20248 D.n8684 D.n8683 0.039
R20249 D.n8662 D.n8661 0.039
R20250 D.n8501 D.n8500 0.039
R20251 D.n8517 D.n8516 0.039
R20252 D.n8519 D.n8517 0.039
R20253 D.n8466 D.n8465 0.039
R20254 D.n8478 D.n8477 0.039
R20255 D.n8480 D.n8478 0.039
R20256 D.n8361 D.n8360 0.039
R20257 D.n8339 D.n8338 0.039
R20258 D.n8212 D.n8211 0.039
R20259 D.n8228 D.n8227 0.039
R20260 D.n8230 D.n8228 0.039
R20261 D.n8309 D.n8308 0.039
R20262 D.n8177 D.n8176 0.039
R20263 D.n8189 D.n8188 0.039
R20264 D.n8191 D.n8189 0.039
R20265 D.n8009 D.n8008 0.039
R20266 D.n8025 D.n8024 0.039
R20267 D.n8027 D.n8025 0.039
R20268 D.n8070 D.n8069 0.039
R20269 D.n7925 D.n7924 0.039
R20270 D.n7972 D.n7971 0.039
R20271 D.n7889 D.n7888 0.039
R20272 D.n7896 D.n7895 0.039
R20273 D.n7916 D.n7915 0.039
R20274 D.n47 D.n26 0.039
R20275 D D.n14144 0.038
R20276 D D.n7884 0.037
R20277 D.n7902 D.n7891 0.035
R20278 D.n7921 D.n7920 0.034
R20279 D.n533 D.n532 0.034
R20280 D.n1160 D.n1159 0.034
R20281 D.n1759 D.n1758 0.034
R20282 D.n2330 D.n2329 0.034
R20283 D.n2873 D.n2872 0.034
R20284 D.n3389 D.n3388 0.034
R20285 D.n3877 D.n3876 0.034
R20286 D.n4337 D.n4336 0.034
R20287 D.n4769 D.n4768 0.034
R20288 D.n5173 D.n5172 0.034
R20289 D.n5549 D.n5548 0.034
R20290 D.n5897 D.n5896 0.034
R20291 D.n6217 D.n6216 0.034
R20292 D.n6509 D.n6508 0.034
R20293 D.n6773 D.n6772 0.034
R20294 D.n7009 D.n7008 0.034
R20295 D.n7217 D.n7216 0.034
R20296 D.n7397 D.n7396 0.034
R20297 D.n7549 D.n7548 0.034
R20298 D.n7673 D.n7672 0.034
R20299 D.n7768 D.n7767 0.034
R20300 D.n7860 D.n7859 0.034
R20301 D.n13669 D.n13668 0.034
R20302 D.n7902 D.n7894 0.033
R20303 D.n7988 D.n7978 0.033
R20304 D.n13679 D.n13661 0.033
R20305 D.n13636 D.n13626 0.033
R20306 D.n12752 D.n12738 0.033
R20307 D.n12713 D.n12703 0.033
R20308 D.n11903 D.n11889 0.033
R20309 D.n11864 D.n11854 0.033
R20310 D.n11140 D.n11126 0.033
R20311 D.n11101 D.n11091 0.033
R20312 D.n10457 D.n10443 0.033
R20313 D.n10418 D.n10408 0.033
R20314 D.n9854 D.n9840 0.033
R20315 D.n9815 D.n9805 0.033
R20316 D.n9325 D.n9311 0.033
R20317 D.n9286 D.n9276 0.033
R20318 D.n8882 D.n8868 0.033
R20319 D.n8843 D.n8833 0.033
R20320 D.n8519 D.n8505 0.033
R20321 D.n8480 D.n8470 0.033
R20322 D.n8230 D.n8216 0.033
R20323 D.n8191 D.n8181 0.033
R20324 D.n8027 D.n8013 0.033
R20325 D.n7823 D.n7822 0.033
R20326 D.n14144 D.n14142 0.032
R20327 D.n511 D.n510 0.031
R20328 D.n7863 D.n7862 0.031
R20329 D.n7864 D.n7863 0.031
R20330 D.n7865 D.n7864 0.031
R20331 D.n7866 D.n7865 0.031
R20332 D.n7867 D.n7866 0.031
R20333 D.n7868 D.n7867 0.031
R20334 D.n7869 D.n7868 0.031
R20335 D.n7870 D.n7869 0.031
R20336 D.n7871 D.n7870 0.031
R20337 D.n7872 D.n7871 0.031
R20338 D.n7873 D.n7872 0.031
R20339 D.n7874 D.n7873 0.031
R20340 D.n7875 D.n7874 0.031
R20341 D.n7876 D.n7875 0.031
R20342 D.n7877 D.n7876 0.031
R20343 D.n7878 D.n7877 0.031
R20344 D.n7879 D.n7878 0.031
R20345 D.n7880 D.n7879 0.031
R20346 D.n7881 D.n7880 0.031
R20347 D.n7882 D.n7881 0.031
R20348 D.n7883 D.n7882 0.031
R20349 D.n7884 D.n7883 0.031
R20350 D.n7933 D.n7928 0.03
R20351 D.n14096 D.n14088 0.03
R20352 D.n14096 D.n14093 0.03
R20353 D.n13183 D.n13181 0.03
R20354 D.n13183 D.n13176 0.03
R20355 D.n12300 D.n12298 0.03
R20356 D.n12300 D.n12293 0.03
R20357 D.n12248 D.n12240 0.03
R20358 D.n12248 D.n12245 0.03
R20359 D.n11449 D.n11441 0.03
R20360 D.n11449 D.n11446 0.03
R20361 D.n10730 D.n10722 0.03
R20362 D.n10730 D.n10727 0.03
R20363 D.n10125 D.n10123 0.03
R20364 D.n10125 D.n10118 0.03
R20365 D.n9562 D.n9560 0.03
R20366 D.n9562 D.n9555 0.03
R20367 D.n9526 D.n9518 0.03
R20368 D.n9526 D.n9523 0.03
R20369 D.n9047 D.n9039 0.03
R20370 D.n9047 D.n9044 0.03
R20371 D.n8670 D.n8668 0.03
R20372 D.n8670 D.n8663 0.03
R20373 D.n8347 D.n8345 0.03
R20374 D.n8347 D.n8340 0.03
R20375 D.n8323 D.n8315 0.03
R20376 D.n8323 D.n8320 0.03
R20377 D.n8084 D.n8076 0.03
R20378 D.n8084 D.n8081 0.03
R20379 D.n7933 D.n7932 0.03
R20380 D.n7917 D.n7908 0.03
R20381 D.n7917 D.n7913 0.03
R20382 D.n13170 D.n13169 0.029
R20383 D.n12287 D.n12286 0.029
R20384 D.n11484 D.n11483 0.029
R20385 D.n10761 D.n10760 0.029
R20386 D.n10112 D.n10111 0.029
R20387 D.n9549 D.n9548 0.029
R20388 D.n9066 D.n9065 0.029
R20389 D.n8657 D.n8656 0.029
R20390 D.n8334 D.n8333 0.029
R20391 D.n8091 D.n8090 0.029
R20392 D.n14142 D.n13644 0.029
R20393 D.n13169 D.n12721 0.029
R20394 D.n12286 D.n11872 0.029
R20395 D.n11483 D.n11109 0.029
R20396 D.n10760 D.n10426 0.029
R20397 D.n10111 D.n9823 0.029
R20398 D.n9548 D.n9294 0.029
R20399 D.n9065 D.n8851 0.029
R20400 D.n8656 D.n8488 0.029
R20401 D.n8333 D.n8199 0.029
R20402 D.n8090 D.n7996 0.029
R20403 D.n25 D.n15 0.029
R20404 D.n23 D.n22 0.028
R20405 D.n41 D.n40 0.028
R20406 D.n23 D.n17 0.027
R20407 D.n13679 D.n13658 0.027
R20408 D.n13636 D.n13623 0.027
R20409 D.n12752 D.n12735 0.027
R20410 D.n12713 D.n12700 0.027
R20411 D.n11903 D.n11886 0.027
R20412 D.n11864 D.n11851 0.027
R20413 D.n11140 D.n11123 0.027
R20414 D.n11101 D.n11088 0.027
R20415 D.n10457 D.n10440 0.027
R20416 D.n10418 D.n10405 0.027
R20417 D.n9854 D.n9837 0.027
R20418 D.n9815 D.n9802 0.027
R20419 D.n9325 D.n9308 0.027
R20420 D.n9286 D.n9273 0.027
R20421 D.n8882 D.n8865 0.027
R20422 D.n8843 D.n8830 0.027
R20423 D.n8519 D.n8502 0.027
R20424 D.n8480 D.n8467 0.027
R20425 D.n8230 D.n8213 0.027
R20426 D.n8191 D.n8178 0.027
R20427 D.n8027 D.n8010 0.027
R20428 D.n7988 D.n7973 0.027
R20429 D.n7902 D.n7900 0.027
R20430 D.n47 D.n27 0.027
R20431 D.n3 D.n0 0.026
R20432 D.n41 D.n35 0.026
R20433 D.n1137 D.n1133 0.025
R20434 D.n1123 D.n1119 0.025
R20435 D.n1109 D.n1105 0.025
R20436 D.n1095 D.n1091 0.025
R20437 D.n1081 D.n1077 0.025
R20438 D.n1067 D.n1063 0.025
R20439 D.n1053 D.n1049 0.025
R20440 D.n1039 D.n1035 0.025
R20441 D.n1025 D.n1021 0.025
R20442 D.n1011 D.n1007 0.025
R20443 D.n997 D.n993 0.025
R20444 D.n983 D.n979 0.025
R20445 D.n969 D.n965 0.025
R20446 D.n955 D.n951 0.025
R20447 D.n941 D.n937 0.025
R20448 D.n927 D.n923 0.025
R20449 D.n913 D.n909 0.025
R20450 D.n899 D.n895 0.025
R20451 D.n885 D.n881 0.025
R20452 D.n871 D.n867 0.025
R20453 D.n857 D.n853 0.025
R20454 D.n843 D.n839 0.025
R20455 D.n829 D.n825 0.025
R20456 D.n815 D.n811 0.025
R20457 D.n801 D.n797 0.025
R20458 D.n787 D.n783 0.025
R20459 D.n773 D.n769 0.025
R20460 D.n759 D.n755 0.025
R20461 D.n745 D.n741 0.025
R20462 D.n731 D.n727 0.025
R20463 D.n717 D.n713 0.025
R20464 D.n703 D.n699 0.025
R20465 D.n689 D.n685 0.025
R20466 D.n675 D.n671 0.025
R20467 D.n661 D.n657 0.025
R20468 D.n647 D.n643 0.025
R20469 D.n633 D.n629 0.025
R20470 D.n619 D.n615 0.025
R20471 D.n605 D.n601 0.025
R20472 D.n591 D.n587 0.025
R20473 D.n577 D.n573 0.025
R20474 D.n563 D.n559 0.025
R20475 D.n549 D.n545 0.025
R20476 D.n535 D.n529 0.025
R20477 D.n1736 D.n1732 0.025
R20478 D.n1722 D.n1718 0.025
R20479 D.n1708 D.n1704 0.025
R20480 D.n1694 D.n1690 0.025
R20481 D.n1680 D.n1676 0.025
R20482 D.n1666 D.n1662 0.025
R20483 D.n1652 D.n1648 0.025
R20484 D.n1638 D.n1634 0.025
R20485 D.n1624 D.n1620 0.025
R20486 D.n1610 D.n1606 0.025
R20487 D.n1596 D.n1592 0.025
R20488 D.n1582 D.n1578 0.025
R20489 D.n1568 D.n1564 0.025
R20490 D.n1554 D.n1550 0.025
R20491 D.n1540 D.n1536 0.025
R20492 D.n1526 D.n1522 0.025
R20493 D.n1512 D.n1508 0.025
R20494 D.n1498 D.n1494 0.025
R20495 D.n1484 D.n1480 0.025
R20496 D.n1470 D.n1466 0.025
R20497 D.n1456 D.n1452 0.025
R20498 D.n1442 D.n1438 0.025
R20499 D.n1428 D.n1424 0.025
R20500 D.n1414 D.n1410 0.025
R20501 D.n1400 D.n1396 0.025
R20502 D.n1386 D.n1382 0.025
R20503 D.n1372 D.n1368 0.025
R20504 D.n1358 D.n1354 0.025
R20505 D.n1344 D.n1340 0.025
R20506 D.n1330 D.n1326 0.025
R20507 D.n1316 D.n1312 0.025
R20508 D.n1302 D.n1298 0.025
R20509 D.n1288 D.n1284 0.025
R20510 D.n1274 D.n1270 0.025
R20511 D.n1260 D.n1256 0.025
R20512 D.n1246 D.n1242 0.025
R20513 D.n1232 D.n1228 0.025
R20514 D.n1218 D.n1214 0.025
R20515 D.n1204 D.n1200 0.025
R20516 D.n1190 D.n1186 0.025
R20517 D.n1176 D.n1172 0.025
R20518 D.n1162 D.n1156 0.025
R20519 D.n2307 D.n2303 0.025
R20520 D.n2293 D.n2289 0.025
R20521 D.n2279 D.n2275 0.025
R20522 D.n2265 D.n2261 0.025
R20523 D.n2251 D.n2247 0.025
R20524 D.n2237 D.n2233 0.025
R20525 D.n2223 D.n2219 0.025
R20526 D.n2209 D.n2205 0.025
R20527 D.n2195 D.n2191 0.025
R20528 D.n2181 D.n2177 0.025
R20529 D.n2167 D.n2163 0.025
R20530 D.n2153 D.n2149 0.025
R20531 D.n2139 D.n2135 0.025
R20532 D.n2125 D.n2121 0.025
R20533 D.n2111 D.n2107 0.025
R20534 D.n2097 D.n2093 0.025
R20535 D.n2083 D.n2079 0.025
R20536 D.n2069 D.n2065 0.025
R20537 D.n2055 D.n2051 0.025
R20538 D.n2041 D.n2037 0.025
R20539 D.n2027 D.n2023 0.025
R20540 D.n2013 D.n2009 0.025
R20541 D.n1999 D.n1995 0.025
R20542 D.n1985 D.n1981 0.025
R20543 D.n1971 D.n1967 0.025
R20544 D.n1957 D.n1953 0.025
R20545 D.n1943 D.n1939 0.025
R20546 D.n1929 D.n1925 0.025
R20547 D.n1915 D.n1911 0.025
R20548 D.n1901 D.n1897 0.025
R20549 D.n1887 D.n1883 0.025
R20550 D.n1873 D.n1869 0.025
R20551 D.n1859 D.n1855 0.025
R20552 D.n1845 D.n1841 0.025
R20553 D.n1831 D.n1827 0.025
R20554 D.n1817 D.n1813 0.025
R20555 D.n1803 D.n1799 0.025
R20556 D.n1789 D.n1785 0.025
R20557 D.n1775 D.n1771 0.025
R20558 D.n1761 D.n1755 0.025
R20559 D.n2850 D.n2846 0.025
R20560 D.n2836 D.n2832 0.025
R20561 D.n2822 D.n2818 0.025
R20562 D.n2808 D.n2804 0.025
R20563 D.n2794 D.n2790 0.025
R20564 D.n2780 D.n2776 0.025
R20565 D.n2766 D.n2762 0.025
R20566 D.n2752 D.n2748 0.025
R20567 D.n2738 D.n2734 0.025
R20568 D.n2724 D.n2720 0.025
R20569 D.n2710 D.n2706 0.025
R20570 D.n2696 D.n2692 0.025
R20571 D.n2682 D.n2678 0.025
R20572 D.n2668 D.n2664 0.025
R20573 D.n2654 D.n2650 0.025
R20574 D.n2640 D.n2636 0.025
R20575 D.n2626 D.n2622 0.025
R20576 D.n2612 D.n2608 0.025
R20577 D.n2598 D.n2594 0.025
R20578 D.n2584 D.n2580 0.025
R20579 D.n2570 D.n2566 0.025
R20580 D.n2556 D.n2552 0.025
R20581 D.n2542 D.n2538 0.025
R20582 D.n2528 D.n2524 0.025
R20583 D.n2514 D.n2510 0.025
R20584 D.n2500 D.n2496 0.025
R20585 D.n2486 D.n2482 0.025
R20586 D.n2472 D.n2468 0.025
R20587 D.n2458 D.n2454 0.025
R20588 D.n2444 D.n2440 0.025
R20589 D.n2430 D.n2426 0.025
R20590 D.n2416 D.n2412 0.025
R20591 D.n2402 D.n2398 0.025
R20592 D.n2388 D.n2384 0.025
R20593 D.n2374 D.n2370 0.025
R20594 D.n2360 D.n2356 0.025
R20595 D.n2346 D.n2342 0.025
R20596 D.n2332 D.n2326 0.025
R20597 D.n3365 D.n3361 0.025
R20598 D.n3351 D.n3347 0.025
R20599 D.n3337 D.n3333 0.025
R20600 D.n3323 D.n3319 0.025
R20601 D.n3309 D.n3305 0.025
R20602 D.n3295 D.n3291 0.025
R20603 D.n3281 D.n3277 0.025
R20604 D.n3267 D.n3263 0.025
R20605 D.n3253 D.n3249 0.025
R20606 D.n3239 D.n3235 0.025
R20607 D.n3225 D.n3221 0.025
R20608 D.n3211 D.n3207 0.025
R20609 D.n3197 D.n3193 0.025
R20610 D.n3183 D.n3179 0.025
R20611 D.n3169 D.n3165 0.025
R20612 D.n3155 D.n3151 0.025
R20613 D.n3141 D.n3137 0.025
R20614 D.n3127 D.n3123 0.025
R20615 D.n3113 D.n3109 0.025
R20616 D.n3099 D.n3095 0.025
R20617 D.n3085 D.n3081 0.025
R20618 D.n3071 D.n3067 0.025
R20619 D.n3057 D.n3053 0.025
R20620 D.n3043 D.n3039 0.025
R20621 D.n3029 D.n3025 0.025
R20622 D.n3015 D.n3011 0.025
R20623 D.n3001 D.n2997 0.025
R20624 D.n2987 D.n2983 0.025
R20625 D.n2973 D.n2969 0.025
R20626 D.n2959 D.n2955 0.025
R20627 D.n2945 D.n2941 0.025
R20628 D.n2931 D.n2927 0.025
R20629 D.n2917 D.n2913 0.025
R20630 D.n2903 D.n2899 0.025
R20631 D.n2889 D.n2885 0.025
R20632 D.n2875 D.n2869 0.025
R20633 D.n3853 D.n3849 0.025
R20634 D.n3839 D.n3835 0.025
R20635 D.n3825 D.n3821 0.025
R20636 D.n3811 D.n3807 0.025
R20637 D.n3797 D.n3793 0.025
R20638 D.n3783 D.n3779 0.025
R20639 D.n3769 D.n3765 0.025
R20640 D.n3755 D.n3751 0.025
R20641 D.n3741 D.n3737 0.025
R20642 D.n3727 D.n3723 0.025
R20643 D.n3713 D.n3709 0.025
R20644 D.n3699 D.n3695 0.025
R20645 D.n3685 D.n3681 0.025
R20646 D.n3671 D.n3667 0.025
R20647 D.n3657 D.n3653 0.025
R20648 D.n3643 D.n3639 0.025
R20649 D.n3629 D.n3625 0.025
R20650 D.n3615 D.n3611 0.025
R20651 D.n3601 D.n3597 0.025
R20652 D.n3587 D.n3583 0.025
R20653 D.n3573 D.n3569 0.025
R20654 D.n3559 D.n3555 0.025
R20655 D.n3545 D.n3541 0.025
R20656 D.n3531 D.n3527 0.025
R20657 D.n3517 D.n3513 0.025
R20658 D.n3503 D.n3499 0.025
R20659 D.n3489 D.n3485 0.025
R20660 D.n3475 D.n3471 0.025
R20661 D.n3461 D.n3457 0.025
R20662 D.n3447 D.n3443 0.025
R20663 D.n3433 D.n3429 0.025
R20664 D.n3419 D.n3415 0.025
R20665 D.n3405 D.n3401 0.025
R20666 D.n3391 D.n3385 0.025
R20667 D.n4313 D.n4309 0.025
R20668 D.n4299 D.n4295 0.025
R20669 D.n4285 D.n4281 0.025
R20670 D.n4271 D.n4267 0.025
R20671 D.n4257 D.n4253 0.025
R20672 D.n4243 D.n4239 0.025
R20673 D.n4229 D.n4225 0.025
R20674 D.n4215 D.n4211 0.025
R20675 D.n4201 D.n4197 0.025
R20676 D.n4187 D.n4183 0.025
R20677 D.n4173 D.n4169 0.025
R20678 D.n4159 D.n4155 0.025
R20679 D.n4145 D.n4141 0.025
R20680 D.n4131 D.n4127 0.025
R20681 D.n4117 D.n4113 0.025
R20682 D.n4103 D.n4099 0.025
R20683 D.n4089 D.n4085 0.025
R20684 D.n4075 D.n4071 0.025
R20685 D.n4061 D.n4057 0.025
R20686 D.n4047 D.n4043 0.025
R20687 D.n4033 D.n4029 0.025
R20688 D.n4019 D.n4015 0.025
R20689 D.n4005 D.n4001 0.025
R20690 D.n3991 D.n3987 0.025
R20691 D.n3977 D.n3973 0.025
R20692 D.n3963 D.n3959 0.025
R20693 D.n3949 D.n3945 0.025
R20694 D.n3935 D.n3931 0.025
R20695 D.n3921 D.n3917 0.025
R20696 D.n3907 D.n3903 0.025
R20697 D.n3893 D.n3889 0.025
R20698 D.n3879 D.n3873 0.025
R20699 D.n4745 D.n4741 0.025
R20700 D.n4731 D.n4727 0.025
R20701 D.n4717 D.n4713 0.025
R20702 D.n4703 D.n4699 0.025
R20703 D.n4689 D.n4685 0.025
R20704 D.n4675 D.n4671 0.025
R20705 D.n4661 D.n4657 0.025
R20706 D.n4647 D.n4643 0.025
R20707 D.n4633 D.n4629 0.025
R20708 D.n4619 D.n4615 0.025
R20709 D.n4605 D.n4601 0.025
R20710 D.n4591 D.n4587 0.025
R20711 D.n4577 D.n4573 0.025
R20712 D.n4563 D.n4559 0.025
R20713 D.n4549 D.n4545 0.025
R20714 D.n4535 D.n4531 0.025
R20715 D.n4521 D.n4517 0.025
R20716 D.n4507 D.n4503 0.025
R20717 D.n4493 D.n4489 0.025
R20718 D.n4479 D.n4475 0.025
R20719 D.n4465 D.n4461 0.025
R20720 D.n4451 D.n4447 0.025
R20721 D.n4437 D.n4433 0.025
R20722 D.n4423 D.n4419 0.025
R20723 D.n4409 D.n4405 0.025
R20724 D.n4395 D.n4391 0.025
R20725 D.n4381 D.n4377 0.025
R20726 D.n4367 D.n4363 0.025
R20727 D.n4353 D.n4349 0.025
R20728 D.n4339 D.n4333 0.025
R20729 D.n5149 D.n5145 0.025
R20730 D.n5135 D.n5131 0.025
R20731 D.n5121 D.n5117 0.025
R20732 D.n5107 D.n5103 0.025
R20733 D.n5093 D.n5089 0.025
R20734 D.n5079 D.n5075 0.025
R20735 D.n5065 D.n5061 0.025
R20736 D.n5051 D.n5047 0.025
R20737 D.n5037 D.n5033 0.025
R20738 D.n5023 D.n5019 0.025
R20739 D.n5009 D.n5005 0.025
R20740 D.n4995 D.n4991 0.025
R20741 D.n4981 D.n4977 0.025
R20742 D.n4967 D.n4963 0.025
R20743 D.n4953 D.n4949 0.025
R20744 D.n4939 D.n4935 0.025
R20745 D.n4925 D.n4921 0.025
R20746 D.n4911 D.n4907 0.025
R20747 D.n4897 D.n4893 0.025
R20748 D.n4883 D.n4879 0.025
R20749 D.n4869 D.n4865 0.025
R20750 D.n4855 D.n4851 0.025
R20751 D.n4841 D.n4837 0.025
R20752 D.n4827 D.n4823 0.025
R20753 D.n4813 D.n4809 0.025
R20754 D.n4799 D.n4795 0.025
R20755 D.n4785 D.n4781 0.025
R20756 D.n4771 D.n4765 0.025
R20757 D.n5525 D.n5521 0.025
R20758 D.n5511 D.n5507 0.025
R20759 D.n5497 D.n5493 0.025
R20760 D.n5483 D.n5479 0.025
R20761 D.n5469 D.n5465 0.025
R20762 D.n5455 D.n5451 0.025
R20763 D.n5441 D.n5437 0.025
R20764 D.n5427 D.n5423 0.025
R20765 D.n5413 D.n5409 0.025
R20766 D.n5399 D.n5395 0.025
R20767 D.n5385 D.n5381 0.025
R20768 D.n5371 D.n5367 0.025
R20769 D.n5357 D.n5353 0.025
R20770 D.n5343 D.n5339 0.025
R20771 D.n5329 D.n5325 0.025
R20772 D.n5315 D.n5311 0.025
R20773 D.n5301 D.n5297 0.025
R20774 D.n5287 D.n5283 0.025
R20775 D.n5273 D.n5269 0.025
R20776 D.n5259 D.n5255 0.025
R20777 D.n5245 D.n5241 0.025
R20778 D.n5231 D.n5227 0.025
R20779 D.n5217 D.n5213 0.025
R20780 D.n5203 D.n5199 0.025
R20781 D.n5189 D.n5185 0.025
R20782 D.n5175 D.n5169 0.025
R20783 D.n5873 D.n5869 0.025
R20784 D.n5859 D.n5855 0.025
R20785 D.n5845 D.n5841 0.025
R20786 D.n5831 D.n5827 0.025
R20787 D.n5817 D.n5813 0.025
R20788 D.n5803 D.n5799 0.025
R20789 D.n5789 D.n5785 0.025
R20790 D.n5775 D.n5771 0.025
R20791 D.n5761 D.n5757 0.025
R20792 D.n5747 D.n5743 0.025
R20793 D.n5733 D.n5729 0.025
R20794 D.n5719 D.n5715 0.025
R20795 D.n5705 D.n5701 0.025
R20796 D.n5691 D.n5687 0.025
R20797 D.n5677 D.n5673 0.025
R20798 D.n5663 D.n5659 0.025
R20799 D.n5649 D.n5645 0.025
R20800 D.n5635 D.n5631 0.025
R20801 D.n5621 D.n5617 0.025
R20802 D.n5607 D.n5603 0.025
R20803 D.n5593 D.n5589 0.025
R20804 D.n5579 D.n5575 0.025
R20805 D.n5565 D.n5561 0.025
R20806 D.n5551 D.n5545 0.025
R20807 D.n6193 D.n6189 0.025
R20808 D.n6179 D.n6175 0.025
R20809 D.n6165 D.n6161 0.025
R20810 D.n6151 D.n6147 0.025
R20811 D.n6137 D.n6133 0.025
R20812 D.n6123 D.n6119 0.025
R20813 D.n6109 D.n6105 0.025
R20814 D.n6095 D.n6091 0.025
R20815 D.n6081 D.n6077 0.025
R20816 D.n6067 D.n6063 0.025
R20817 D.n6053 D.n6049 0.025
R20818 D.n6039 D.n6035 0.025
R20819 D.n6025 D.n6021 0.025
R20820 D.n6011 D.n6007 0.025
R20821 D.n5997 D.n5993 0.025
R20822 D.n5983 D.n5979 0.025
R20823 D.n5969 D.n5965 0.025
R20824 D.n5955 D.n5951 0.025
R20825 D.n5941 D.n5937 0.025
R20826 D.n5927 D.n5923 0.025
R20827 D.n5913 D.n5909 0.025
R20828 D.n5899 D.n5893 0.025
R20829 D.n6485 D.n6481 0.025
R20830 D.n6471 D.n6467 0.025
R20831 D.n6457 D.n6453 0.025
R20832 D.n6443 D.n6439 0.025
R20833 D.n6429 D.n6425 0.025
R20834 D.n6415 D.n6411 0.025
R20835 D.n6401 D.n6397 0.025
R20836 D.n6387 D.n6383 0.025
R20837 D.n6373 D.n6369 0.025
R20838 D.n6359 D.n6355 0.025
R20839 D.n6345 D.n6341 0.025
R20840 D.n6331 D.n6327 0.025
R20841 D.n6317 D.n6313 0.025
R20842 D.n6303 D.n6299 0.025
R20843 D.n6289 D.n6285 0.025
R20844 D.n6275 D.n6271 0.025
R20845 D.n6261 D.n6257 0.025
R20846 D.n6247 D.n6243 0.025
R20847 D.n6233 D.n6229 0.025
R20848 D.n6219 D.n6213 0.025
R20849 D.n6749 D.n6745 0.025
R20850 D.n6735 D.n6731 0.025
R20851 D.n6721 D.n6717 0.025
R20852 D.n6707 D.n6703 0.025
R20853 D.n6693 D.n6689 0.025
R20854 D.n6679 D.n6675 0.025
R20855 D.n6665 D.n6661 0.025
R20856 D.n6651 D.n6647 0.025
R20857 D.n6637 D.n6633 0.025
R20858 D.n6623 D.n6619 0.025
R20859 D.n6609 D.n6605 0.025
R20860 D.n6595 D.n6591 0.025
R20861 D.n6581 D.n6577 0.025
R20862 D.n6567 D.n6563 0.025
R20863 D.n6553 D.n6549 0.025
R20864 D.n6539 D.n6535 0.025
R20865 D.n6525 D.n6521 0.025
R20866 D.n6511 D.n6505 0.025
R20867 D.n6985 D.n6981 0.025
R20868 D.n6971 D.n6967 0.025
R20869 D.n6957 D.n6953 0.025
R20870 D.n6943 D.n6939 0.025
R20871 D.n6929 D.n6925 0.025
R20872 D.n6915 D.n6911 0.025
R20873 D.n6901 D.n6897 0.025
R20874 D.n6887 D.n6883 0.025
R20875 D.n6873 D.n6869 0.025
R20876 D.n6859 D.n6855 0.025
R20877 D.n6845 D.n6841 0.025
R20878 D.n6831 D.n6827 0.025
R20879 D.n6817 D.n6813 0.025
R20880 D.n6803 D.n6799 0.025
R20881 D.n6789 D.n6785 0.025
R20882 D.n6775 D.n6769 0.025
R20883 D.n7193 D.n7189 0.025
R20884 D.n7179 D.n7175 0.025
R20885 D.n7165 D.n7161 0.025
R20886 D.n7151 D.n7147 0.025
R20887 D.n7137 D.n7133 0.025
R20888 D.n7123 D.n7119 0.025
R20889 D.n7109 D.n7105 0.025
R20890 D.n7095 D.n7091 0.025
R20891 D.n7081 D.n7077 0.025
R20892 D.n7067 D.n7063 0.025
R20893 D.n7053 D.n7049 0.025
R20894 D.n7039 D.n7035 0.025
R20895 D.n7025 D.n7021 0.025
R20896 D.n7011 D.n7005 0.025
R20897 D.n7373 D.n7369 0.025
R20898 D.n7359 D.n7355 0.025
R20899 D.n7345 D.n7341 0.025
R20900 D.n7331 D.n7327 0.025
R20901 D.n7317 D.n7313 0.025
R20902 D.n7303 D.n7299 0.025
R20903 D.n7289 D.n7285 0.025
R20904 D.n7275 D.n7271 0.025
R20905 D.n7261 D.n7257 0.025
R20906 D.n7247 D.n7243 0.025
R20907 D.n7233 D.n7229 0.025
R20908 D.n7219 D.n7213 0.025
R20909 D.n7525 D.n7521 0.025
R20910 D.n7511 D.n7507 0.025
R20911 D.n7497 D.n7493 0.025
R20912 D.n7483 D.n7479 0.025
R20913 D.n7469 D.n7465 0.025
R20914 D.n7455 D.n7451 0.025
R20915 D.n7441 D.n7437 0.025
R20916 D.n7427 D.n7423 0.025
R20917 D.n7413 D.n7409 0.025
R20918 D.n7399 D.n7393 0.025
R20919 D.n7649 D.n7645 0.025
R20920 D.n7635 D.n7631 0.025
R20921 D.n7621 D.n7617 0.025
R20922 D.n7607 D.n7603 0.025
R20923 D.n7593 D.n7589 0.025
R20924 D.n7579 D.n7575 0.025
R20925 D.n7565 D.n7561 0.025
R20926 D.n7551 D.n7545 0.025
R20927 D.n7745 D.n7741 0.025
R20928 D.n7731 D.n7727 0.025
R20929 D.n7717 D.n7713 0.025
R20930 D.n7703 D.n7699 0.025
R20931 D.n7689 D.n7685 0.025
R20932 D.n7675 D.n7669 0.025
R20933 D.n7814 D.n7810 0.025
R20934 D.n7798 D.n7794 0.025
R20935 D.n7784 D.n7780 0.025
R20936 D.n7770 D.n7764 0.025
R20937 D.n505 D.n504 0.024
R20938 D.n26 D.n25 0.023
R20939 D.n7983 D.n7980 0.023
R20940 D.n7985 D.n7984 0.023
R20941 D.n13654 D.n13647 0.023
R20942 D.n13656 D.n13655 0.023
R20943 D.n13674 D.n13663 0.023
R20944 D.n13676 D.n13675 0.023
R20945 D.n13619 D.n13616 0.023
R20946 D.n13621 D.n13620 0.023
R20947 D.n13631 D.n13628 0.023
R20948 D.n13633 D.n13632 0.023
R20949 D.n12731 D.n12724 0.023
R20950 D.n12733 D.n12732 0.023
R20951 D.n12747 D.n12740 0.023
R20952 D.n12749 D.n12748 0.023
R20953 D.n12696 D.n12693 0.023
R20954 D.n12698 D.n12697 0.023
R20955 D.n12708 D.n12705 0.023
R20956 D.n12710 D.n12709 0.023
R20957 D.n11882 D.n11875 0.023
R20958 D.n11884 D.n11883 0.023
R20959 D.n11898 D.n11891 0.023
R20960 D.n11900 D.n11899 0.023
R20961 D.n11847 D.n11844 0.023
R20962 D.n11849 D.n11848 0.023
R20963 D.n11859 D.n11856 0.023
R20964 D.n11861 D.n11860 0.023
R20965 D.n11119 D.n11112 0.023
R20966 D.n11121 D.n11120 0.023
R20967 D.n11135 D.n11128 0.023
R20968 D.n11137 D.n11136 0.023
R20969 D.n11084 D.n11081 0.023
R20970 D.n11086 D.n11085 0.023
R20971 D.n11096 D.n11093 0.023
R20972 D.n11098 D.n11097 0.023
R20973 D.n10436 D.n10429 0.023
R20974 D.n10438 D.n10437 0.023
R20975 D.n10452 D.n10445 0.023
R20976 D.n10454 D.n10453 0.023
R20977 D.n10401 D.n10398 0.023
R20978 D.n10403 D.n10402 0.023
R20979 D.n10413 D.n10410 0.023
R20980 D.n10415 D.n10414 0.023
R20981 D.n9833 D.n9826 0.023
R20982 D.n9835 D.n9834 0.023
R20983 D.n9849 D.n9842 0.023
R20984 D.n9851 D.n9850 0.023
R20985 D.n9798 D.n9795 0.023
R20986 D.n9800 D.n9799 0.023
R20987 D.n9810 D.n9807 0.023
R20988 D.n9812 D.n9811 0.023
R20989 D.n9304 D.n9297 0.023
R20990 D.n9306 D.n9305 0.023
R20991 D.n9320 D.n9313 0.023
R20992 D.n9322 D.n9321 0.023
R20993 D.n9269 D.n9266 0.023
R20994 D.n9271 D.n9270 0.023
R20995 D.n9281 D.n9278 0.023
R20996 D.n9283 D.n9282 0.023
R20997 D.n8861 D.n8854 0.023
R20998 D.n8863 D.n8862 0.023
R20999 D.n8877 D.n8870 0.023
R21000 D.n8879 D.n8878 0.023
R21001 D.n8826 D.n8823 0.023
R21002 D.n8828 D.n8827 0.023
R21003 D.n8838 D.n8835 0.023
R21004 D.n8840 D.n8839 0.023
R21005 D.n8498 D.n8491 0.023
R21006 D.n8500 D.n8499 0.023
R21007 D.n8514 D.n8507 0.023
R21008 D.n8516 D.n8515 0.023
R21009 D.n8463 D.n8460 0.023
R21010 D.n8465 D.n8464 0.023
R21011 D.n8475 D.n8472 0.023
R21012 D.n8477 D.n8476 0.023
R21013 D.n8209 D.n8202 0.023
R21014 D.n8211 D.n8210 0.023
R21015 D.n8225 D.n8218 0.023
R21016 D.n8227 D.n8226 0.023
R21017 D.n8174 D.n8171 0.023
R21018 D.n8176 D.n8175 0.023
R21019 D.n8186 D.n8183 0.023
R21020 D.n8188 D.n8187 0.023
R21021 D.n8006 D.n7999 0.023
R21022 D.n8008 D.n8007 0.023
R21023 D.n8022 D.n8015 0.023
R21024 D.n8024 D.n8023 0.023
R21025 D.n7971 D.n7970 0.023
R21026 D.n7969 D.n7966 0.023
R21027 D.n44 D.n43 0.023
R21028 D.n1141 D.n1140 0.023
R21029 D.n549 D.n547 0.023
R21030 D.n563 D.n561 0.023
R21031 D.n577 D.n575 0.023
R21032 D.n591 D.n589 0.023
R21033 D.n605 D.n603 0.023
R21034 D.n619 D.n617 0.023
R21035 D.n633 D.n631 0.023
R21036 D.n647 D.n645 0.023
R21037 D.n661 D.n659 0.023
R21038 D.n675 D.n673 0.023
R21039 D.n689 D.n687 0.023
R21040 D.n703 D.n701 0.023
R21041 D.n717 D.n715 0.023
R21042 D.n731 D.n729 0.023
R21043 D.n745 D.n743 0.023
R21044 D.n759 D.n757 0.023
R21045 D.n773 D.n771 0.023
R21046 D.n787 D.n785 0.023
R21047 D.n801 D.n799 0.023
R21048 D.n815 D.n813 0.023
R21049 D.n829 D.n827 0.023
R21050 D.n843 D.n841 0.023
R21051 D.n857 D.n855 0.023
R21052 D.n871 D.n869 0.023
R21053 D.n885 D.n883 0.023
R21054 D.n899 D.n897 0.023
R21055 D.n913 D.n911 0.023
R21056 D.n927 D.n925 0.023
R21057 D.n941 D.n939 0.023
R21058 D.n955 D.n953 0.023
R21059 D.n969 D.n967 0.023
R21060 D.n983 D.n981 0.023
R21061 D.n997 D.n995 0.023
R21062 D.n1011 D.n1009 0.023
R21063 D.n1025 D.n1023 0.023
R21064 D.n1039 D.n1037 0.023
R21065 D.n1053 D.n1051 0.023
R21066 D.n1067 D.n1065 0.023
R21067 D.n1081 D.n1079 0.023
R21068 D.n1095 D.n1093 0.023
R21069 D.n1109 D.n1107 0.023
R21070 D.n1123 D.n1121 0.023
R21071 D.n1137 D.n1135 0.023
R21072 D.n1740 D.n1739 0.023
R21073 D.n1176 D.n1174 0.023
R21074 D.n1190 D.n1188 0.023
R21075 D.n1204 D.n1202 0.023
R21076 D.n1218 D.n1216 0.023
R21077 D.n1232 D.n1230 0.023
R21078 D.n1246 D.n1244 0.023
R21079 D.n1260 D.n1258 0.023
R21080 D.n1274 D.n1272 0.023
R21081 D.n1288 D.n1286 0.023
R21082 D.n1302 D.n1300 0.023
R21083 D.n1316 D.n1314 0.023
R21084 D.n1330 D.n1328 0.023
R21085 D.n1344 D.n1342 0.023
R21086 D.n1358 D.n1356 0.023
R21087 D.n1372 D.n1370 0.023
R21088 D.n1386 D.n1384 0.023
R21089 D.n1400 D.n1398 0.023
R21090 D.n1414 D.n1412 0.023
R21091 D.n1428 D.n1426 0.023
R21092 D.n1442 D.n1440 0.023
R21093 D.n1456 D.n1454 0.023
R21094 D.n1470 D.n1468 0.023
R21095 D.n1484 D.n1482 0.023
R21096 D.n1498 D.n1496 0.023
R21097 D.n1512 D.n1510 0.023
R21098 D.n1526 D.n1524 0.023
R21099 D.n1540 D.n1538 0.023
R21100 D.n1554 D.n1552 0.023
R21101 D.n1568 D.n1566 0.023
R21102 D.n1582 D.n1580 0.023
R21103 D.n1596 D.n1594 0.023
R21104 D.n1610 D.n1608 0.023
R21105 D.n1624 D.n1622 0.023
R21106 D.n1638 D.n1636 0.023
R21107 D.n1652 D.n1650 0.023
R21108 D.n1666 D.n1664 0.023
R21109 D.n1680 D.n1678 0.023
R21110 D.n1694 D.n1692 0.023
R21111 D.n1708 D.n1706 0.023
R21112 D.n1722 D.n1720 0.023
R21113 D.n1736 D.n1734 0.023
R21114 D.n2311 D.n2310 0.023
R21115 D.n1775 D.n1773 0.023
R21116 D.n1789 D.n1787 0.023
R21117 D.n1803 D.n1801 0.023
R21118 D.n1817 D.n1815 0.023
R21119 D.n1831 D.n1829 0.023
R21120 D.n1845 D.n1843 0.023
R21121 D.n1859 D.n1857 0.023
R21122 D.n1873 D.n1871 0.023
R21123 D.n1887 D.n1885 0.023
R21124 D.n1901 D.n1899 0.023
R21125 D.n1915 D.n1913 0.023
R21126 D.n1929 D.n1927 0.023
R21127 D.n1943 D.n1941 0.023
R21128 D.n1957 D.n1955 0.023
R21129 D.n1971 D.n1969 0.023
R21130 D.n1985 D.n1983 0.023
R21131 D.n1999 D.n1997 0.023
R21132 D.n2013 D.n2011 0.023
R21133 D.n2027 D.n2025 0.023
R21134 D.n2041 D.n2039 0.023
R21135 D.n2055 D.n2053 0.023
R21136 D.n2069 D.n2067 0.023
R21137 D.n2083 D.n2081 0.023
R21138 D.n2097 D.n2095 0.023
R21139 D.n2111 D.n2109 0.023
R21140 D.n2125 D.n2123 0.023
R21141 D.n2139 D.n2137 0.023
R21142 D.n2153 D.n2151 0.023
R21143 D.n2167 D.n2165 0.023
R21144 D.n2181 D.n2179 0.023
R21145 D.n2195 D.n2193 0.023
R21146 D.n2209 D.n2207 0.023
R21147 D.n2223 D.n2221 0.023
R21148 D.n2237 D.n2235 0.023
R21149 D.n2251 D.n2249 0.023
R21150 D.n2265 D.n2263 0.023
R21151 D.n2279 D.n2277 0.023
R21152 D.n2293 D.n2291 0.023
R21153 D.n2307 D.n2305 0.023
R21154 D.n2854 D.n2853 0.023
R21155 D.n2346 D.n2344 0.023
R21156 D.n2360 D.n2358 0.023
R21157 D.n2374 D.n2372 0.023
R21158 D.n2388 D.n2386 0.023
R21159 D.n2402 D.n2400 0.023
R21160 D.n2416 D.n2414 0.023
R21161 D.n2430 D.n2428 0.023
R21162 D.n2444 D.n2442 0.023
R21163 D.n2458 D.n2456 0.023
R21164 D.n2472 D.n2470 0.023
R21165 D.n2486 D.n2484 0.023
R21166 D.n2500 D.n2498 0.023
R21167 D.n2514 D.n2512 0.023
R21168 D.n2528 D.n2526 0.023
R21169 D.n2542 D.n2540 0.023
R21170 D.n2556 D.n2554 0.023
R21171 D.n2570 D.n2568 0.023
R21172 D.n2584 D.n2582 0.023
R21173 D.n2598 D.n2596 0.023
R21174 D.n2612 D.n2610 0.023
R21175 D.n2626 D.n2624 0.023
R21176 D.n2640 D.n2638 0.023
R21177 D.n2654 D.n2652 0.023
R21178 D.n2668 D.n2666 0.023
R21179 D.n2682 D.n2680 0.023
R21180 D.n2696 D.n2694 0.023
R21181 D.n2710 D.n2708 0.023
R21182 D.n2724 D.n2722 0.023
R21183 D.n2738 D.n2736 0.023
R21184 D.n2752 D.n2750 0.023
R21185 D.n2766 D.n2764 0.023
R21186 D.n2780 D.n2778 0.023
R21187 D.n2794 D.n2792 0.023
R21188 D.n2808 D.n2806 0.023
R21189 D.n2822 D.n2820 0.023
R21190 D.n2836 D.n2834 0.023
R21191 D.n2850 D.n2848 0.023
R21192 D.n3369 D.n3368 0.023
R21193 D.n2889 D.n2887 0.023
R21194 D.n2903 D.n2901 0.023
R21195 D.n2917 D.n2915 0.023
R21196 D.n2931 D.n2929 0.023
R21197 D.n2945 D.n2943 0.023
R21198 D.n2959 D.n2957 0.023
R21199 D.n2973 D.n2971 0.023
R21200 D.n2987 D.n2985 0.023
R21201 D.n3001 D.n2999 0.023
R21202 D.n3015 D.n3013 0.023
R21203 D.n3029 D.n3027 0.023
R21204 D.n3043 D.n3041 0.023
R21205 D.n3057 D.n3055 0.023
R21206 D.n3071 D.n3069 0.023
R21207 D.n3085 D.n3083 0.023
R21208 D.n3099 D.n3097 0.023
R21209 D.n3113 D.n3111 0.023
R21210 D.n3127 D.n3125 0.023
R21211 D.n3141 D.n3139 0.023
R21212 D.n3155 D.n3153 0.023
R21213 D.n3169 D.n3167 0.023
R21214 D.n3183 D.n3181 0.023
R21215 D.n3197 D.n3195 0.023
R21216 D.n3211 D.n3209 0.023
R21217 D.n3225 D.n3223 0.023
R21218 D.n3239 D.n3237 0.023
R21219 D.n3253 D.n3251 0.023
R21220 D.n3267 D.n3265 0.023
R21221 D.n3281 D.n3279 0.023
R21222 D.n3295 D.n3293 0.023
R21223 D.n3309 D.n3307 0.023
R21224 D.n3323 D.n3321 0.023
R21225 D.n3337 D.n3335 0.023
R21226 D.n3351 D.n3349 0.023
R21227 D.n3365 D.n3363 0.023
R21228 D.n3857 D.n3856 0.023
R21229 D.n3405 D.n3403 0.023
R21230 D.n3419 D.n3417 0.023
R21231 D.n3433 D.n3431 0.023
R21232 D.n3447 D.n3445 0.023
R21233 D.n3461 D.n3459 0.023
R21234 D.n3475 D.n3473 0.023
R21235 D.n3489 D.n3487 0.023
R21236 D.n3503 D.n3501 0.023
R21237 D.n3517 D.n3515 0.023
R21238 D.n3531 D.n3529 0.023
R21239 D.n3545 D.n3543 0.023
R21240 D.n3559 D.n3557 0.023
R21241 D.n3573 D.n3571 0.023
R21242 D.n3587 D.n3585 0.023
R21243 D.n3601 D.n3599 0.023
R21244 D.n3615 D.n3613 0.023
R21245 D.n3629 D.n3627 0.023
R21246 D.n3643 D.n3641 0.023
R21247 D.n3657 D.n3655 0.023
R21248 D.n3671 D.n3669 0.023
R21249 D.n3685 D.n3683 0.023
R21250 D.n3699 D.n3697 0.023
R21251 D.n3713 D.n3711 0.023
R21252 D.n3727 D.n3725 0.023
R21253 D.n3741 D.n3739 0.023
R21254 D.n3755 D.n3753 0.023
R21255 D.n3769 D.n3767 0.023
R21256 D.n3783 D.n3781 0.023
R21257 D.n3797 D.n3795 0.023
R21258 D.n3811 D.n3809 0.023
R21259 D.n3825 D.n3823 0.023
R21260 D.n3839 D.n3837 0.023
R21261 D.n3853 D.n3851 0.023
R21262 D.n4317 D.n4316 0.023
R21263 D.n3893 D.n3891 0.023
R21264 D.n3907 D.n3905 0.023
R21265 D.n3921 D.n3919 0.023
R21266 D.n3935 D.n3933 0.023
R21267 D.n3949 D.n3947 0.023
R21268 D.n3963 D.n3961 0.023
R21269 D.n3977 D.n3975 0.023
R21270 D.n3991 D.n3989 0.023
R21271 D.n4005 D.n4003 0.023
R21272 D.n4019 D.n4017 0.023
R21273 D.n4033 D.n4031 0.023
R21274 D.n4047 D.n4045 0.023
R21275 D.n4061 D.n4059 0.023
R21276 D.n4075 D.n4073 0.023
R21277 D.n4089 D.n4087 0.023
R21278 D.n4103 D.n4101 0.023
R21279 D.n4117 D.n4115 0.023
R21280 D.n4131 D.n4129 0.023
R21281 D.n4145 D.n4143 0.023
R21282 D.n4159 D.n4157 0.023
R21283 D.n4173 D.n4171 0.023
R21284 D.n4187 D.n4185 0.023
R21285 D.n4201 D.n4199 0.023
R21286 D.n4215 D.n4213 0.023
R21287 D.n4229 D.n4227 0.023
R21288 D.n4243 D.n4241 0.023
R21289 D.n4257 D.n4255 0.023
R21290 D.n4271 D.n4269 0.023
R21291 D.n4285 D.n4283 0.023
R21292 D.n4299 D.n4297 0.023
R21293 D.n4313 D.n4311 0.023
R21294 D.n4749 D.n4748 0.023
R21295 D.n4353 D.n4351 0.023
R21296 D.n4367 D.n4365 0.023
R21297 D.n4381 D.n4379 0.023
R21298 D.n4395 D.n4393 0.023
R21299 D.n4409 D.n4407 0.023
R21300 D.n4423 D.n4421 0.023
R21301 D.n4437 D.n4435 0.023
R21302 D.n4451 D.n4449 0.023
R21303 D.n4465 D.n4463 0.023
R21304 D.n4479 D.n4477 0.023
R21305 D.n4493 D.n4491 0.023
R21306 D.n4507 D.n4505 0.023
R21307 D.n4521 D.n4519 0.023
R21308 D.n4535 D.n4533 0.023
R21309 D.n4549 D.n4547 0.023
R21310 D.n4563 D.n4561 0.023
R21311 D.n4577 D.n4575 0.023
R21312 D.n4591 D.n4589 0.023
R21313 D.n4605 D.n4603 0.023
R21314 D.n4619 D.n4617 0.023
R21315 D.n4633 D.n4631 0.023
R21316 D.n4647 D.n4645 0.023
R21317 D.n4661 D.n4659 0.023
R21318 D.n4675 D.n4673 0.023
R21319 D.n4689 D.n4687 0.023
R21320 D.n4703 D.n4701 0.023
R21321 D.n4717 D.n4715 0.023
R21322 D.n4731 D.n4729 0.023
R21323 D.n4745 D.n4743 0.023
R21324 D.n5153 D.n5152 0.023
R21325 D.n4785 D.n4783 0.023
R21326 D.n4799 D.n4797 0.023
R21327 D.n4813 D.n4811 0.023
R21328 D.n4827 D.n4825 0.023
R21329 D.n4841 D.n4839 0.023
R21330 D.n4855 D.n4853 0.023
R21331 D.n4869 D.n4867 0.023
R21332 D.n4883 D.n4881 0.023
R21333 D.n4897 D.n4895 0.023
R21334 D.n4911 D.n4909 0.023
R21335 D.n4925 D.n4923 0.023
R21336 D.n4939 D.n4937 0.023
R21337 D.n4953 D.n4951 0.023
R21338 D.n4967 D.n4965 0.023
R21339 D.n4981 D.n4979 0.023
R21340 D.n4995 D.n4993 0.023
R21341 D.n5009 D.n5007 0.023
R21342 D.n5023 D.n5021 0.023
R21343 D.n5037 D.n5035 0.023
R21344 D.n5051 D.n5049 0.023
R21345 D.n5065 D.n5063 0.023
R21346 D.n5079 D.n5077 0.023
R21347 D.n5093 D.n5091 0.023
R21348 D.n5107 D.n5105 0.023
R21349 D.n5121 D.n5119 0.023
R21350 D.n5135 D.n5133 0.023
R21351 D.n5149 D.n5147 0.023
R21352 D.n5529 D.n5528 0.023
R21353 D.n5189 D.n5187 0.023
R21354 D.n5203 D.n5201 0.023
R21355 D.n5217 D.n5215 0.023
R21356 D.n5231 D.n5229 0.023
R21357 D.n5245 D.n5243 0.023
R21358 D.n5259 D.n5257 0.023
R21359 D.n5273 D.n5271 0.023
R21360 D.n5287 D.n5285 0.023
R21361 D.n5301 D.n5299 0.023
R21362 D.n5315 D.n5313 0.023
R21363 D.n5329 D.n5327 0.023
R21364 D.n5343 D.n5341 0.023
R21365 D.n5357 D.n5355 0.023
R21366 D.n5371 D.n5369 0.023
R21367 D.n5385 D.n5383 0.023
R21368 D.n5399 D.n5397 0.023
R21369 D.n5413 D.n5411 0.023
R21370 D.n5427 D.n5425 0.023
R21371 D.n5441 D.n5439 0.023
R21372 D.n5455 D.n5453 0.023
R21373 D.n5469 D.n5467 0.023
R21374 D.n5483 D.n5481 0.023
R21375 D.n5497 D.n5495 0.023
R21376 D.n5511 D.n5509 0.023
R21377 D.n5525 D.n5523 0.023
R21378 D.n5877 D.n5876 0.023
R21379 D.n5565 D.n5563 0.023
R21380 D.n5579 D.n5577 0.023
R21381 D.n5593 D.n5591 0.023
R21382 D.n5607 D.n5605 0.023
R21383 D.n5621 D.n5619 0.023
R21384 D.n5635 D.n5633 0.023
R21385 D.n5649 D.n5647 0.023
R21386 D.n5663 D.n5661 0.023
R21387 D.n5677 D.n5675 0.023
R21388 D.n5691 D.n5689 0.023
R21389 D.n5705 D.n5703 0.023
R21390 D.n5719 D.n5717 0.023
R21391 D.n5733 D.n5731 0.023
R21392 D.n5747 D.n5745 0.023
R21393 D.n5761 D.n5759 0.023
R21394 D.n5775 D.n5773 0.023
R21395 D.n5789 D.n5787 0.023
R21396 D.n5803 D.n5801 0.023
R21397 D.n5817 D.n5815 0.023
R21398 D.n5831 D.n5829 0.023
R21399 D.n5845 D.n5843 0.023
R21400 D.n5859 D.n5857 0.023
R21401 D.n5873 D.n5871 0.023
R21402 D.n6197 D.n6196 0.023
R21403 D.n5913 D.n5911 0.023
R21404 D.n5927 D.n5925 0.023
R21405 D.n5941 D.n5939 0.023
R21406 D.n5955 D.n5953 0.023
R21407 D.n5969 D.n5967 0.023
R21408 D.n5983 D.n5981 0.023
R21409 D.n5997 D.n5995 0.023
R21410 D.n6011 D.n6009 0.023
R21411 D.n6025 D.n6023 0.023
R21412 D.n6039 D.n6037 0.023
R21413 D.n6053 D.n6051 0.023
R21414 D.n6067 D.n6065 0.023
R21415 D.n6081 D.n6079 0.023
R21416 D.n6095 D.n6093 0.023
R21417 D.n6109 D.n6107 0.023
R21418 D.n6123 D.n6121 0.023
R21419 D.n6137 D.n6135 0.023
R21420 D.n6151 D.n6149 0.023
R21421 D.n6165 D.n6163 0.023
R21422 D.n6179 D.n6177 0.023
R21423 D.n6193 D.n6191 0.023
R21424 D.n6489 D.n6488 0.023
R21425 D.n6233 D.n6231 0.023
R21426 D.n6247 D.n6245 0.023
R21427 D.n6261 D.n6259 0.023
R21428 D.n6275 D.n6273 0.023
R21429 D.n6289 D.n6287 0.023
R21430 D.n6303 D.n6301 0.023
R21431 D.n6317 D.n6315 0.023
R21432 D.n6331 D.n6329 0.023
R21433 D.n6345 D.n6343 0.023
R21434 D.n6359 D.n6357 0.023
R21435 D.n6373 D.n6371 0.023
R21436 D.n6387 D.n6385 0.023
R21437 D.n6401 D.n6399 0.023
R21438 D.n6415 D.n6413 0.023
R21439 D.n6429 D.n6427 0.023
R21440 D.n6443 D.n6441 0.023
R21441 D.n6457 D.n6455 0.023
R21442 D.n6471 D.n6469 0.023
R21443 D.n6485 D.n6483 0.023
R21444 D.n6753 D.n6752 0.023
R21445 D.n6525 D.n6523 0.023
R21446 D.n6539 D.n6537 0.023
R21447 D.n6553 D.n6551 0.023
R21448 D.n6567 D.n6565 0.023
R21449 D.n6581 D.n6579 0.023
R21450 D.n6595 D.n6593 0.023
R21451 D.n6609 D.n6607 0.023
R21452 D.n6623 D.n6621 0.023
R21453 D.n6637 D.n6635 0.023
R21454 D.n6651 D.n6649 0.023
R21455 D.n6665 D.n6663 0.023
R21456 D.n6679 D.n6677 0.023
R21457 D.n6693 D.n6691 0.023
R21458 D.n6707 D.n6705 0.023
R21459 D.n6721 D.n6719 0.023
R21460 D.n6735 D.n6733 0.023
R21461 D.n6749 D.n6747 0.023
R21462 D.n6989 D.n6988 0.023
R21463 D.n6789 D.n6787 0.023
R21464 D.n6803 D.n6801 0.023
R21465 D.n6817 D.n6815 0.023
R21466 D.n6831 D.n6829 0.023
R21467 D.n6845 D.n6843 0.023
R21468 D.n6859 D.n6857 0.023
R21469 D.n6873 D.n6871 0.023
R21470 D.n6887 D.n6885 0.023
R21471 D.n6901 D.n6899 0.023
R21472 D.n6915 D.n6913 0.023
R21473 D.n6929 D.n6927 0.023
R21474 D.n6943 D.n6941 0.023
R21475 D.n6957 D.n6955 0.023
R21476 D.n6971 D.n6969 0.023
R21477 D.n6985 D.n6983 0.023
R21478 D.n7197 D.n7196 0.023
R21479 D.n7025 D.n7023 0.023
R21480 D.n7039 D.n7037 0.023
R21481 D.n7053 D.n7051 0.023
R21482 D.n7067 D.n7065 0.023
R21483 D.n7081 D.n7079 0.023
R21484 D.n7095 D.n7093 0.023
R21485 D.n7109 D.n7107 0.023
R21486 D.n7123 D.n7121 0.023
R21487 D.n7137 D.n7135 0.023
R21488 D.n7151 D.n7149 0.023
R21489 D.n7165 D.n7163 0.023
R21490 D.n7179 D.n7177 0.023
R21491 D.n7193 D.n7191 0.023
R21492 D.n7377 D.n7376 0.023
R21493 D.n7233 D.n7231 0.023
R21494 D.n7247 D.n7245 0.023
R21495 D.n7261 D.n7259 0.023
R21496 D.n7275 D.n7273 0.023
R21497 D.n7289 D.n7287 0.023
R21498 D.n7303 D.n7301 0.023
R21499 D.n7317 D.n7315 0.023
R21500 D.n7331 D.n7329 0.023
R21501 D.n7345 D.n7343 0.023
R21502 D.n7359 D.n7357 0.023
R21503 D.n7373 D.n7371 0.023
R21504 D.n7529 D.n7528 0.023
R21505 D.n7413 D.n7411 0.023
R21506 D.n7427 D.n7425 0.023
R21507 D.n7441 D.n7439 0.023
R21508 D.n7455 D.n7453 0.023
R21509 D.n7469 D.n7467 0.023
R21510 D.n7483 D.n7481 0.023
R21511 D.n7497 D.n7495 0.023
R21512 D.n7511 D.n7509 0.023
R21513 D.n7525 D.n7523 0.023
R21514 D.n7653 D.n7652 0.023
R21515 D.n7565 D.n7563 0.023
R21516 D.n7579 D.n7577 0.023
R21517 D.n7593 D.n7591 0.023
R21518 D.n7607 D.n7605 0.023
R21519 D.n7621 D.n7619 0.023
R21520 D.n7635 D.n7633 0.023
R21521 D.n7649 D.n7647 0.023
R21522 D.n7749 D.n7748 0.023
R21523 D.n7689 D.n7687 0.023
R21524 D.n7703 D.n7701 0.023
R21525 D.n7717 D.n7715 0.023
R21526 D.n7731 D.n7729 0.023
R21527 D.n7745 D.n7743 0.023
R21528 D.n7784 D.n7782 0.023
R21529 D.n7798 D.n7796 0.023
R21530 D.n7814 D.n7812 0.023
R21531 D.n7919 D.n7918 0.023
R21532 D.n7887 D.n7886 0.021
R21533 D.n7915 D.n7914 0.021
R21534 D.n46 D.n44 0.021
R21535 D.n13641 D.n13638 0.02
R21536 D.n12718 D.n12715 0.02
R21537 D.n11869 D.n11866 0.02
R21538 D.n11106 D.n11103 0.02
R21539 D.n10423 D.n10420 0.02
R21540 D.n9820 D.n9817 0.02
R21541 D.n9291 D.n9288 0.02
R21542 D.n8848 D.n8845 0.02
R21543 D.n8485 D.n8482 0.02
R21544 D.n8196 D.n8193 0.02
R21545 D.n7993 D.n7990 0.02
R21546 D.n1141 D.n512 0.019
R21547 D.n1740 D.n1142 0.019
R21548 D.n2311 D.n1741 0.019
R21549 D.n2854 D.n2312 0.019
R21550 D.n3369 D.n2855 0.019
R21551 D.n3857 D.n3371 0.019
R21552 D.n4317 D.n3859 0.019
R21553 D.n4749 D.n4319 0.019
R21554 D.n5153 D.n4751 0.019
R21555 D.n5529 D.n5155 0.019
R21556 D.n5877 D.n5531 0.019
R21557 D.n6197 D.n5879 0.019
R21558 D.n6489 D.n6199 0.019
R21559 D.n6753 D.n6491 0.019
R21560 D.n6989 D.n6755 0.019
R21561 D.n7197 D.n6991 0.019
R21562 D.n7377 D.n7199 0.019
R21563 D.n7529 D.n7379 0.019
R21564 D.n7653 D.n7531 0.019
R21565 D.n7749 D.n7655 0.019
R21566 D.n7918 D.n7917 0.017
R21567 D.n7842 D.n7841 0.016
R21568 D.n7849 D.n7848 0.016
R21569 D.n47 D.n46 0.016
R21570 D.n7933 D.n7926 0.016
R21571 D.n14096 D.n14086 0.016
R21572 D.n14096 D.n14095 0.016
R21573 D.n13183 D.n13182 0.016
R21574 D.n13184 D.n13183 0.016
R21575 D.n12300 D.n12299 0.016
R21576 D.n12301 D.n12300 0.016
R21577 D.n12248 D.n12238 0.016
R21578 D.n12248 D.n12247 0.016
R21579 D.n11449 D.n11439 0.016
R21580 D.n11449 D.n11448 0.016
R21581 D.n10730 D.n10720 0.016
R21582 D.n10730 D.n10729 0.016
R21583 D.n10125 D.n10124 0.016
R21584 D.n10126 D.n10125 0.016
R21585 D.n9562 D.n9561 0.016
R21586 D.n9563 D.n9562 0.016
R21587 D.n9526 D.n9516 0.016
R21588 D.n9526 D.n9525 0.016
R21589 D.n9047 D.n9037 0.016
R21590 D.n9047 D.n9046 0.016
R21591 D.n8670 D.n8669 0.016
R21592 D.n8671 D.n8670 0.016
R21593 D.n8347 D.n8346 0.016
R21594 D.n8348 D.n8347 0.016
R21595 D.n8323 D.n8313 0.016
R21596 D.n8323 D.n8322 0.016
R21597 D.n8084 D.n8074 0.016
R21598 D.n8084 D.n8083 0.016
R21599 D.n7934 D.n7933 0.016
R21600 D.n7917 D.n7907 0.016
R21601 D.n7917 D.n7916 0.016
R21602 D.n13698 D.n13697 0.016
R21603 D.n13716 D.n13715 0.016
R21604 D.n13734 D.n13733 0.016
R21605 D.n13752 D.n13751 0.016
R21606 D.n13770 D.n13769 0.016
R21607 D.n13788 D.n13787 0.016
R21608 D.n13806 D.n13805 0.016
R21609 D.n13824 D.n13823 0.016
R21610 D.n13842 D.n13841 0.016
R21611 D.n13860 D.n13859 0.016
R21612 D.n13878 D.n13877 0.016
R21613 D.n13896 D.n13895 0.016
R21614 D.n13914 D.n13913 0.016
R21615 D.n13932 D.n13931 0.016
R21616 D.n13950 D.n13949 0.016
R21617 D.n13968 D.n13967 0.016
R21618 D.n13986 D.n13985 0.016
R21619 D.n14004 D.n14003 0.016
R21620 D.n14022 D.n14021 0.016
R21621 D.n14040 D.n14039 0.016
R21622 D.n14058 D.n14057 0.016
R21623 D.n13602 D.n13601 0.016
R21624 D.n13582 D.n13581 0.016
R21625 D.n13562 D.n13561 0.016
R21626 D.n13542 D.n13541 0.016
R21627 D.n13522 D.n13521 0.016
R21628 D.n13502 D.n13501 0.016
R21629 D.n13482 D.n13481 0.016
R21630 D.n13462 D.n13461 0.016
R21631 D.n13442 D.n13441 0.016
R21632 D.n13422 D.n13421 0.016
R21633 D.n13402 D.n13401 0.016
R21634 D.n13382 D.n13381 0.016
R21635 D.n13362 D.n13361 0.016
R21636 D.n13342 D.n13341 0.016
R21637 D.n13322 D.n13321 0.016
R21638 D.n13302 D.n13301 0.016
R21639 D.n13282 D.n13281 0.016
R21640 D.n13262 D.n13261 0.016
R21641 D.n13242 D.n13241 0.016
R21642 D.n13222 D.n13221 0.016
R21643 D.n12771 D.n12770 0.016
R21644 D.n12789 D.n12788 0.016
R21645 D.n12807 D.n12806 0.016
R21646 D.n12825 D.n12824 0.016
R21647 D.n12843 D.n12842 0.016
R21648 D.n12861 D.n12860 0.016
R21649 D.n12879 D.n12878 0.016
R21650 D.n12897 D.n12896 0.016
R21651 D.n12915 D.n12914 0.016
R21652 D.n12933 D.n12932 0.016
R21653 D.n12951 D.n12950 0.016
R21654 D.n12969 D.n12968 0.016
R21655 D.n12987 D.n12986 0.016
R21656 D.n13005 D.n13004 0.016
R21657 D.n13023 D.n13022 0.016
R21658 D.n13041 D.n13040 0.016
R21659 D.n13059 D.n13058 0.016
R21660 D.n13077 D.n13076 0.016
R21661 D.n13095 D.n13094 0.016
R21662 D.n12679 D.n12678 0.016
R21663 D.n12659 D.n12658 0.016
R21664 D.n12639 D.n12638 0.016
R21665 D.n12619 D.n12618 0.016
R21666 D.n12599 D.n12598 0.016
R21667 D.n12579 D.n12578 0.016
R21668 D.n12559 D.n12558 0.016
R21669 D.n12539 D.n12538 0.016
R21670 D.n12519 D.n12518 0.016
R21671 D.n12499 D.n12498 0.016
R21672 D.n12479 D.n12478 0.016
R21673 D.n12459 D.n12458 0.016
R21674 D.n12439 D.n12438 0.016
R21675 D.n12419 D.n12418 0.016
R21676 D.n12399 D.n12398 0.016
R21677 D.n12379 D.n12378 0.016
R21678 D.n12359 D.n12358 0.016
R21679 D.n12339 D.n12338 0.016
R21680 D.n11922 D.n11921 0.016
R21681 D.n11940 D.n11939 0.016
R21682 D.n11958 D.n11957 0.016
R21683 D.n11976 D.n11975 0.016
R21684 D.n11994 D.n11993 0.016
R21685 D.n12012 D.n12011 0.016
R21686 D.n12030 D.n12029 0.016
R21687 D.n12048 D.n12047 0.016
R21688 D.n12066 D.n12065 0.016
R21689 D.n12084 D.n12083 0.016
R21690 D.n12102 D.n12101 0.016
R21691 D.n12120 D.n12119 0.016
R21692 D.n12138 D.n12137 0.016
R21693 D.n12156 D.n12155 0.016
R21694 D.n12174 D.n12173 0.016
R21695 D.n12192 D.n12191 0.016
R21696 D.n12210 D.n12209 0.016
R21697 D.n11830 D.n11829 0.016
R21698 D.n11810 D.n11809 0.016
R21699 D.n11790 D.n11789 0.016
R21700 D.n11770 D.n11769 0.016
R21701 D.n11750 D.n11749 0.016
R21702 D.n11730 D.n11729 0.016
R21703 D.n11710 D.n11709 0.016
R21704 D.n11690 D.n11689 0.016
R21705 D.n11670 D.n11669 0.016
R21706 D.n11650 D.n11649 0.016
R21707 D.n11630 D.n11629 0.016
R21708 D.n11610 D.n11609 0.016
R21709 D.n11590 D.n11589 0.016
R21710 D.n11570 D.n11569 0.016
R21711 D.n11550 D.n11549 0.016
R21712 D.n11530 D.n11529 0.016
R21713 D.n11159 D.n11158 0.016
R21714 D.n11177 D.n11176 0.016
R21715 D.n11195 D.n11194 0.016
R21716 D.n11213 D.n11212 0.016
R21717 D.n11231 D.n11230 0.016
R21718 D.n11249 D.n11248 0.016
R21719 D.n11267 D.n11266 0.016
R21720 D.n11285 D.n11284 0.016
R21721 D.n11303 D.n11302 0.016
R21722 D.n11321 D.n11320 0.016
R21723 D.n11339 D.n11338 0.016
R21724 D.n11357 D.n11356 0.016
R21725 D.n11375 D.n11374 0.016
R21726 D.n11393 D.n11392 0.016
R21727 D.n11411 D.n11410 0.016
R21728 D.n11067 D.n11066 0.016
R21729 D.n11047 D.n11046 0.016
R21730 D.n11027 D.n11026 0.016
R21731 D.n11007 D.n11006 0.016
R21732 D.n10987 D.n10986 0.016
R21733 D.n10967 D.n10966 0.016
R21734 D.n10947 D.n10946 0.016
R21735 D.n10927 D.n10926 0.016
R21736 D.n10907 D.n10906 0.016
R21737 D.n10887 D.n10886 0.016
R21738 D.n10867 D.n10866 0.016
R21739 D.n10847 D.n10846 0.016
R21740 D.n10827 D.n10826 0.016
R21741 D.n10807 D.n10806 0.016
R21742 D.n10476 D.n10475 0.016
R21743 D.n10494 D.n10493 0.016
R21744 D.n10512 D.n10511 0.016
R21745 D.n10530 D.n10529 0.016
R21746 D.n10548 D.n10547 0.016
R21747 D.n10566 D.n10565 0.016
R21748 D.n10584 D.n10583 0.016
R21749 D.n10602 D.n10601 0.016
R21750 D.n10620 D.n10619 0.016
R21751 D.n10638 D.n10637 0.016
R21752 D.n10656 D.n10655 0.016
R21753 D.n10674 D.n10673 0.016
R21754 D.n10692 D.n10691 0.016
R21755 D.n10384 D.n10383 0.016
R21756 D.n10364 D.n10363 0.016
R21757 D.n10344 D.n10343 0.016
R21758 D.n10324 D.n10323 0.016
R21759 D.n10304 D.n10303 0.016
R21760 D.n10284 D.n10283 0.016
R21761 D.n10264 D.n10263 0.016
R21762 D.n10244 D.n10243 0.016
R21763 D.n10224 D.n10223 0.016
R21764 D.n10204 D.n10203 0.016
R21765 D.n10184 D.n10183 0.016
R21766 D.n10164 D.n10163 0.016
R21767 D.n9873 D.n9872 0.016
R21768 D.n9891 D.n9890 0.016
R21769 D.n9909 D.n9908 0.016
R21770 D.n9927 D.n9926 0.016
R21771 D.n9945 D.n9944 0.016
R21772 D.n9963 D.n9962 0.016
R21773 D.n9981 D.n9980 0.016
R21774 D.n9999 D.n9998 0.016
R21775 D.n10017 D.n10016 0.016
R21776 D.n10035 D.n10034 0.016
R21777 D.n10053 D.n10052 0.016
R21778 D.n9781 D.n9780 0.016
R21779 D.n9761 D.n9760 0.016
R21780 D.n9741 D.n9740 0.016
R21781 D.n9721 D.n9720 0.016
R21782 D.n9701 D.n9700 0.016
R21783 D.n9681 D.n9680 0.016
R21784 D.n9661 D.n9660 0.016
R21785 D.n9641 D.n9640 0.016
R21786 D.n9621 D.n9620 0.016
R21787 D.n9601 D.n9600 0.016
R21788 D.n9344 D.n9343 0.016
R21789 D.n9362 D.n9361 0.016
R21790 D.n9380 D.n9379 0.016
R21791 D.n9398 D.n9397 0.016
R21792 D.n9416 D.n9415 0.016
R21793 D.n9434 D.n9433 0.016
R21794 D.n9452 D.n9451 0.016
R21795 D.n9470 D.n9469 0.016
R21796 D.n9488 D.n9487 0.016
R21797 D.n9252 D.n9251 0.016
R21798 D.n9232 D.n9231 0.016
R21799 D.n9212 D.n9211 0.016
R21800 D.n9192 D.n9191 0.016
R21801 D.n9172 D.n9171 0.016
R21802 D.n9152 D.n9151 0.016
R21803 D.n9132 D.n9131 0.016
R21804 D.n9112 D.n9111 0.016
R21805 D.n8901 D.n8900 0.016
R21806 D.n8919 D.n8918 0.016
R21807 D.n8937 D.n8936 0.016
R21808 D.n8955 D.n8954 0.016
R21809 D.n8973 D.n8972 0.016
R21810 D.n8991 D.n8990 0.016
R21811 D.n9009 D.n9008 0.016
R21812 D.n8809 D.n8808 0.016
R21813 D.n8789 D.n8788 0.016
R21814 D.n8769 D.n8768 0.016
R21815 D.n8749 D.n8748 0.016
R21816 D.n8729 D.n8728 0.016
R21817 D.n8709 D.n8708 0.016
R21818 D.n8538 D.n8537 0.016
R21819 D.n8556 D.n8555 0.016
R21820 D.n8574 D.n8573 0.016
R21821 D.n8592 D.n8591 0.016
R21822 D.n8610 D.n8609 0.016
R21823 D.n8446 D.n8445 0.016
R21824 D.n8426 D.n8425 0.016
R21825 D.n8406 D.n8405 0.016
R21826 D.n8386 D.n8385 0.016
R21827 D.n8249 D.n8248 0.016
R21828 D.n8267 D.n8266 0.016
R21829 D.n8285 D.n8284 0.016
R21830 D.n8157 D.n8156 0.016
R21831 D.n8137 D.n8136 0.016
R21832 D.n8046 D.n8045 0.016
R21833 D.n7962 D.n7961 0.016
R21834 D.n13689 D.n13680 0.016
R21835 D.n13707 D.n13699 0.016
R21836 D.n13725 D.n13717 0.016
R21837 D.n13743 D.n13735 0.016
R21838 D.n13761 D.n13753 0.016
R21839 D.n13779 D.n13771 0.016
R21840 D.n13797 D.n13789 0.016
R21841 D.n13815 D.n13807 0.016
R21842 D.n13833 D.n13825 0.016
R21843 D.n13851 D.n13843 0.016
R21844 D.n13869 D.n13861 0.016
R21845 D.n13887 D.n13879 0.016
R21846 D.n13905 D.n13897 0.016
R21847 D.n13923 D.n13915 0.016
R21848 D.n13941 D.n13933 0.016
R21849 D.n13959 D.n13951 0.016
R21850 D.n13977 D.n13969 0.016
R21851 D.n13995 D.n13987 0.016
R21852 D.n14013 D.n14005 0.016
R21853 D.n14031 D.n14023 0.016
R21854 D.n14049 D.n14041 0.016
R21855 D.n14067 D.n14059 0.016
R21856 D.n13612 D.n13605 0.016
R21857 D.n13592 D.n13585 0.016
R21858 D.n13572 D.n13565 0.016
R21859 D.n13552 D.n13545 0.016
R21860 D.n13532 D.n13525 0.016
R21861 D.n13512 D.n13505 0.016
R21862 D.n13492 D.n13485 0.016
R21863 D.n13472 D.n13465 0.016
R21864 D.n13452 D.n13445 0.016
R21865 D.n13432 D.n13425 0.016
R21866 D.n13412 D.n13405 0.016
R21867 D.n13392 D.n13385 0.016
R21868 D.n13372 D.n13365 0.016
R21869 D.n13352 D.n13345 0.016
R21870 D.n13332 D.n13325 0.016
R21871 D.n13312 D.n13305 0.016
R21872 D.n13292 D.n13285 0.016
R21873 D.n13272 D.n13265 0.016
R21874 D.n13252 D.n13245 0.016
R21875 D.n13232 D.n13225 0.016
R21876 D.n13212 D.n13205 0.016
R21877 D.n12762 D.n12753 0.016
R21878 D.n12780 D.n12772 0.016
R21879 D.n12798 D.n12790 0.016
R21880 D.n12816 D.n12808 0.016
R21881 D.n12834 D.n12826 0.016
R21882 D.n12852 D.n12844 0.016
R21883 D.n12870 D.n12862 0.016
R21884 D.n12888 D.n12880 0.016
R21885 D.n12906 D.n12898 0.016
R21886 D.n12924 D.n12916 0.016
R21887 D.n12942 D.n12934 0.016
R21888 D.n12960 D.n12952 0.016
R21889 D.n12978 D.n12970 0.016
R21890 D.n12996 D.n12988 0.016
R21891 D.n13014 D.n13006 0.016
R21892 D.n13032 D.n13024 0.016
R21893 D.n13050 D.n13042 0.016
R21894 D.n13068 D.n13060 0.016
R21895 D.n13086 D.n13078 0.016
R21896 D.n13104 D.n13096 0.016
R21897 D.n12689 D.n12682 0.016
R21898 D.n12669 D.n12662 0.016
R21899 D.n12649 D.n12642 0.016
R21900 D.n12629 D.n12622 0.016
R21901 D.n12609 D.n12602 0.016
R21902 D.n12589 D.n12582 0.016
R21903 D.n12569 D.n12562 0.016
R21904 D.n12549 D.n12542 0.016
R21905 D.n12529 D.n12522 0.016
R21906 D.n12509 D.n12502 0.016
R21907 D.n12489 D.n12482 0.016
R21908 D.n12469 D.n12462 0.016
R21909 D.n12449 D.n12442 0.016
R21910 D.n12429 D.n12422 0.016
R21911 D.n12409 D.n12402 0.016
R21912 D.n12389 D.n12382 0.016
R21913 D.n12369 D.n12362 0.016
R21914 D.n12349 D.n12342 0.016
R21915 D.n12329 D.n12322 0.016
R21916 D.n11913 D.n11904 0.016
R21917 D.n11931 D.n11923 0.016
R21918 D.n11949 D.n11941 0.016
R21919 D.n11967 D.n11959 0.016
R21920 D.n11985 D.n11977 0.016
R21921 D.n12003 D.n11995 0.016
R21922 D.n12021 D.n12013 0.016
R21923 D.n12039 D.n12031 0.016
R21924 D.n12057 D.n12049 0.016
R21925 D.n12075 D.n12067 0.016
R21926 D.n12093 D.n12085 0.016
R21927 D.n12111 D.n12103 0.016
R21928 D.n12129 D.n12121 0.016
R21929 D.n12147 D.n12139 0.016
R21930 D.n12165 D.n12157 0.016
R21931 D.n12183 D.n12175 0.016
R21932 D.n12201 D.n12193 0.016
R21933 D.n12219 D.n12211 0.016
R21934 D.n11840 D.n11833 0.016
R21935 D.n11820 D.n11813 0.016
R21936 D.n11800 D.n11793 0.016
R21937 D.n11780 D.n11773 0.016
R21938 D.n11760 D.n11753 0.016
R21939 D.n11740 D.n11733 0.016
R21940 D.n11720 D.n11713 0.016
R21941 D.n11700 D.n11693 0.016
R21942 D.n11680 D.n11673 0.016
R21943 D.n11660 D.n11653 0.016
R21944 D.n11640 D.n11633 0.016
R21945 D.n11620 D.n11613 0.016
R21946 D.n11600 D.n11593 0.016
R21947 D.n11580 D.n11573 0.016
R21948 D.n11560 D.n11553 0.016
R21949 D.n11540 D.n11533 0.016
R21950 D.n11520 D.n11513 0.016
R21951 D.n11150 D.n11141 0.016
R21952 D.n11168 D.n11160 0.016
R21953 D.n11186 D.n11178 0.016
R21954 D.n11204 D.n11196 0.016
R21955 D.n11222 D.n11214 0.016
R21956 D.n11240 D.n11232 0.016
R21957 D.n11258 D.n11250 0.016
R21958 D.n11276 D.n11268 0.016
R21959 D.n11294 D.n11286 0.016
R21960 D.n11312 D.n11304 0.016
R21961 D.n11330 D.n11322 0.016
R21962 D.n11348 D.n11340 0.016
R21963 D.n11366 D.n11358 0.016
R21964 D.n11384 D.n11376 0.016
R21965 D.n11402 D.n11394 0.016
R21966 D.n11420 D.n11412 0.016
R21967 D.n11077 D.n11070 0.016
R21968 D.n11057 D.n11050 0.016
R21969 D.n11037 D.n11030 0.016
R21970 D.n11017 D.n11010 0.016
R21971 D.n10997 D.n10990 0.016
R21972 D.n10977 D.n10970 0.016
R21973 D.n10957 D.n10950 0.016
R21974 D.n10937 D.n10930 0.016
R21975 D.n10917 D.n10910 0.016
R21976 D.n10897 D.n10890 0.016
R21977 D.n10877 D.n10870 0.016
R21978 D.n10857 D.n10850 0.016
R21979 D.n10837 D.n10830 0.016
R21980 D.n10817 D.n10810 0.016
R21981 D.n10797 D.n10790 0.016
R21982 D.n10467 D.n10458 0.016
R21983 D.n10485 D.n10477 0.016
R21984 D.n10503 D.n10495 0.016
R21985 D.n10521 D.n10513 0.016
R21986 D.n10539 D.n10531 0.016
R21987 D.n10557 D.n10549 0.016
R21988 D.n10575 D.n10567 0.016
R21989 D.n10593 D.n10585 0.016
R21990 D.n10611 D.n10603 0.016
R21991 D.n10629 D.n10621 0.016
R21992 D.n10647 D.n10639 0.016
R21993 D.n10665 D.n10657 0.016
R21994 D.n10683 D.n10675 0.016
R21995 D.n10701 D.n10693 0.016
R21996 D.n10394 D.n10387 0.016
R21997 D.n10374 D.n10367 0.016
R21998 D.n10354 D.n10347 0.016
R21999 D.n10334 D.n10327 0.016
R22000 D.n10314 D.n10307 0.016
R22001 D.n10294 D.n10287 0.016
R22002 D.n10274 D.n10267 0.016
R22003 D.n10254 D.n10247 0.016
R22004 D.n10234 D.n10227 0.016
R22005 D.n10214 D.n10207 0.016
R22006 D.n10194 D.n10187 0.016
R22007 D.n10174 D.n10167 0.016
R22008 D.n10154 D.n10147 0.016
R22009 D.n9864 D.n9855 0.016
R22010 D.n9882 D.n9874 0.016
R22011 D.n9900 D.n9892 0.016
R22012 D.n9918 D.n9910 0.016
R22013 D.n9936 D.n9928 0.016
R22014 D.n9954 D.n9946 0.016
R22015 D.n9972 D.n9964 0.016
R22016 D.n9990 D.n9982 0.016
R22017 D.n10008 D.n10000 0.016
R22018 D.n10026 D.n10018 0.016
R22019 D.n10044 D.n10036 0.016
R22020 D.n10062 D.n10054 0.016
R22021 D.n9791 D.n9784 0.016
R22022 D.n9771 D.n9764 0.016
R22023 D.n9751 D.n9744 0.016
R22024 D.n9731 D.n9724 0.016
R22025 D.n9711 D.n9704 0.016
R22026 D.n9691 D.n9684 0.016
R22027 D.n9671 D.n9664 0.016
R22028 D.n9651 D.n9644 0.016
R22029 D.n9631 D.n9624 0.016
R22030 D.n9611 D.n9604 0.016
R22031 D.n9591 D.n9584 0.016
R22032 D.n9335 D.n9326 0.016
R22033 D.n9353 D.n9345 0.016
R22034 D.n9371 D.n9363 0.016
R22035 D.n9389 D.n9381 0.016
R22036 D.n9407 D.n9399 0.016
R22037 D.n9425 D.n9417 0.016
R22038 D.n9443 D.n9435 0.016
R22039 D.n9461 D.n9453 0.016
R22040 D.n9479 D.n9471 0.016
R22041 D.n9497 D.n9489 0.016
R22042 D.n9262 D.n9255 0.016
R22043 D.n9242 D.n9235 0.016
R22044 D.n9222 D.n9215 0.016
R22045 D.n9202 D.n9195 0.016
R22046 D.n9182 D.n9175 0.016
R22047 D.n9162 D.n9155 0.016
R22048 D.n9142 D.n9135 0.016
R22049 D.n9122 D.n9115 0.016
R22050 D.n9102 D.n9095 0.016
R22051 D.n8892 D.n8883 0.016
R22052 D.n8910 D.n8902 0.016
R22053 D.n8928 D.n8920 0.016
R22054 D.n8946 D.n8938 0.016
R22055 D.n8964 D.n8956 0.016
R22056 D.n8982 D.n8974 0.016
R22057 D.n9000 D.n8992 0.016
R22058 D.n9018 D.n9010 0.016
R22059 D.n8819 D.n8812 0.016
R22060 D.n8799 D.n8792 0.016
R22061 D.n8779 D.n8772 0.016
R22062 D.n8759 D.n8752 0.016
R22063 D.n8739 D.n8732 0.016
R22064 D.n8719 D.n8712 0.016
R22065 D.n8699 D.n8692 0.016
R22066 D.n8529 D.n8520 0.016
R22067 D.n8547 D.n8539 0.016
R22068 D.n8565 D.n8557 0.016
R22069 D.n8583 D.n8575 0.016
R22070 D.n8601 D.n8593 0.016
R22071 D.n8619 D.n8611 0.016
R22072 D.n8456 D.n8449 0.016
R22073 D.n8436 D.n8429 0.016
R22074 D.n8416 D.n8409 0.016
R22075 D.n8396 D.n8389 0.016
R22076 D.n8376 D.n8369 0.016
R22077 D.n8240 D.n8231 0.016
R22078 D.n8258 D.n8250 0.016
R22079 D.n8276 D.n8268 0.016
R22080 D.n8294 D.n8286 0.016
R22081 D.n8167 D.n8160 0.016
R22082 D.n8147 D.n8140 0.016
R22083 D.n8127 D.n8120 0.016
R22084 D.n8037 D.n8028 0.016
R22085 D.n8055 D.n8047 0.016
R22086 D.n57 D.n56 0.016
R22087 D.n66 D.n65 0.016
R22088 D.n75 D.n74 0.016
R22089 D.n84 D.n83 0.016
R22090 D.n93 D.n92 0.016
R22091 D.n102 D.n101 0.016
R22092 D.n111 D.n110 0.016
R22093 D.n120 D.n119 0.016
R22094 D.n129 D.n128 0.016
R22095 D.n138 D.n137 0.016
R22096 D.n147 D.n146 0.016
R22097 D.n156 D.n155 0.016
R22098 D.n165 D.n164 0.016
R22099 D.n174 D.n173 0.016
R22100 D.n183 D.n182 0.016
R22101 D.n192 D.n191 0.016
R22102 D.n201 D.n200 0.016
R22103 D.n210 D.n209 0.016
R22104 D.n219 D.n218 0.016
R22105 D.n228 D.n227 0.016
R22106 D.n237 D.n236 0.016
R22107 D.n246 D.n245 0.016
R22108 D.n255 D.n254 0.016
R22109 D.n264 D.n263 0.016
R22110 D.n273 D.n272 0.016
R22111 D.n282 D.n281 0.016
R22112 D.n291 D.n290 0.016
R22113 D.n300 D.n299 0.016
R22114 D.n309 D.n308 0.016
R22115 D.n318 D.n317 0.016
R22116 D.n327 D.n326 0.016
R22117 D.n336 D.n335 0.016
R22118 D.n345 D.n344 0.016
R22119 D.n354 D.n353 0.016
R22120 D.n363 D.n362 0.016
R22121 D.n372 D.n371 0.016
R22122 D.n381 D.n380 0.016
R22123 D.n390 D.n389 0.016
R22124 D.n399 D.n398 0.016
R22125 D.n408 D.n407 0.016
R22126 D.n417 D.n416 0.016
R22127 D.n426 D.n425 0.016
R22128 D.n435 D.n434 0.016
R22129 D.n1137 D.n1125 0.016
R22130 D.n1123 D.n1111 0.016
R22131 D.n1109 D.n1097 0.016
R22132 D.n1095 D.n1083 0.016
R22133 D.n1081 D.n1069 0.016
R22134 D.n1067 D.n1055 0.016
R22135 D.n1053 D.n1041 0.016
R22136 D.n1039 D.n1027 0.016
R22137 D.n1025 D.n1013 0.016
R22138 D.n1011 D.n999 0.016
R22139 D.n997 D.n985 0.016
R22140 D.n983 D.n971 0.016
R22141 D.n969 D.n957 0.016
R22142 D.n955 D.n943 0.016
R22143 D.n941 D.n929 0.016
R22144 D.n927 D.n915 0.016
R22145 D.n913 D.n901 0.016
R22146 D.n899 D.n887 0.016
R22147 D.n885 D.n873 0.016
R22148 D.n871 D.n859 0.016
R22149 D.n857 D.n845 0.016
R22150 D.n843 D.n831 0.016
R22151 D.n829 D.n817 0.016
R22152 D.n815 D.n803 0.016
R22153 D.n801 D.n789 0.016
R22154 D.n787 D.n775 0.016
R22155 D.n773 D.n761 0.016
R22156 D.n759 D.n747 0.016
R22157 D.n745 D.n733 0.016
R22158 D.n731 D.n719 0.016
R22159 D.n717 D.n705 0.016
R22160 D.n703 D.n691 0.016
R22161 D.n689 D.n677 0.016
R22162 D.n675 D.n663 0.016
R22163 D.n661 D.n649 0.016
R22164 D.n647 D.n635 0.016
R22165 D.n633 D.n621 0.016
R22166 D.n619 D.n607 0.016
R22167 D.n605 D.n593 0.016
R22168 D.n591 D.n579 0.016
R22169 D.n577 D.n565 0.016
R22170 D.n563 D.n551 0.016
R22171 D.n1736 D.n1724 0.016
R22172 D.n1722 D.n1710 0.016
R22173 D.n1708 D.n1696 0.016
R22174 D.n1694 D.n1682 0.016
R22175 D.n1680 D.n1668 0.016
R22176 D.n1666 D.n1654 0.016
R22177 D.n1652 D.n1640 0.016
R22178 D.n1638 D.n1626 0.016
R22179 D.n1624 D.n1612 0.016
R22180 D.n1610 D.n1598 0.016
R22181 D.n1596 D.n1584 0.016
R22182 D.n1582 D.n1570 0.016
R22183 D.n1568 D.n1556 0.016
R22184 D.n1554 D.n1542 0.016
R22185 D.n1540 D.n1528 0.016
R22186 D.n1526 D.n1514 0.016
R22187 D.n1512 D.n1500 0.016
R22188 D.n1498 D.n1486 0.016
R22189 D.n1484 D.n1472 0.016
R22190 D.n1470 D.n1458 0.016
R22191 D.n1456 D.n1444 0.016
R22192 D.n1442 D.n1430 0.016
R22193 D.n1428 D.n1416 0.016
R22194 D.n1414 D.n1402 0.016
R22195 D.n1400 D.n1388 0.016
R22196 D.n1386 D.n1374 0.016
R22197 D.n1372 D.n1360 0.016
R22198 D.n1358 D.n1346 0.016
R22199 D.n1344 D.n1332 0.016
R22200 D.n1330 D.n1318 0.016
R22201 D.n1316 D.n1304 0.016
R22202 D.n1302 D.n1290 0.016
R22203 D.n1288 D.n1276 0.016
R22204 D.n1274 D.n1262 0.016
R22205 D.n1260 D.n1248 0.016
R22206 D.n1246 D.n1234 0.016
R22207 D.n1232 D.n1220 0.016
R22208 D.n1218 D.n1206 0.016
R22209 D.n1204 D.n1192 0.016
R22210 D.n1190 D.n1178 0.016
R22211 D.n2307 D.n2295 0.016
R22212 D.n2293 D.n2281 0.016
R22213 D.n2279 D.n2267 0.016
R22214 D.n2265 D.n2253 0.016
R22215 D.n2251 D.n2239 0.016
R22216 D.n2237 D.n2225 0.016
R22217 D.n2223 D.n2211 0.016
R22218 D.n2209 D.n2197 0.016
R22219 D.n2195 D.n2183 0.016
R22220 D.n2181 D.n2169 0.016
R22221 D.n2167 D.n2155 0.016
R22222 D.n2153 D.n2141 0.016
R22223 D.n2139 D.n2127 0.016
R22224 D.n2125 D.n2113 0.016
R22225 D.n2111 D.n2099 0.016
R22226 D.n2097 D.n2085 0.016
R22227 D.n2083 D.n2071 0.016
R22228 D.n2069 D.n2057 0.016
R22229 D.n2055 D.n2043 0.016
R22230 D.n2041 D.n2029 0.016
R22231 D.n2027 D.n2015 0.016
R22232 D.n2013 D.n2001 0.016
R22233 D.n1999 D.n1987 0.016
R22234 D.n1985 D.n1973 0.016
R22235 D.n1971 D.n1959 0.016
R22236 D.n1957 D.n1945 0.016
R22237 D.n1943 D.n1931 0.016
R22238 D.n1929 D.n1917 0.016
R22239 D.n1915 D.n1903 0.016
R22240 D.n1901 D.n1889 0.016
R22241 D.n1887 D.n1875 0.016
R22242 D.n1873 D.n1861 0.016
R22243 D.n1859 D.n1847 0.016
R22244 D.n1845 D.n1833 0.016
R22245 D.n1831 D.n1819 0.016
R22246 D.n1817 D.n1805 0.016
R22247 D.n1803 D.n1791 0.016
R22248 D.n1789 D.n1777 0.016
R22249 D.n2850 D.n2838 0.016
R22250 D.n2836 D.n2824 0.016
R22251 D.n2822 D.n2810 0.016
R22252 D.n2808 D.n2796 0.016
R22253 D.n2794 D.n2782 0.016
R22254 D.n2780 D.n2768 0.016
R22255 D.n2766 D.n2754 0.016
R22256 D.n2752 D.n2740 0.016
R22257 D.n2738 D.n2726 0.016
R22258 D.n2724 D.n2712 0.016
R22259 D.n2710 D.n2698 0.016
R22260 D.n2696 D.n2684 0.016
R22261 D.n2682 D.n2670 0.016
R22262 D.n2668 D.n2656 0.016
R22263 D.n2654 D.n2642 0.016
R22264 D.n2640 D.n2628 0.016
R22265 D.n2626 D.n2614 0.016
R22266 D.n2612 D.n2600 0.016
R22267 D.n2598 D.n2586 0.016
R22268 D.n2584 D.n2572 0.016
R22269 D.n2570 D.n2558 0.016
R22270 D.n2556 D.n2544 0.016
R22271 D.n2542 D.n2530 0.016
R22272 D.n2528 D.n2516 0.016
R22273 D.n2514 D.n2502 0.016
R22274 D.n2500 D.n2488 0.016
R22275 D.n2486 D.n2474 0.016
R22276 D.n2472 D.n2460 0.016
R22277 D.n2458 D.n2446 0.016
R22278 D.n2444 D.n2432 0.016
R22279 D.n2430 D.n2418 0.016
R22280 D.n2416 D.n2404 0.016
R22281 D.n2402 D.n2390 0.016
R22282 D.n2388 D.n2376 0.016
R22283 D.n2374 D.n2362 0.016
R22284 D.n2360 D.n2348 0.016
R22285 D.n3365 D.n3353 0.016
R22286 D.n3351 D.n3339 0.016
R22287 D.n3337 D.n3325 0.016
R22288 D.n3323 D.n3311 0.016
R22289 D.n3309 D.n3297 0.016
R22290 D.n3295 D.n3283 0.016
R22291 D.n3281 D.n3269 0.016
R22292 D.n3267 D.n3255 0.016
R22293 D.n3253 D.n3241 0.016
R22294 D.n3239 D.n3227 0.016
R22295 D.n3225 D.n3213 0.016
R22296 D.n3211 D.n3199 0.016
R22297 D.n3197 D.n3185 0.016
R22298 D.n3183 D.n3171 0.016
R22299 D.n3169 D.n3157 0.016
R22300 D.n3155 D.n3143 0.016
R22301 D.n3141 D.n3129 0.016
R22302 D.n3127 D.n3115 0.016
R22303 D.n3113 D.n3101 0.016
R22304 D.n3099 D.n3087 0.016
R22305 D.n3085 D.n3073 0.016
R22306 D.n3071 D.n3059 0.016
R22307 D.n3057 D.n3045 0.016
R22308 D.n3043 D.n3031 0.016
R22309 D.n3029 D.n3017 0.016
R22310 D.n3015 D.n3003 0.016
R22311 D.n3001 D.n2989 0.016
R22312 D.n2987 D.n2975 0.016
R22313 D.n2973 D.n2961 0.016
R22314 D.n2959 D.n2947 0.016
R22315 D.n2945 D.n2933 0.016
R22316 D.n2931 D.n2919 0.016
R22317 D.n2917 D.n2905 0.016
R22318 D.n2903 D.n2891 0.016
R22319 D.n3853 D.n3841 0.016
R22320 D.n3839 D.n3827 0.016
R22321 D.n3825 D.n3813 0.016
R22322 D.n3811 D.n3799 0.016
R22323 D.n3797 D.n3785 0.016
R22324 D.n3783 D.n3771 0.016
R22325 D.n3769 D.n3757 0.016
R22326 D.n3755 D.n3743 0.016
R22327 D.n3741 D.n3729 0.016
R22328 D.n3727 D.n3715 0.016
R22329 D.n3713 D.n3701 0.016
R22330 D.n3699 D.n3687 0.016
R22331 D.n3685 D.n3673 0.016
R22332 D.n3671 D.n3659 0.016
R22333 D.n3657 D.n3645 0.016
R22334 D.n3643 D.n3631 0.016
R22335 D.n3629 D.n3617 0.016
R22336 D.n3615 D.n3603 0.016
R22337 D.n3601 D.n3589 0.016
R22338 D.n3587 D.n3575 0.016
R22339 D.n3573 D.n3561 0.016
R22340 D.n3559 D.n3547 0.016
R22341 D.n3545 D.n3533 0.016
R22342 D.n3531 D.n3519 0.016
R22343 D.n3517 D.n3505 0.016
R22344 D.n3503 D.n3491 0.016
R22345 D.n3489 D.n3477 0.016
R22346 D.n3475 D.n3463 0.016
R22347 D.n3461 D.n3449 0.016
R22348 D.n3447 D.n3435 0.016
R22349 D.n3433 D.n3421 0.016
R22350 D.n3419 D.n3407 0.016
R22351 D.n4313 D.n4301 0.016
R22352 D.n4299 D.n4287 0.016
R22353 D.n4285 D.n4273 0.016
R22354 D.n4271 D.n4259 0.016
R22355 D.n4257 D.n4245 0.016
R22356 D.n4243 D.n4231 0.016
R22357 D.n4229 D.n4217 0.016
R22358 D.n4215 D.n4203 0.016
R22359 D.n4201 D.n4189 0.016
R22360 D.n4187 D.n4175 0.016
R22361 D.n4173 D.n4161 0.016
R22362 D.n4159 D.n4147 0.016
R22363 D.n4145 D.n4133 0.016
R22364 D.n4131 D.n4119 0.016
R22365 D.n4117 D.n4105 0.016
R22366 D.n4103 D.n4091 0.016
R22367 D.n4089 D.n4077 0.016
R22368 D.n4075 D.n4063 0.016
R22369 D.n4061 D.n4049 0.016
R22370 D.n4047 D.n4035 0.016
R22371 D.n4033 D.n4021 0.016
R22372 D.n4019 D.n4007 0.016
R22373 D.n4005 D.n3993 0.016
R22374 D.n3991 D.n3979 0.016
R22375 D.n3977 D.n3965 0.016
R22376 D.n3963 D.n3951 0.016
R22377 D.n3949 D.n3937 0.016
R22378 D.n3935 D.n3923 0.016
R22379 D.n3921 D.n3909 0.016
R22380 D.n3907 D.n3895 0.016
R22381 D.n4745 D.n4733 0.016
R22382 D.n4731 D.n4719 0.016
R22383 D.n4717 D.n4705 0.016
R22384 D.n4703 D.n4691 0.016
R22385 D.n4689 D.n4677 0.016
R22386 D.n4675 D.n4663 0.016
R22387 D.n4661 D.n4649 0.016
R22388 D.n4647 D.n4635 0.016
R22389 D.n4633 D.n4621 0.016
R22390 D.n4619 D.n4607 0.016
R22391 D.n4605 D.n4593 0.016
R22392 D.n4591 D.n4579 0.016
R22393 D.n4577 D.n4565 0.016
R22394 D.n4563 D.n4551 0.016
R22395 D.n4549 D.n4537 0.016
R22396 D.n4535 D.n4523 0.016
R22397 D.n4521 D.n4509 0.016
R22398 D.n4507 D.n4495 0.016
R22399 D.n4493 D.n4481 0.016
R22400 D.n4479 D.n4467 0.016
R22401 D.n4465 D.n4453 0.016
R22402 D.n4451 D.n4439 0.016
R22403 D.n4437 D.n4425 0.016
R22404 D.n4423 D.n4411 0.016
R22405 D.n4409 D.n4397 0.016
R22406 D.n4395 D.n4383 0.016
R22407 D.n4381 D.n4369 0.016
R22408 D.n4367 D.n4355 0.016
R22409 D.n5149 D.n5137 0.016
R22410 D.n5135 D.n5123 0.016
R22411 D.n5121 D.n5109 0.016
R22412 D.n5107 D.n5095 0.016
R22413 D.n5093 D.n5081 0.016
R22414 D.n5079 D.n5067 0.016
R22415 D.n5065 D.n5053 0.016
R22416 D.n5051 D.n5039 0.016
R22417 D.n5037 D.n5025 0.016
R22418 D.n5023 D.n5011 0.016
R22419 D.n5009 D.n4997 0.016
R22420 D.n4995 D.n4983 0.016
R22421 D.n4981 D.n4969 0.016
R22422 D.n4967 D.n4955 0.016
R22423 D.n4953 D.n4941 0.016
R22424 D.n4939 D.n4927 0.016
R22425 D.n4925 D.n4913 0.016
R22426 D.n4911 D.n4899 0.016
R22427 D.n4897 D.n4885 0.016
R22428 D.n4883 D.n4871 0.016
R22429 D.n4869 D.n4857 0.016
R22430 D.n4855 D.n4843 0.016
R22431 D.n4841 D.n4829 0.016
R22432 D.n4827 D.n4815 0.016
R22433 D.n4813 D.n4801 0.016
R22434 D.n4799 D.n4787 0.016
R22435 D.n5525 D.n5513 0.016
R22436 D.n5511 D.n5499 0.016
R22437 D.n5497 D.n5485 0.016
R22438 D.n5483 D.n5471 0.016
R22439 D.n5469 D.n5457 0.016
R22440 D.n5455 D.n5443 0.016
R22441 D.n5441 D.n5429 0.016
R22442 D.n5427 D.n5415 0.016
R22443 D.n5413 D.n5401 0.016
R22444 D.n5399 D.n5387 0.016
R22445 D.n5385 D.n5373 0.016
R22446 D.n5371 D.n5359 0.016
R22447 D.n5357 D.n5345 0.016
R22448 D.n5343 D.n5331 0.016
R22449 D.n5329 D.n5317 0.016
R22450 D.n5315 D.n5303 0.016
R22451 D.n5301 D.n5289 0.016
R22452 D.n5287 D.n5275 0.016
R22453 D.n5273 D.n5261 0.016
R22454 D.n5259 D.n5247 0.016
R22455 D.n5245 D.n5233 0.016
R22456 D.n5231 D.n5219 0.016
R22457 D.n5217 D.n5205 0.016
R22458 D.n5203 D.n5191 0.016
R22459 D.n5873 D.n5861 0.016
R22460 D.n5859 D.n5847 0.016
R22461 D.n5845 D.n5833 0.016
R22462 D.n5831 D.n5819 0.016
R22463 D.n5817 D.n5805 0.016
R22464 D.n5803 D.n5791 0.016
R22465 D.n5789 D.n5777 0.016
R22466 D.n5775 D.n5763 0.016
R22467 D.n5761 D.n5749 0.016
R22468 D.n5747 D.n5735 0.016
R22469 D.n5733 D.n5721 0.016
R22470 D.n5719 D.n5707 0.016
R22471 D.n5705 D.n5693 0.016
R22472 D.n5691 D.n5679 0.016
R22473 D.n5677 D.n5665 0.016
R22474 D.n5663 D.n5651 0.016
R22475 D.n5649 D.n5637 0.016
R22476 D.n5635 D.n5623 0.016
R22477 D.n5621 D.n5609 0.016
R22478 D.n5607 D.n5595 0.016
R22479 D.n5593 D.n5581 0.016
R22480 D.n5579 D.n5567 0.016
R22481 D.n6193 D.n6181 0.016
R22482 D.n6179 D.n6167 0.016
R22483 D.n6165 D.n6153 0.016
R22484 D.n6151 D.n6139 0.016
R22485 D.n6137 D.n6125 0.016
R22486 D.n6123 D.n6111 0.016
R22487 D.n6109 D.n6097 0.016
R22488 D.n6095 D.n6083 0.016
R22489 D.n6081 D.n6069 0.016
R22490 D.n6067 D.n6055 0.016
R22491 D.n6053 D.n6041 0.016
R22492 D.n6039 D.n6027 0.016
R22493 D.n6025 D.n6013 0.016
R22494 D.n6011 D.n5999 0.016
R22495 D.n5997 D.n5985 0.016
R22496 D.n5983 D.n5971 0.016
R22497 D.n5969 D.n5957 0.016
R22498 D.n5955 D.n5943 0.016
R22499 D.n5941 D.n5929 0.016
R22500 D.n5927 D.n5915 0.016
R22501 D.n6485 D.n6473 0.016
R22502 D.n6471 D.n6459 0.016
R22503 D.n6457 D.n6445 0.016
R22504 D.n6443 D.n6431 0.016
R22505 D.n6429 D.n6417 0.016
R22506 D.n6415 D.n6403 0.016
R22507 D.n6401 D.n6389 0.016
R22508 D.n6387 D.n6375 0.016
R22509 D.n6373 D.n6361 0.016
R22510 D.n6359 D.n6347 0.016
R22511 D.n6345 D.n6333 0.016
R22512 D.n6331 D.n6319 0.016
R22513 D.n6317 D.n6305 0.016
R22514 D.n6303 D.n6291 0.016
R22515 D.n6289 D.n6277 0.016
R22516 D.n6275 D.n6263 0.016
R22517 D.n6261 D.n6249 0.016
R22518 D.n6247 D.n6235 0.016
R22519 D.n6749 D.n6737 0.016
R22520 D.n6735 D.n6723 0.016
R22521 D.n6721 D.n6709 0.016
R22522 D.n6707 D.n6695 0.016
R22523 D.n6693 D.n6681 0.016
R22524 D.n6679 D.n6667 0.016
R22525 D.n6665 D.n6653 0.016
R22526 D.n6651 D.n6639 0.016
R22527 D.n6637 D.n6625 0.016
R22528 D.n6623 D.n6611 0.016
R22529 D.n6609 D.n6597 0.016
R22530 D.n6595 D.n6583 0.016
R22531 D.n6581 D.n6569 0.016
R22532 D.n6567 D.n6555 0.016
R22533 D.n6553 D.n6541 0.016
R22534 D.n6539 D.n6527 0.016
R22535 D.n6985 D.n6973 0.016
R22536 D.n6971 D.n6959 0.016
R22537 D.n6957 D.n6945 0.016
R22538 D.n6943 D.n6931 0.016
R22539 D.n6929 D.n6917 0.016
R22540 D.n6915 D.n6903 0.016
R22541 D.n6901 D.n6889 0.016
R22542 D.n6887 D.n6875 0.016
R22543 D.n6873 D.n6861 0.016
R22544 D.n6859 D.n6847 0.016
R22545 D.n6845 D.n6833 0.016
R22546 D.n6831 D.n6819 0.016
R22547 D.n6817 D.n6805 0.016
R22548 D.n6803 D.n6791 0.016
R22549 D.n7193 D.n7181 0.016
R22550 D.n7179 D.n7167 0.016
R22551 D.n7165 D.n7153 0.016
R22552 D.n7151 D.n7139 0.016
R22553 D.n7137 D.n7125 0.016
R22554 D.n7123 D.n7111 0.016
R22555 D.n7109 D.n7097 0.016
R22556 D.n7095 D.n7083 0.016
R22557 D.n7081 D.n7069 0.016
R22558 D.n7067 D.n7055 0.016
R22559 D.n7053 D.n7041 0.016
R22560 D.n7039 D.n7027 0.016
R22561 D.n7373 D.n7361 0.016
R22562 D.n7359 D.n7347 0.016
R22563 D.n7345 D.n7333 0.016
R22564 D.n7331 D.n7319 0.016
R22565 D.n7317 D.n7305 0.016
R22566 D.n7303 D.n7291 0.016
R22567 D.n7289 D.n7277 0.016
R22568 D.n7275 D.n7263 0.016
R22569 D.n7261 D.n7249 0.016
R22570 D.n7247 D.n7235 0.016
R22571 D.n7525 D.n7513 0.016
R22572 D.n7511 D.n7499 0.016
R22573 D.n7497 D.n7485 0.016
R22574 D.n7483 D.n7471 0.016
R22575 D.n7469 D.n7457 0.016
R22576 D.n7455 D.n7443 0.016
R22577 D.n7441 D.n7429 0.016
R22578 D.n7427 D.n7415 0.016
R22579 D.n7649 D.n7637 0.016
R22580 D.n7635 D.n7623 0.016
R22581 D.n7621 D.n7609 0.016
R22582 D.n7607 D.n7595 0.016
R22583 D.n7593 D.n7581 0.016
R22584 D.n7579 D.n7567 0.016
R22585 D.n7745 D.n7733 0.016
R22586 D.n7731 D.n7719 0.016
R22587 D.n7717 D.n7705 0.016
R22588 D.n7703 D.n7691 0.016
R22589 D.n7814 D.n7800 0.016
R22590 D.n7798 D.n7786 0.016
R22591 D.n1141 D.n520 0.016
R22592 D.n1740 D.n1147 0.016
R22593 D.n2311 D.n1746 0.016
R22594 D.n2854 D.n2317 0.016
R22595 D.n3369 D.n2860 0.016
R22596 D.n3857 D.n3376 0.016
R22597 D.n4317 D.n3864 0.016
R22598 D.n4749 D.n4324 0.016
R22599 D.n5153 D.n4756 0.016
R22600 D.n5529 D.n5160 0.016
R22601 D.n5877 D.n5536 0.016
R22602 D.n6197 D.n5884 0.016
R22603 D.n6489 D.n6204 0.016
R22604 D.n6753 D.n6496 0.016
R22605 D.n6989 D.n6760 0.016
R22606 D.n7197 D.n6996 0.016
R22607 D.n7377 D.n7204 0.016
R22608 D.n7529 D.n7384 0.016
R22609 D.n7653 D.n7536 0.016
R22610 D.n7749 D.n7660 0.016
R22611 D.n7816 D.n7755 0.016
R22612 D.n7849 D.n7846 0.016
R22613 D.n7856 D.n7851 0.016
R22614 D.n7856 D.n7855 0.016
R22615 D.n13172 D.n13171 0.015
R22616 D.n12289 D.n12288 0.015
R22617 D.n11486 D.n11485 0.015
R22618 D.n10763 D.n10762 0.015
R22619 D.n10114 D.n10113 0.015
R22620 D.n9551 D.n9550 0.015
R22621 D.n9068 D.n9067 0.015
R22622 D.n8659 D.n8658 0.015
R22623 D.n8336 D.n8335 0.015
R22624 D.n8093 D.n8092 0.015
R22625 D.n7975 D.n7974 0.015
R22626 D.n7949 D.n7948 0.015
R22627 D.n14085 D.n14084 0.015
R22628 D.n14070 D.n14069 0.015
R22629 D.n13199 D.n13198 0.015
R22630 D.n13187 D.n13185 0.015
R22631 D.n13126 D.n13125 0.015
R22632 D.n13106 D.n13105 0.015
R22633 D.n12316 D.n12315 0.015
R22634 D.n12304 D.n12302 0.015
R22635 D.n12237 D.n12236 0.015
R22636 D.n12222 D.n12221 0.015
R22637 D.n11507 D.n11506 0.015
R22638 D.n11497 D.n11496 0.015
R22639 D.n11438 D.n11437 0.015
R22640 D.n11423 D.n11422 0.015
R22641 D.n10784 D.n10783 0.015
R22642 D.n10774 D.n10773 0.015
R22643 D.n10719 D.n10718 0.015
R22644 D.n10704 D.n10703 0.015
R22645 D.n10141 D.n10140 0.015
R22646 D.n10129 D.n10127 0.015
R22647 D.n10084 D.n10083 0.015
R22648 D.n10064 D.n10063 0.015
R22649 D.n9578 D.n9577 0.015
R22650 D.n9566 D.n9564 0.015
R22651 D.n9515 D.n9514 0.015
R22652 D.n9500 D.n9499 0.015
R22653 D.n9089 D.n9088 0.015
R22654 D.n9079 D.n9078 0.015
R22655 D.n9036 D.n9035 0.015
R22656 D.n9021 D.n9020 0.015
R22657 D.n8686 D.n8685 0.015
R22658 D.n8674 D.n8672 0.015
R22659 D.n8641 D.n8640 0.015
R22660 D.n8621 D.n8620 0.015
R22661 D.n8363 D.n8362 0.015
R22662 D.n8351 D.n8349 0.015
R22663 D.n8312 D.n8311 0.015
R22664 D.n8297 D.n8296 0.015
R22665 D.n8114 D.n8113 0.015
R22666 D.n8104 D.n8103 0.015
R22667 D.n8073 D.n8072 0.015
R22668 D.n8058 D.n8057 0.015
R22669 D.n7937 D.n7935 0.015
R22670 D.n502 D.n13 0.014
R22671 D.n42 D.n41 0.013
R22672 D.n24 D.n23 0.013
R22673 D.n547 D.n546 0.013
R22674 D.n561 D.n560 0.013
R22675 D.n575 D.n574 0.013
R22676 D.n589 D.n588 0.013
R22677 D.n603 D.n602 0.013
R22678 D.n617 D.n616 0.013
R22679 D.n631 D.n630 0.013
R22680 D.n645 D.n644 0.013
R22681 D.n659 D.n658 0.013
R22682 D.n673 D.n672 0.013
R22683 D.n687 D.n686 0.013
R22684 D.n701 D.n700 0.013
R22685 D.n715 D.n714 0.013
R22686 D.n729 D.n728 0.013
R22687 D.n743 D.n742 0.013
R22688 D.n757 D.n756 0.013
R22689 D.n771 D.n770 0.013
R22690 D.n785 D.n784 0.013
R22691 D.n799 D.n798 0.013
R22692 D.n813 D.n812 0.013
R22693 D.n827 D.n826 0.013
R22694 D.n841 D.n840 0.013
R22695 D.n855 D.n854 0.013
R22696 D.n869 D.n868 0.013
R22697 D.n883 D.n882 0.013
R22698 D.n897 D.n896 0.013
R22699 D.n911 D.n910 0.013
R22700 D.n925 D.n924 0.013
R22701 D.n939 D.n938 0.013
R22702 D.n953 D.n952 0.013
R22703 D.n967 D.n966 0.013
R22704 D.n981 D.n980 0.013
R22705 D.n995 D.n994 0.013
R22706 D.n1009 D.n1008 0.013
R22707 D.n1023 D.n1022 0.013
R22708 D.n1037 D.n1036 0.013
R22709 D.n1051 D.n1050 0.013
R22710 D.n1065 D.n1064 0.013
R22711 D.n1079 D.n1078 0.013
R22712 D.n1093 D.n1092 0.013
R22713 D.n1107 D.n1106 0.013
R22714 D.n1121 D.n1120 0.013
R22715 D.n1135 D.n1134 0.013
R22716 D.n1140 D.n1139 0.013
R22717 D.n1174 D.n1173 0.013
R22718 D.n1188 D.n1187 0.013
R22719 D.n1202 D.n1201 0.013
R22720 D.n1216 D.n1215 0.013
R22721 D.n1230 D.n1229 0.013
R22722 D.n1244 D.n1243 0.013
R22723 D.n1258 D.n1257 0.013
R22724 D.n1272 D.n1271 0.013
R22725 D.n1286 D.n1285 0.013
R22726 D.n1300 D.n1299 0.013
R22727 D.n1314 D.n1313 0.013
R22728 D.n1328 D.n1327 0.013
R22729 D.n1342 D.n1341 0.013
R22730 D.n1356 D.n1355 0.013
R22731 D.n1370 D.n1369 0.013
R22732 D.n1384 D.n1383 0.013
R22733 D.n1398 D.n1397 0.013
R22734 D.n1412 D.n1411 0.013
R22735 D.n1426 D.n1425 0.013
R22736 D.n1440 D.n1439 0.013
R22737 D.n1454 D.n1453 0.013
R22738 D.n1468 D.n1467 0.013
R22739 D.n1482 D.n1481 0.013
R22740 D.n1496 D.n1495 0.013
R22741 D.n1510 D.n1509 0.013
R22742 D.n1524 D.n1523 0.013
R22743 D.n1538 D.n1537 0.013
R22744 D.n1552 D.n1551 0.013
R22745 D.n1566 D.n1565 0.013
R22746 D.n1580 D.n1579 0.013
R22747 D.n1594 D.n1593 0.013
R22748 D.n1608 D.n1607 0.013
R22749 D.n1622 D.n1621 0.013
R22750 D.n1636 D.n1635 0.013
R22751 D.n1650 D.n1649 0.013
R22752 D.n1664 D.n1663 0.013
R22753 D.n1678 D.n1677 0.013
R22754 D.n1692 D.n1691 0.013
R22755 D.n1706 D.n1705 0.013
R22756 D.n1720 D.n1719 0.013
R22757 D.n1734 D.n1733 0.013
R22758 D.n1739 D.n1738 0.013
R22759 D.n1773 D.n1772 0.013
R22760 D.n1787 D.n1786 0.013
R22761 D.n1801 D.n1800 0.013
R22762 D.n1815 D.n1814 0.013
R22763 D.n1829 D.n1828 0.013
R22764 D.n1843 D.n1842 0.013
R22765 D.n1857 D.n1856 0.013
R22766 D.n1871 D.n1870 0.013
R22767 D.n1885 D.n1884 0.013
R22768 D.n1899 D.n1898 0.013
R22769 D.n1913 D.n1912 0.013
R22770 D.n1927 D.n1926 0.013
R22771 D.n1941 D.n1940 0.013
R22772 D.n1955 D.n1954 0.013
R22773 D.n1969 D.n1968 0.013
R22774 D.n1983 D.n1982 0.013
R22775 D.n1997 D.n1996 0.013
R22776 D.n2011 D.n2010 0.013
R22777 D.n2025 D.n2024 0.013
R22778 D.n2039 D.n2038 0.013
R22779 D.n2053 D.n2052 0.013
R22780 D.n2067 D.n2066 0.013
R22781 D.n2081 D.n2080 0.013
R22782 D.n2095 D.n2094 0.013
R22783 D.n2109 D.n2108 0.013
R22784 D.n2123 D.n2122 0.013
R22785 D.n2137 D.n2136 0.013
R22786 D.n2151 D.n2150 0.013
R22787 D.n2165 D.n2164 0.013
R22788 D.n2179 D.n2178 0.013
R22789 D.n2193 D.n2192 0.013
R22790 D.n2207 D.n2206 0.013
R22791 D.n2221 D.n2220 0.013
R22792 D.n2235 D.n2234 0.013
R22793 D.n2249 D.n2248 0.013
R22794 D.n2263 D.n2262 0.013
R22795 D.n2277 D.n2276 0.013
R22796 D.n2291 D.n2290 0.013
R22797 D.n2305 D.n2304 0.013
R22798 D.n2310 D.n2309 0.013
R22799 D.n2344 D.n2343 0.013
R22800 D.n2358 D.n2357 0.013
R22801 D.n2372 D.n2371 0.013
R22802 D.n2386 D.n2385 0.013
R22803 D.n2400 D.n2399 0.013
R22804 D.n2414 D.n2413 0.013
R22805 D.n2428 D.n2427 0.013
R22806 D.n2442 D.n2441 0.013
R22807 D.n2456 D.n2455 0.013
R22808 D.n2470 D.n2469 0.013
R22809 D.n2484 D.n2483 0.013
R22810 D.n2498 D.n2497 0.013
R22811 D.n2512 D.n2511 0.013
R22812 D.n2526 D.n2525 0.013
R22813 D.n2540 D.n2539 0.013
R22814 D.n2554 D.n2553 0.013
R22815 D.n2568 D.n2567 0.013
R22816 D.n2582 D.n2581 0.013
R22817 D.n2596 D.n2595 0.013
R22818 D.n2610 D.n2609 0.013
R22819 D.n2624 D.n2623 0.013
R22820 D.n2638 D.n2637 0.013
R22821 D.n2652 D.n2651 0.013
R22822 D.n2666 D.n2665 0.013
R22823 D.n2680 D.n2679 0.013
R22824 D.n2694 D.n2693 0.013
R22825 D.n2708 D.n2707 0.013
R22826 D.n2722 D.n2721 0.013
R22827 D.n2736 D.n2735 0.013
R22828 D.n2750 D.n2749 0.013
R22829 D.n2764 D.n2763 0.013
R22830 D.n2778 D.n2777 0.013
R22831 D.n2792 D.n2791 0.013
R22832 D.n2806 D.n2805 0.013
R22833 D.n2820 D.n2819 0.013
R22834 D.n2834 D.n2833 0.013
R22835 D.n2848 D.n2847 0.013
R22836 D.n2853 D.n2852 0.013
R22837 D.n2887 D.n2886 0.013
R22838 D.n2901 D.n2900 0.013
R22839 D.n2915 D.n2914 0.013
R22840 D.n2929 D.n2928 0.013
R22841 D.n2943 D.n2942 0.013
R22842 D.n2957 D.n2956 0.013
R22843 D.n2971 D.n2970 0.013
R22844 D.n2985 D.n2984 0.013
R22845 D.n2999 D.n2998 0.013
R22846 D.n3013 D.n3012 0.013
R22847 D.n3027 D.n3026 0.013
R22848 D.n3041 D.n3040 0.013
R22849 D.n3055 D.n3054 0.013
R22850 D.n3069 D.n3068 0.013
R22851 D.n3083 D.n3082 0.013
R22852 D.n3097 D.n3096 0.013
R22853 D.n3111 D.n3110 0.013
R22854 D.n3125 D.n3124 0.013
R22855 D.n3139 D.n3138 0.013
R22856 D.n3153 D.n3152 0.013
R22857 D.n3167 D.n3166 0.013
R22858 D.n3181 D.n3180 0.013
R22859 D.n3195 D.n3194 0.013
R22860 D.n3209 D.n3208 0.013
R22861 D.n3223 D.n3222 0.013
R22862 D.n3237 D.n3236 0.013
R22863 D.n3251 D.n3250 0.013
R22864 D.n3265 D.n3264 0.013
R22865 D.n3279 D.n3278 0.013
R22866 D.n3293 D.n3292 0.013
R22867 D.n3307 D.n3306 0.013
R22868 D.n3321 D.n3320 0.013
R22869 D.n3335 D.n3334 0.013
R22870 D.n3349 D.n3348 0.013
R22871 D.n3363 D.n3362 0.013
R22872 D.n3368 D.n3367 0.013
R22873 D.n3403 D.n3402 0.013
R22874 D.n3417 D.n3416 0.013
R22875 D.n3431 D.n3430 0.013
R22876 D.n3445 D.n3444 0.013
R22877 D.n3459 D.n3458 0.013
R22878 D.n3473 D.n3472 0.013
R22879 D.n3487 D.n3486 0.013
R22880 D.n3501 D.n3500 0.013
R22881 D.n3515 D.n3514 0.013
R22882 D.n3529 D.n3528 0.013
R22883 D.n3543 D.n3542 0.013
R22884 D.n3557 D.n3556 0.013
R22885 D.n3571 D.n3570 0.013
R22886 D.n3585 D.n3584 0.013
R22887 D.n3599 D.n3598 0.013
R22888 D.n3613 D.n3612 0.013
R22889 D.n3627 D.n3626 0.013
R22890 D.n3641 D.n3640 0.013
R22891 D.n3655 D.n3654 0.013
R22892 D.n3669 D.n3668 0.013
R22893 D.n3683 D.n3682 0.013
R22894 D.n3697 D.n3696 0.013
R22895 D.n3711 D.n3710 0.013
R22896 D.n3725 D.n3724 0.013
R22897 D.n3739 D.n3738 0.013
R22898 D.n3753 D.n3752 0.013
R22899 D.n3767 D.n3766 0.013
R22900 D.n3781 D.n3780 0.013
R22901 D.n3795 D.n3794 0.013
R22902 D.n3809 D.n3808 0.013
R22903 D.n3823 D.n3822 0.013
R22904 D.n3837 D.n3836 0.013
R22905 D.n3851 D.n3850 0.013
R22906 D.n3856 D.n3855 0.013
R22907 D.n3891 D.n3890 0.013
R22908 D.n3905 D.n3904 0.013
R22909 D.n3919 D.n3918 0.013
R22910 D.n3933 D.n3932 0.013
R22911 D.n3947 D.n3946 0.013
R22912 D.n3961 D.n3960 0.013
R22913 D.n3975 D.n3974 0.013
R22914 D.n3989 D.n3988 0.013
R22915 D.n4003 D.n4002 0.013
R22916 D.n4017 D.n4016 0.013
R22917 D.n4031 D.n4030 0.013
R22918 D.n4045 D.n4044 0.013
R22919 D.n4059 D.n4058 0.013
R22920 D.n4073 D.n4072 0.013
R22921 D.n4087 D.n4086 0.013
R22922 D.n4101 D.n4100 0.013
R22923 D.n4115 D.n4114 0.013
R22924 D.n4129 D.n4128 0.013
R22925 D.n4143 D.n4142 0.013
R22926 D.n4157 D.n4156 0.013
R22927 D.n4171 D.n4170 0.013
R22928 D.n4185 D.n4184 0.013
R22929 D.n4199 D.n4198 0.013
R22930 D.n4213 D.n4212 0.013
R22931 D.n4227 D.n4226 0.013
R22932 D.n4241 D.n4240 0.013
R22933 D.n4255 D.n4254 0.013
R22934 D.n4269 D.n4268 0.013
R22935 D.n4283 D.n4282 0.013
R22936 D.n4297 D.n4296 0.013
R22937 D.n4311 D.n4310 0.013
R22938 D.n4316 D.n4315 0.013
R22939 D.n4351 D.n4350 0.013
R22940 D.n4365 D.n4364 0.013
R22941 D.n4379 D.n4378 0.013
R22942 D.n4393 D.n4392 0.013
R22943 D.n4407 D.n4406 0.013
R22944 D.n4421 D.n4420 0.013
R22945 D.n4435 D.n4434 0.013
R22946 D.n4449 D.n4448 0.013
R22947 D.n4463 D.n4462 0.013
R22948 D.n4477 D.n4476 0.013
R22949 D.n4491 D.n4490 0.013
R22950 D.n4505 D.n4504 0.013
R22951 D.n4519 D.n4518 0.013
R22952 D.n4533 D.n4532 0.013
R22953 D.n4547 D.n4546 0.013
R22954 D.n4561 D.n4560 0.013
R22955 D.n4575 D.n4574 0.013
R22956 D.n4589 D.n4588 0.013
R22957 D.n4603 D.n4602 0.013
R22958 D.n4617 D.n4616 0.013
R22959 D.n4631 D.n4630 0.013
R22960 D.n4645 D.n4644 0.013
R22961 D.n4659 D.n4658 0.013
R22962 D.n4673 D.n4672 0.013
R22963 D.n4687 D.n4686 0.013
R22964 D.n4701 D.n4700 0.013
R22965 D.n4715 D.n4714 0.013
R22966 D.n4729 D.n4728 0.013
R22967 D.n4743 D.n4742 0.013
R22968 D.n4748 D.n4747 0.013
R22969 D.n4783 D.n4782 0.013
R22970 D.n4797 D.n4796 0.013
R22971 D.n4811 D.n4810 0.013
R22972 D.n4825 D.n4824 0.013
R22973 D.n4839 D.n4838 0.013
R22974 D.n4853 D.n4852 0.013
R22975 D.n4867 D.n4866 0.013
R22976 D.n4881 D.n4880 0.013
R22977 D.n4895 D.n4894 0.013
R22978 D.n4909 D.n4908 0.013
R22979 D.n4923 D.n4922 0.013
R22980 D.n4937 D.n4936 0.013
R22981 D.n4951 D.n4950 0.013
R22982 D.n4965 D.n4964 0.013
R22983 D.n4979 D.n4978 0.013
R22984 D.n4993 D.n4992 0.013
R22985 D.n5007 D.n5006 0.013
R22986 D.n5021 D.n5020 0.013
R22987 D.n5035 D.n5034 0.013
R22988 D.n5049 D.n5048 0.013
R22989 D.n5063 D.n5062 0.013
R22990 D.n5077 D.n5076 0.013
R22991 D.n5091 D.n5090 0.013
R22992 D.n5105 D.n5104 0.013
R22993 D.n5119 D.n5118 0.013
R22994 D.n5133 D.n5132 0.013
R22995 D.n5147 D.n5146 0.013
R22996 D.n5152 D.n5151 0.013
R22997 D.n5187 D.n5186 0.013
R22998 D.n5201 D.n5200 0.013
R22999 D.n5215 D.n5214 0.013
R23000 D.n5229 D.n5228 0.013
R23001 D.n5243 D.n5242 0.013
R23002 D.n5257 D.n5256 0.013
R23003 D.n5271 D.n5270 0.013
R23004 D.n5285 D.n5284 0.013
R23005 D.n5299 D.n5298 0.013
R23006 D.n5313 D.n5312 0.013
R23007 D.n5327 D.n5326 0.013
R23008 D.n5341 D.n5340 0.013
R23009 D.n5355 D.n5354 0.013
R23010 D.n5369 D.n5368 0.013
R23011 D.n5383 D.n5382 0.013
R23012 D.n5397 D.n5396 0.013
R23013 D.n5411 D.n5410 0.013
R23014 D.n5425 D.n5424 0.013
R23015 D.n5439 D.n5438 0.013
R23016 D.n5453 D.n5452 0.013
R23017 D.n5467 D.n5466 0.013
R23018 D.n5481 D.n5480 0.013
R23019 D.n5495 D.n5494 0.013
R23020 D.n5509 D.n5508 0.013
R23021 D.n5523 D.n5522 0.013
R23022 D.n5528 D.n5527 0.013
R23023 D.n5563 D.n5562 0.013
R23024 D.n5577 D.n5576 0.013
R23025 D.n5591 D.n5590 0.013
R23026 D.n5605 D.n5604 0.013
R23027 D.n5619 D.n5618 0.013
R23028 D.n5633 D.n5632 0.013
R23029 D.n5647 D.n5646 0.013
R23030 D.n5661 D.n5660 0.013
R23031 D.n5675 D.n5674 0.013
R23032 D.n5689 D.n5688 0.013
R23033 D.n5703 D.n5702 0.013
R23034 D.n5717 D.n5716 0.013
R23035 D.n5731 D.n5730 0.013
R23036 D.n5745 D.n5744 0.013
R23037 D.n5759 D.n5758 0.013
R23038 D.n5773 D.n5772 0.013
R23039 D.n5787 D.n5786 0.013
R23040 D.n5801 D.n5800 0.013
R23041 D.n5815 D.n5814 0.013
R23042 D.n5829 D.n5828 0.013
R23043 D.n5843 D.n5842 0.013
R23044 D.n5857 D.n5856 0.013
R23045 D.n5871 D.n5870 0.013
R23046 D.n5876 D.n5875 0.013
R23047 D.n5911 D.n5910 0.013
R23048 D.n5925 D.n5924 0.013
R23049 D.n5939 D.n5938 0.013
R23050 D.n5953 D.n5952 0.013
R23051 D.n5967 D.n5966 0.013
R23052 D.n5981 D.n5980 0.013
R23053 D.n5995 D.n5994 0.013
R23054 D.n6009 D.n6008 0.013
R23055 D.n6023 D.n6022 0.013
R23056 D.n6037 D.n6036 0.013
R23057 D.n6051 D.n6050 0.013
R23058 D.n6065 D.n6064 0.013
R23059 D.n6079 D.n6078 0.013
R23060 D.n6093 D.n6092 0.013
R23061 D.n6107 D.n6106 0.013
R23062 D.n6121 D.n6120 0.013
R23063 D.n6135 D.n6134 0.013
R23064 D.n6149 D.n6148 0.013
R23065 D.n6163 D.n6162 0.013
R23066 D.n6177 D.n6176 0.013
R23067 D.n6191 D.n6190 0.013
R23068 D.n6196 D.n6195 0.013
R23069 D.n6231 D.n6230 0.013
R23070 D.n6245 D.n6244 0.013
R23071 D.n6259 D.n6258 0.013
R23072 D.n6273 D.n6272 0.013
R23073 D.n6287 D.n6286 0.013
R23074 D.n6301 D.n6300 0.013
R23075 D.n6315 D.n6314 0.013
R23076 D.n6329 D.n6328 0.013
R23077 D.n6343 D.n6342 0.013
R23078 D.n6357 D.n6356 0.013
R23079 D.n6371 D.n6370 0.013
R23080 D.n6385 D.n6384 0.013
R23081 D.n6399 D.n6398 0.013
R23082 D.n6413 D.n6412 0.013
R23083 D.n6427 D.n6426 0.013
R23084 D.n6441 D.n6440 0.013
R23085 D.n6455 D.n6454 0.013
R23086 D.n6469 D.n6468 0.013
R23087 D.n6483 D.n6482 0.013
R23088 D.n6488 D.n6487 0.013
R23089 D.n6523 D.n6522 0.013
R23090 D.n6537 D.n6536 0.013
R23091 D.n6551 D.n6550 0.013
R23092 D.n6565 D.n6564 0.013
R23093 D.n6579 D.n6578 0.013
R23094 D.n6593 D.n6592 0.013
R23095 D.n6607 D.n6606 0.013
R23096 D.n6621 D.n6620 0.013
R23097 D.n6635 D.n6634 0.013
R23098 D.n6649 D.n6648 0.013
R23099 D.n6663 D.n6662 0.013
R23100 D.n6677 D.n6676 0.013
R23101 D.n6691 D.n6690 0.013
R23102 D.n6705 D.n6704 0.013
R23103 D.n6719 D.n6718 0.013
R23104 D.n6733 D.n6732 0.013
R23105 D.n6747 D.n6746 0.013
R23106 D.n6752 D.n6751 0.013
R23107 D.n6787 D.n6786 0.013
R23108 D.n6801 D.n6800 0.013
R23109 D.n6815 D.n6814 0.013
R23110 D.n6829 D.n6828 0.013
R23111 D.n6843 D.n6842 0.013
R23112 D.n6857 D.n6856 0.013
R23113 D.n6871 D.n6870 0.013
R23114 D.n6885 D.n6884 0.013
R23115 D.n6899 D.n6898 0.013
R23116 D.n6913 D.n6912 0.013
R23117 D.n6927 D.n6926 0.013
R23118 D.n6941 D.n6940 0.013
R23119 D.n6955 D.n6954 0.013
R23120 D.n6969 D.n6968 0.013
R23121 D.n6983 D.n6982 0.013
R23122 D.n6988 D.n6987 0.013
R23123 D.n7023 D.n7022 0.013
R23124 D.n7037 D.n7036 0.013
R23125 D.n7051 D.n7050 0.013
R23126 D.n7065 D.n7064 0.013
R23127 D.n7079 D.n7078 0.013
R23128 D.n7093 D.n7092 0.013
R23129 D.n7107 D.n7106 0.013
R23130 D.n7121 D.n7120 0.013
R23131 D.n7135 D.n7134 0.013
R23132 D.n7149 D.n7148 0.013
R23133 D.n7163 D.n7162 0.013
R23134 D.n7177 D.n7176 0.013
R23135 D.n7191 D.n7190 0.013
R23136 D.n7196 D.n7195 0.013
R23137 D.n7231 D.n7230 0.013
R23138 D.n7245 D.n7244 0.013
R23139 D.n7259 D.n7258 0.013
R23140 D.n7273 D.n7272 0.013
R23141 D.n7287 D.n7286 0.013
R23142 D.n7301 D.n7300 0.013
R23143 D.n7315 D.n7314 0.013
R23144 D.n7329 D.n7328 0.013
R23145 D.n7343 D.n7342 0.013
R23146 D.n7357 D.n7356 0.013
R23147 D.n7371 D.n7370 0.013
R23148 D.n7376 D.n7375 0.013
R23149 D.n7411 D.n7410 0.013
R23150 D.n7425 D.n7424 0.013
R23151 D.n7439 D.n7438 0.013
R23152 D.n7453 D.n7452 0.013
R23153 D.n7467 D.n7466 0.013
R23154 D.n7481 D.n7480 0.013
R23155 D.n7495 D.n7494 0.013
R23156 D.n7509 D.n7508 0.013
R23157 D.n7523 D.n7522 0.013
R23158 D.n7528 D.n7527 0.013
R23159 D.n7563 D.n7562 0.013
R23160 D.n7577 D.n7576 0.013
R23161 D.n7591 D.n7590 0.013
R23162 D.n7605 D.n7604 0.013
R23163 D.n7619 D.n7618 0.013
R23164 D.n7633 D.n7632 0.013
R23165 D.n7647 D.n7646 0.013
R23166 D.n7652 D.n7651 0.013
R23167 D.n7687 D.n7686 0.013
R23168 D.n7701 D.n7700 0.013
R23169 D.n7715 D.n7714 0.013
R23170 D.n7729 D.n7728 0.013
R23171 D.n7743 D.n7742 0.013
R23172 D.n7748 D.n7747 0.013
R23173 D.n7782 D.n7781 0.013
R23174 D.n7796 D.n7795 0.013
R23175 D.n7812 D.n7811 0.013
R23176 D.n13658 D.n13657 0.012
R23177 D.n13623 D.n13622 0.012
R23178 D.n12735 D.n12734 0.012
R23179 D.n12700 D.n12699 0.012
R23180 D.n11886 D.n11885 0.012
R23181 D.n11851 D.n11850 0.012
R23182 D.n11123 D.n11122 0.012
R23183 D.n11088 D.n11087 0.012
R23184 D.n10440 D.n10439 0.012
R23185 D.n10405 D.n10404 0.012
R23186 D.n9837 D.n9836 0.012
R23187 D.n9802 D.n9801 0.012
R23188 D.n9308 D.n9307 0.012
R23189 D.n9273 D.n9272 0.012
R23190 D.n8865 D.n8864 0.012
R23191 D.n8830 D.n8829 0.012
R23192 D.n8502 D.n8501 0.012
R23193 D.n8467 D.n8466 0.012
R23194 D.n8213 D.n8212 0.012
R23195 D.n8178 D.n8177 0.012
R23196 D.n8010 D.n8009 0.012
R23197 D.n7973 D.n7972 0.012
R23198 D.n453 D.n452 0.011
R23199 D.n7843 D.n7842 0.011
R23200 D.n13689 D.n13688 0.011
R23201 D.n13707 D.n13706 0.011
R23202 D.n13725 D.n13724 0.011
R23203 D.n13743 D.n13742 0.011
R23204 D.n13761 D.n13760 0.011
R23205 D.n13779 D.n13778 0.011
R23206 D.n13797 D.n13796 0.011
R23207 D.n13815 D.n13814 0.011
R23208 D.n13833 D.n13832 0.011
R23209 D.n13851 D.n13850 0.011
R23210 D.n13869 D.n13868 0.011
R23211 D.n13887 D.n13886 0.011
R23212 D.n13905 D.n13904 0.011
R23213 D.n13923 D.n13922 0.011
R23214 D.n13941 D.n13940 0.011
R23215 D.n13959 D.n13958 0.011
R23216 D.n13977 D.n13976 0.011
R23217 D.n13995 D.n13994 0.011
R23218 D.n14013 D.n14012 0.011
R23219 D.n14031 D.n14030 0.011
R23220 D.n14049 D.n14048 0.011
R23221 D.n14067 D.n14066 0.011
R23222 D.n13613 D.n13612 0.011
R23223 D.n13593 D.n13592 0.011
R23224 D.n13573 D.n13572 0.011
R23225 D.n13553 D.n13552 0.011
R23226 D.n13533 D.n13532 0.011
R23227 D.n13513 D.n13512 0.011
R23228 D.n13493 D.n13492 0.011
R23229 D.n13473 D.n13472 0.011
R23230 D.n13453 D.n13452 0.011
R23231 D.n13433 D.n13432 0.011
R23232 D.n13413 D.n13412 0.011
R23233 D.n13393 D.n13392 0.011
R23234 D.n13373 D.n13372 0.011
R23235 D.n13353 D.n13352 0.011
R23236 D.n13333 D.n13332 0.011
R23237 D.n13313 D.n13312 0.011
R23238 D.n13293 D.n13292 0.011
R23239 D.n13273 D.n13272 0.011
R23240 D.n13253 D.n13252 0.011
R23241 D.n13233 D.n13232 0.011
R23242 D.n13213 D.n13212 0.011
R23243 D.n12762 D.n12761 0.011
R23244 D.n12780 D.n12779 0.011
R23245 D.n12798 D.n12797 0.011
R23246 D.n12816 D.n12815 0.011
R23247 D.n12834 D.n12833 0.011
R23248 D.n12852 D.n12851 0.011
R23249 D.n12870 D.n12869 0.011
R23250 D.n12888 D.n12887 0.011
R23251 D.n12906 D.n12905 0.011
R23252 D.n12924 D.n12923 0.011
R23253 D.n12942 D.n12941 0.011
R23254 D.n12960 D.n12959 0.011
R23255 D.n12978 D.n12977 0.011
R23256 D.n12996 D.n12995 0.011
R23257 D.n13014 D.n13013 0.011
R23258 D.n13032 D.n13031 0.011
R23259 D.n13050 D.n13049 0.011
R23260 D.n13068 D.n13067 0.011
R23261 D.n13086 D.n13085 0.011
R23262 D.n13104 D.n13103 0.011
R23263 D.n12690 D.n12689 0.011
R23264 D.n12670 D.n12669 0.011
R23265 D.n12650 D.n12649 0.011
R23266 D.n12630 D.n12629 0.011
R23267 D.n12610 D.n12609 0.011
R23268 D.n12590 D.n12589 0.011
R23269 D.n12570 D.n12569 0.011
R23270 D.n12550 D.n12549 0.011
R23271 D.n12530 D.n12529 0.011
R23272 D.n12510 D.n12509 0.011
R23273 D.n12490 D.n12489 0.011
R23274 D.n12470 D.n12469 0.011
R23275 D.n12450 D.n12449 0.011
R23276 D.n12430 D.n12429 0.011
R23277 D.n12410 D.n12409 0.011
R23278 D.n12390 D.n12389 0.011
R23279 D.n12370 D.n12369 0.011
R23280 D.n12350 D.n12349 0.011
R23281 D.n12330 D.n12329 0.011
R23282 D.n11913 D.n11912 0.011
R23283 D.n11931 D.n11930 0.011
R23284 D.n11949 D.n11948 0.011
R23285 D.n11967 D.n11966 0.011
R23286 D.n11985 D.n11984 0.011
R23287 D.n12003 D.n12002 0.011
R23288 D.n12021 D.n12020 0.011
R23289 D.n12039 D.n12038 0.011
R23290 D.n12057 D.n12056 0.011
R23291 D.n12075 D.n12074 0.011
R23292 D.n12093 D.n12092 0.011
R23293 D.n12111 D.n12110 0.011
R23294 D.n12129 D.n12128 0.011
R23295 D.n12147 D.n12146 0.011
R23296 D.n12165 D.n12164 0.011
R23297 D.n12183 D.n12182 0.011
R23298 D.n12201 D.n12200 0.011
R23299 D.n12219 D.n12218 0.011
R23300 D.n11841 D.n11840 0.011
R23301 D.n11821 D.n11820 0.011
R23302 D.n11801 D.n11800 0.011
R23303 D.n11781 D.n11780 0.011
R23304 D.n11761 D.n11760 0.011
R23305 D.n11741 D.n11740 0.011
R23306 D.n11721 D.n11720 0.011
R23307 D.n11701 D.n11700 0.011
R23308 D.n11681 D.n11680 0.011
R23309 D.n11661 D.n11660 0.011
R23310 D.n11641 D.n11640 0.011
R23311 D.n11621 D.n11620 0.011
R23312 D.n11601 D.n11600 0.011
R23313 D.n11581 D.n11580 0.011
R23314 D.n11561 D.n11560 0.011
R23315 D.n11541 D.n11540 0.011
R23316 D.n11521 D.n11520 0.011
R23317 D.n11150 D.n11149 0.011
R23318 D.n11168 D.n11167 0.011
R23319 D.n11186 D.n11185 0.011
R23320 D.n11204 D.n11203 0.011
R23321 D.n11222 D.n11221 0.011
R23322 D.n11240 D.n11239 0.011
R23323 D.n11258 D.n11257 0.011
R23324 D.n11276 D.n11275 0.011
R23325 D.n11294 D.n11293 0.011
R23326 D.n11312 D.n11311 0.011
R23327 D.n11330 D.n11329 0.011
R23328 D.n11348 D.n11347 0.011
R23329 D.n11366 D.n11365 0.011
R23330 D.n11384 D.n11383 0.011
R23331 D.n11402 D.n11401 0.011
R23332 D.n11420 D.n11419 0.011
R23333 D.n11078 D.n11077 0.011
R23334 D.n11058 D.n11057 0.011
R23335 D.n11038 D.n11037 0.011
R23336 D.n11018 D.n11017 0.011
R23337 D.n10998 D.n10997 0.011
R23338 D.n10978 D.n10977 0.011
R23339 D.n10958 D.n10957 0.011
R23340 D.n10938 D.n10937 0.011
R23341 D.n10918 D.n10917 0.011
R23342 D.n10898 D.n10897 0.011
R23343 D.n10878 D.n10877 0.011
R23344 D.n10858 D.n10857 0.011
R23345 D.n10838 D.n10837 0.011
R23346 D.n10818 D.n10817 0.011
R23347 D.n10798 D.n10797 0.011
R23348 D.n10467 D.n10466 0.011
R23349 D.n10485 D.n10484 0.011
R23350 D.n10503 D.n10502 0.011
R23351 D.n10521 D.n10520 0.011
R23352 D.n10539 D.n10538 0.011
R23353 D.n10557 D.n10556 0.011
R23354 D.n10575 D.n10574 0.011
R23355 D.n10593 D.n10592 0.011
R23356 D.n10611 D.n10610 0.011
R23357 D.n10629 D.n10628 0.011
R23358 D.n10647 D.n10646 0.011
R23359 D.n10665 D.n10664 0.011
R23360 D.n10683 D.n10682 0.011
R23361 D.n10701 D.n10700 0.011
R23362 D.n10395 D.n10394 0.011
R23363 D.n10375 D.n10374 0.011
R23364 D.n10355 D.n10354 0.011
R23365 D.n10335 D.n10334 0.011
R23366 D.n10315 D.n10314 0.011
R23367 D.n10295 D.n10294 0.011
R23368 D.n10275 D.n10274 0.011
R23369 D.n10255 D.n10254 0.011
R23370 D.n10235 D.n10234 0.011
R23371 D.n10215 D.n10214 0.011
R23372 D.n10195 D.n10194 0.011
R23373 D.n10175 D.n10174 0.011
R23374 D.n10155 D.n10154 0.011
R23375 D.n9864 D.n9863 0.011
R23376 D.n9882 D.n9881 0.011
R23377 D.n9900 D.n9899 0.011
R23378 D.n9918 D.n9917 0.011
R23379 D.n9936 D.n9935 0.011
R23380 D.n9954 D.n9953 0.011
R23381 D.n9972 D.n9971 0.011
R23382 D.n9990 D.n9989 0.011
R23383 D.n10008 D.n10007 0.011
R23384 D.n10026 D.n10025 0.011
R23385 D.n10044 D.n10043 0.011
R23386 D.n10062 D.n10061 0.011
R23387 D.n9792 D.n9791 0.011
R23388 D.n9772 D.n9771 0.011
R23389 D.n9752 D.n9751 0.011
R23390 D.n9732 D.n9731 0.011
R23391 D.n9712 D.n9711 0.011
R23392 D.n9692 D.n9691 0.011
R23393 D.n9672 D.n9671 0.011
R23394 D.n9652 D.n9651 0.011
R23395 D.n9632 D.n9631 0.011
R23396 D.n9612 D.n9611 0.011
R23397 D.n9592 D.n9591 0.011
R23398 D.n9335 D.n9334 0.011
R23399 D.n9353 D.n9352 0.011
R23400 D.n9371 D.n9370 0.011
R23401 D.n9389 D.n9388 0.011
R23402 D.n9407 D.n9406 0.011
R23403 D.n9425 D.n9424 0.011
R23404 D.n9443 D.n9442 0.011
R23405 D.n9461 D.n9460 0.011
R23406 D.n9479 D.n9478 0.011
R23407 D.n9497 D.n9496 0.011
R23408 D.n9263 D.n9262 0.011
R23409 D.n9243 D.n9242 0.011
R23410 D.n9223 D.n9222 0.011
R23411 D.n9203 D.n9202 0.011
R23412 D.n9183 D.n9182 0.011
R23413 D.n9163 D.n9162 0.011
R23414 D.n9143 D.n9142 0.011
R23415 D.n9123 D.n9122 0.011
R23416 D.n9103 D.n9102 0.011
R23417 D.n8892 D.n8891 0.011
R23418 D.n8910 D.n8909 0.011
R23419 D.n8928 D.n8927 0.011
R23420 D.n8946 D.n8945 0.011
R23421 D.n8964 D.n8963 0.011
R23422 D.n8982 D.n8981 0.011
R23423 D.n9000 D.n8999 0.011
R23424 D.n9018 D.n9017 0.011
R23425 D.n8820 D.n8819 0.011
R23426 D.n8800 D.n8799 0.011
R23427 D.n8780 D.n8779 0.011
R23428 D.n8760 D.n8759 0.011
R23429 D.n8740 D.n8739 0.011
R23430 D.n8720 D.n8719 0.011
R23431 D.n8700 D.n8699 0.011
R23432 D.n8529 D.n8528 0.011
R23433 D.n8547 D.n8546 0.011
R23434 D.n8565 D.n8564 0.011
R23435 D.n8583 D.n8582 0.011
R23436 D.n8601 D.n8600 0.011
R23437 D.n8619 D.n8618 0.011
R23438 D.n8457 D.n8456 0.011
R23439 D.n8437 D.n8436 0.011
R23440 D.n8417 D.n8416 0.011
R23441 D.n8397 D.n8396 0.011
R23442 D.n8377 D.n8376 0.011
R23443 D.n8240 D.n8239 0.011
R23444 D.n8258 D.n8257 0.011
R23445 D.n8276 D.n8275 0.011
R23446 D.n8294 D.n8293 0.011
R23447 D.n8168 D.n8167 0.011
R23448 D.n8148 D.n8147 0.011
R23449 D.n8128 D.n8127 0.011
R23450 D.n8037 D.n8036 0.011
R23451 D.n8055 D.n8054 0.011
R23452 D.n7963 D.n7962 0.011
R23453 D.n444 D.n443 0.011
R23454 D.n435 D.n427 0.011
R23455 D.n426 D.n418 0.011
R23456 D.n417 D.n409 0.011
R23457 D.n408 D.n400 0.011
R23458 D.n399 D.n391 0.011
R23459 D.n390 D.n382 0.011
R23460 D.n381 D.n373 0.011
R23461 D.n372 D.n364 0.011
R23462 D.n363 D.n355 0.011
R23463 D.n354 D.n346 0.011
R23464 D.n345 D.n337 0.011
R23465 D.n336 D.n328 0.011
R23466 D.n327 D.n319 0.011
R23467 D.n318 D.n310 0.011
R23468 D.n309 D.n301 0.011
R23469 D.n300 D.n292 0.011
R23470 D.n291 D.n283 0.011
R23471 D.n282 D.n274 0.011
R23472 D.n273 D.n265 0.011
R23473 D.n264 D.n256 0.011
R23474 D.n255 D.n247 0.011
R23475 D.n246 D.n238 0.011
R23476 D.n237 D.n229 0.011
R23477 D.n228 D.n220 0.011
R23478 D.n219 D.n211 0.011
R23479 D.n210 D.n202 0.011
R23480 D.n201 D.n193 0.011
R23481 D.n192 D.n184 0.011
R23482 D.n183 D.n175 0.011
R23483 D.n174 D.n166 0.011
R23484 D.n165 D.n157 0.011
R23485 D.n156 D.n148 0.011
R23486 D.n147 D.n139 0.011
R23487 D.n138 D.n130 0.011
R23488 D.n129 D.n121 0.011
R23489 D.n120 D.n112 0.011
R23490 D.n111 D.n103 0.011
R23491 D.n102 D.n94 0.011
R23492 D.n93 D.n85 0.011
R23493 D.n84 D.n76 0.011
R23494 D.n75 D.n67 0.011
R23495 D.n66 D.n58 0.011
R23496 D.n57 D.n49 0.011
R23497 D.n7833 D.n7832 0.011
R23498 D.n7816 D.n7750 0.011
R23499 D.n2 D.n1 0.01
R23500 D.n13698 D.n13690 0.01
R23501 D.n13716 D.n13708 0.01
R23502 D.n13734 D.n13726 0.01
R23503 D.n13752 D.n13744 0.01
R23504 D.n13770 D.n13762 0.01
R23505 D.n13788 D.n13780 0.01
R23506 D.n13806 D.n13798 0.01
R23507 D.n13824 D.n13816 0.01
R23508 D.n13842 D.n13834 0.01
R23509 D.n13860 D.n13852 0.01
R23510 D.n13878 D.n13870 0.01
R23511 D.n13896 D.n13888 0.01
R23512 D.n13914 D.n13906 0.01
R23513 D.n13932 D.n13924 0.01
R23514 D.n13950 D.n13942 0.01
R23515 D.n13968 D.n13960 0.01
R23516 D.n13986 D.n13978 0.01
R23517 D.n14004 D.n13996 0.01
R23518 D.n14022 D.n14014 0.01
R23519 D.n14040 D.n14032 0.01
R23520 D.n14058 D.n14050 0.01
R23521 D.n13603 D.n13602 0.01
R23522 D.n13583 D.n13582 0.01
R23523 D.n13563 D.n13562 0.01
R23524 D.n13543 D.n13542 0.01
R23525 D.n13523 D.n13522 0.01
R23526 D.n13503 D.n13502 0.01
R23527 D.n13483 D.n13482 0.01
R23528 D.n13463 D.n13462 0.01
R23529 D.n13443 D.n13442 0.01
R23530 D.n13423 D.n13422 0.01
R23531 D.n13403 D.n13402 0.01
R23532 D.n13383 D.n13382 0.01
R23533 D.n13363 D.n13362 0.01
R23534 D.n13343 D.n13342 0.01
R23535 D.n13323 D.n13322 0.01
R23536 D.n13303 D.n13302 0.01
R23537 D.n13283 D.n13282 0.01
R23538 D.n13263 D.n13262 0.01
R23539 D.n13243 D.n13242 0.01
R23540 D.n13223 D.n13222 0.01
R23541 D.n12771 D.n12763 0.01
R23542 D.n12789 D.n12781 0.01
R23543 D.n12807 D.n12799 0.01
R23544 D.n12825 D.n12817 0.01
R23545 D.n12843 D.n12835 0.01
R23546 D.n12861 D.n12853 0.01
R23547 D.n12879 D.n12871 0.01
R23548 D.n12897 D.n12889 0.01
R23549 D.n12915 D.n12907 0.01
R23550 D.n12933 D.n12925 0.01
R23551 D.n12951 D.n12943 0.01
R23552 D.n12969 D.n12961 0.01
R23553 D.n12987 D.n12979 0.01
R23554 D.n13005 D.n12997 0.01
R23555 D.n13023 D.n13015 0.01
R23556 D.n13041 D.n13033 0.01
R23557 D.n13059 D.n13051 0.01
R23558 D.n13077 D.n13069 0.01
R23559 D.n13095 D.n13087 0.01
R23560 D.n12680 D.n12679 0.01
R23561 D.n12660 D.n12659 0.01
R23562 D.n12640 D.n12639 0.01
R23563 D.n12620 D.n12619 0.01
R23564 D.n12600 D.n12599 0.01
R23565 D.n12580 D.n12579 0.01
R23566 D.n12560 D.n12559 0.01
R23567 D.n12540 D.n12539 0.01
R23568 D.n12520 D.n12519 0.01
R23569 D.n12500 D.n12499 0.01
R23570 D.n12480 D.n12479 0.01
R23571 D.n12460 D.n12459 0.01
R23572 D.n12440 D.n12439 0.01
R23573 D.n12420 D.n12419 0.01
R23574 D.n12400 D.n12399 0.01
R23575 D.n12380 D.n12379 0.01
R23576 D.n12360 D.n12359 0.01
R23577 D.n12340 D.n12339 0.01
R23578 D.n11922 D.n11914 0.01
R23579 D.n11940 D.n11932 0.01
R23580 D.n11958 D.n11950 0.01
R23581 D.n11976 D.n11968 0.01
R23582 D.n11994 D.n11986 0.01
R23583 D.n12012 D.n12004 0.01
R23584 D.n12030 D.n12022 0.01
R23585 D.n12048 D.n12040 0.01
R23586 D.n12066 D.n12058 0.01
R23587 D.n12084 D.n12076 0.01
R23588 D.n12102 D.n12094 0.01
R23589 D.n12120 D.n12112 0.01
R23590 D.n12138 D.n12130 0.01
R23591 D.n12156 D.n12148 0.01
R23592 D.n12174 D.n12166 0.01
R23593 D.n12192 D.n12184 0.01
R23594 D.n12210 D.n12202 0.01
R23595 D.n11831 D.n11830 0.01
R23596 D.n11811 D.n11810 0.01
R23597 D.n11791 D.n11790 0.01
R23598 D.n11771 D.n11770 0.01
R23599 D.n11751 D.n11750 0.01
R23600 D.n11731 D.n11730 0.01
R23601 D.n11711 D.n11710 0.01
R23602 D.n11691 D.n11690 0.01
R23603 D.n11671 D.n11670 0.01
R23604 D.n11651 D.n11650 0.01
R23605 D.n11631 D.n11630 0.01
R23606 D.n11611 D.n11610 0.01
R23607 D.n11591 D.n11590 0.01
R23608 D.n11571 D.n11570 0.01
R23609 D.n11551 D.n11550 0.01
R23610 D.n11531 D.n11530 0.01
R23611 D.n11159 D.n11151 0.01
R23612 D.n11177 D.n11169 0.01
R23613 D.n11195 D.n11187 0.01
R23614 D.n11213 D.n11205 0.01
R23615 D.n11231 D.n11223 0.01
R23616 D.n11249 D.n11241 0.01
R23617 D.n11267 D.n11259 0.01
R23618 D.n11285 D.n11277 0.01
R23619 D.n11303 D.n11295 0.01
R23620 D.n11321 D.n11313 0.01
R23621 D.n11339 D.n11331 0.01
R23622 D.n11357 D.n11349 0.01
R23623 D.n11375 D.n11367 0.01
R23624 D.n11393 D.n11385 0.01
R23625 D.n11411 D.n11403 0.01
R23626 D.n11068 D.n11067 0.01
R23627 D.n11048 D.n11047 0.01
R23628 D.n11028 D.n11027 0.01
R23629 D.n11008 D.n11007 0.01
R23630 D.n10988 D.n10987 0.01
R23631 D.n10968 D.n10967 0.01
R23632 D.n10948 D.n10947 0.01
R23633 D.n10928 D.n10927 0.01
R23634 D.n10908 D.n10907 0.01
R23635 D.n10888 D.n10887 0.01
R23636 D.n10868 D.n10867 0.01
R23637 D.n10848 D.n10847 0.01
R23638 D.n10828 D.n10827 0.01
R23639 D.n10808 D.n10807 0.01
R23640 D.n10476 D.n10468 0.01
R23641 D.n10494 D.n10486 0.01
R23642 D.n10512 D.n10504 0.01
R23643 D.n10530 D.n10522 0.01
R23644 D.n10548 D.n10540 0.01
R23645 D.n10566 D.n10558 0.01
R23646 D.n10584 D.n10576 0.01
R23647 D.n10602 D.n10594 0.01
R23648 D.n10620 D.n10612 0.01
R23649 D.n10638 D.n10630 0.01
R23650 D.n10656 D.n10648 0.01
R23651 D.n10674 D.n10666 0.01
R23652 D.n10692 D.n10684 0.01
R23653 D.n10385 D.n10384 0.01
R23654 D.n10365 D.n10364 0.01
R23655 D.n10345 D.n10344 0.01
R23656 D.n10325 D.n10324 0.01
R23657 D.n10305 D.n10304 0.01
R23658 D.n10285 D.n10284 0.01
R23659 D.n10265 D.n10264 0.01
R23660 D.n10245 D.n10244 0.01
R23661 D.n10225 D.n10224 0.01
R23662 D.n10205 D.n10204 0.01
R23663 D.n10185 D.n10184 0.01
R23664 D.n10165 D.n10164 0.01
R23665 D.n9873 D.n9865 0.01
R23666 D.n9891 D.n9883 0.01
R23667 D.n9909 D.n9901 0.01
R23668 D.n9927 D.n9919 0.01
R23669 D.n9945 D.n9937 0.01
R23670 D.n9963 D.n9955 0.01
R23671 D.n9981 D.n9973 0.01
R23672 D.n9999 D.n9991 0.01
R23673 D.n10017 D.n10009 0.01
R23674 D.n10035 D.n10027 0.01
R23675 D.n10053 D.n10045 0.01
R23676 D.n9782 D.n9781 0.01
R23677 D.n9762 D.n9761 0.01
R23678 D.n9742 D.n9741 0.01
R23679 D.n9722 D.n9721 0.01
R23680 D.n9702 D.n9701 0.01
R23681 D.n9682 D.n9681 0.01
R23682 D.n9662 D.n9661 0.01
R23683 D.n9642 D.n9641 0.01
R23684 D.n9622 D.n9621 0.01
R23685 D.n9602 D.n9601 0.01
R23686 D.n9344 D.n9336 0.01
R23687 D.n9362 D.n9354 0.01
R23688 D.n9380 D.n9372 0.01
R23689 D.n9398 D.n9390 0.01
R23690 D.n9416 D.n9408 0.01
R23691 D.n9434 D.n9426 0.01
R23692 D.n9452 D.n9444 0.01
R23693 D.n9470 D.n9462 0.01
R23694 D.n9488 D.n9480 0.01
R23695 D.n9253 D.n9252 0.01
R23696 D.n9233 D.n9232 0.01
R23697 D.n9213 D.n9212 0.01
R23698 D.n9193 D.n9192 0.01
R23699 D.n9173 D.n9172 0.01
R23700 D.n9153 D.n9152 0.01
R23701 D.n9133 D.n9132 0.01
R23702 D.n9113 D.n9112 0.01
R23703 D.n8901 D.n8893 0.01
R23704 D.n8919 D.n8911 0.01
R23705 D.n8937 D.n8929 0.01
R23706 D.n8955 D.n8947 0.01
R23707 D.n8973 D.n8965 0.01
R23708 D.n8991 D.n8983 0.01
R23709 D.n9009 D.n9001 0.01
R23710 D.n8810 D.n8809 0.01
R23711 D.n8790 D.n8789 0.01
R23712 D.n8770 D.n8769 0.01
R23713 D.n8750 D.n8749 0.01
R23714 D.n8730 D.n8729 0.01
R23715 D.n8710 D.n8709 0.01
R23716 D.n8538 D.n8530 0.01
R23717 D.n8556 D.n8548 0.01
R23718 D.n8574 D.n8566 0.01
R23719 D.n8592 D.n8584 0.01
R23720 D.n8610 D.n8602 0.01
R23721 D.n8447 D.n8446 0.01
R23722 D.n8427 D.n8426 0.01
R23723 D.n8407 D.n8406 0.01
R23724 D.n8387 D.n8386 0.01
R23725 D.n8249 D.n8241 0.01
R23726 D.n8267 D.n8259 0.01
R23727 D.n8285 D.n8277 0.01
R23728 D.n8158 D.n8157 0.01
R23729 D.n8138 D.n8137 0.01
R23730 D.n8046 D.n8038 0.01
R23731 D.n8003 D.n8002 0.01
R23732 D.n8019 D.n8018 0.01
R23733 D.n13652 D.n13649 0.01
R23734 D.n13672 D.n13669 0.01
R23735 D.n13651 D.n13650 0.01
R23736 D.n13671 D.n13670 0.01
R23737 D.n12729 D.n12726 0.01
R23738 D.n12745 D.n12742 0.01
R23739 D.n12728 D.n12727 0.01
R23740 D.n12744 D.n12743 0.01
R23741 D.n11880 D.n11877 0.01
R23742 D.n11896 D.n11893 0.01
R23743 D.n11879 D.n11878 0.01
R23744 D.n11895 D.n11894 0.01
R23745 D.n11117 D.n11114 0.01
R23746 D.n11133 D.n11130 0.01
R23747 D.n11116 D.n11115 0.01
R23748 D.n11132 D.n11131 0.01
R23749 D.n10434 D.n10431 0.01
R23750 D.n10450 D.n10447 0.01
R23751 D.n10433 D.n10432 0.01
R23752 D.n10449 D.n10448 0.01
R23753 D.n9831 D.n9828 0.01
R23754 D.n9847 D.n9844 0.01
R23755 D.n9830 D.n9829 0.01
R23756 D.n9846 D.n9845 0.01
R23757 D.n9302 D.n9299 0.01
R23758 D.n9318 D.n9315 0.01
R23759 D.n9301 D.n9300 0.01
R23760 D.n9317 D.n9316 0.01
R23761 D.n8859 D.n8856 0.01
R23762 D.n8875 D.n8872 0.01
R23763 D.n8858 D.n8857 0.01
R23764 D.n8874 D.n8873 0.01
R23765 D.n8496 D.n8493 0.01
R23766 D.n8512 D.n8509 0.01
R23767 D.n8495 D.n8494 0.01
R23768 D.n8511 D.n8510 0.01
R23769 D.n8207 D.n8204 0.01
R23770 D.n8223 D.n8220 0.01
R23771 D.n8206 D.n8205 0.01
R23772 D.n8222 D.n8221 0.01
R23773 D.n8004 D.n8001 0.01
R23774 D.n8020 D.n8017 0.01
R23775 D.n535 D.n534 0.01
R23776 D.n1162 D.n1161 0.01
R23777 D.n1761 D.n1760 0.01
R23778 D.n2332 D.n2331 0.01
R23779 D.n2875 D.n2874 0.01
R23780 D.n3391 D.n3390 0.01
R23781 D.n3879 D.n3878 0.01
R23782 D.n4339 D.n4338 0.01
R23783 D.n4771 D.n4770 0.01
R23784 D.n5175 D.n5174 0.01
R23785 D.n5551 D.n5550 0.01
R23786 D.n5899 D.n5898 0.01
R23787 D.n6219 D.n6218 0.01
R23788 D.n6511 D.n6510 0.01
R23789 D.n6775 D.n6774 0.01
R23790 D.n7011 D.n7010 0.01
R23791 D.n7219 D.n7218 0.01
R23792 D.n7399 D.n7398 0.01
R23793 D.n7551 D.n7550 0.01
R23794 D.n7675 D.n7674 0.01
R23795 D.n7770 D.n7769 0.01
R23796 D.n14081 D.n14080 0.009
R23797 D.n13202 D.n13201 0.009
R23798 D.n13117 D.n13116 0.009
R23799 D.n12319 D.n12318 0.009
R23800 D.n12232 D.n12231 0.009
R23801 D.n11510 D.n11509 0.009
R23802 D.n11433 D.n11432 0.009
R23803 D.n10787 D.n10786 0.009
R23804 D.n10714 D.n10713 0.009
R23805 D.n10144 D.n10143 0.009
R23806 D.n10075 D.n10074 0.009
R23807 D.n9581 D.n9580 0.009
R23808 D.n9510 D.n9509 0.009
R23809 D.n9092 D.n9091 0.009
R23810 D.n9031 D.n9030 0.009
R23811 D.n8689 D.n8688 0.009
R23812 D.n8632 D.n8631 0.009
R23813 D.n8366 D.n8365 0.009
R23814 D.n8307 D.n8306 0.009
R23815 D.n8117 D.n8116 0.009
R23816 D.n8068 D.n8067 0.009
R23817 D.n13667 D.n13666 0.009
R23818 D.n509 D.n508 0.009
R23819 D.n13637 D.n13636 0.009
R23820 D.n12714 D.n12713 0.009
R23821 D.n11865 D.n11864 0.009
R23822 D.n11102 D.n11101 0.009
R23823 D.n10419 D.n10418 0.009
R23824 D.n9816 D.n9815 0.009
R23825 D.n9287 D.n9286 0.009
R23826 D.n8844 D.n8843 0.009
R23827 D.n8481 D.n8480 0.009
R23828 D.n8192 D.n8191 0.009
R23829 D.n7989 D.n7988 0.009
R23830 D.n7952 D.n7951 0.009
R23831 D.n22 D.n21 0.008
R23832 D.n14081 D.n14072 0.008
R23833 D.n13203 D.n13202 0.008
R23834 D.n13117 D.n13108 0.008
R23835 D.n12320 D.n12319 0.008
R23836 D.n12232 D.n12224 0.008
R23837 D.n11511 D.n11510 0.008
R23838 D.n11433 D.n11425 0.008
R23839 D.n10788 D.n10787 0.008
R23840 D.n10714 D.n10706 0.008
R23841 D.n10145 D.n10144 0.008
R23842 D.n10075 D.n10066 0.008
R23843 D.n9582 D.n9581 0.008
R23844 D.n9510 D.n9502 0.008
R23845 D.n9093 D.n9092 0.008
R23846 D.n9031 D.n9023 0.008
R23847 D.n8690 D.n8689 0.008
R23848 D.n8632 D.n8623 0.008
R23849 D.n8367 D.n8366 0.008
R23850 D.n8307 D.n8299 0.008
R23851 D.n8118 D.n8117 0.008
R23852 D.n8068 D.n8060 0.008
R23853 D.n7953 D.n7952 0.008
R23854 D.n13127 D.n13124 0.007
R23855 D.n13127 D.n13119 0.007
R23856 D.n11495 D.n11494 0.007
R23857 D.n11495 D.n11489 0.007
R23858 D.n10772 D.n10771 0.007
R23859 D.n10772 D.n10766 0.007
R23860 D.n10085 D.n10082 0.007
R23861 D.n10085 D.n10077 0.007
R23862 D.n9077 D.n9076 0.007
R23863 D.n9077 D.n9071 0.007
R23864 D.n8642 D.n8639 0.007
R23865 D.n8642 D.n8634 0.007
R23866 D.n8102 D.n8101 0.007
R23867 D.n8102 D.n8096 0.007
R23868 D.n453 D.n445 0.006
R23869 D.n22 D.n19 0.006
R23870 D.n508 D.n502 0.006
R23871 D.n40 D.n37 0.006
R23872 D.n40 D.n39 0.006
R23873 D.n7906 D.n7905 0.006
R23874 D.n535 D.n521 0.006
R23875 D.n1162 D.n1148 0.006
R23876 D.n1761 D.n1747 0.006
R23877 D.n2332 D.n2318 0.006
R23878 D.n2875 D.n2861 0.006
R23879 D.n3391 D.n3377 0.006
R23880 D.n3879 D.n3865 0.006
R23881 D.n4339 D.n4325 0.006
R23882 D.n4771 D.n4757 0.006
R23883 D.n5175 D.n5161 0.006
R23884 D.n5551 D.n5537 0.006
R23885 D.n5899 D.n5885 0.006
R23886 D.n6219 D.n6205 0.006
R23887 D.n6511 D.n6497 0.006
R23888 D.n6775 D.n6761 0.006
R23889 D.n7011 D.n6997 0.006
R23890 D.n7219 D.n7205 0.006
R23891 D.n7399 D.n7385 0.006
R23892 D.n7551 D.n7537 0.006
R23893 D.n7675 D.n7661 0.006
R23894 D.n7770 D.n7756 0.006
R23895 D.n444 D.n436 0.006
R23896 D.n549 D.n537 0.006
R23897 D.n1176 D.n1164 0.006
R23898 D.n1775 D.n1763 0.006
R23899 D.n2346 D.n2334 0.006
R23900 D.n2889 D.n2877 0.006
R23901 D.n3405 D.n3393 0.006
R23902 D.n3893 D.n3881 0.006
R23903 D.n4353 D.n4341 0.006
R23904 D.n4785 D.n4773 0.006
R23905 D.n5189 D.n5177 0.006
R23906 D.n5565 D.n5553 0.006
R23907 D.n5913 D.n5901 0.006
R23908 D.n6233 D.n6221 0.006
R23909 D.n6525 D.n6513 0.006
R23910 D.n6789 D.n6777 0.006
R23911 D.n7025 D.n7013 0.006
R23912 D.n7233 D.n7221 0.006
R23913 D.n7413 D.n7401 0.006
R23914 D.n7565 D.n7553 0.006
R23915 D.n7689 D.n7677 0.006
R23916 D.n7784 D.n7772 0.006
R23917 D.n7832 D.n7831 0.005
R23918 D.n510 D.n509 0.005
R23919 D.n13641 D.n13640 0.005
R23920 D.n12718 D.n12717 0.005
R23921 D.n11869 D.n11868 0.005
R23922 D.n11106 D.n11105 0.005
R23923 D.n10423 D.n10422 0.005
R23924 D.n9820 D.n9819 0.005
R23925 D.n9291 D.n9290 0.005
R23926 D.n8848 D.n8847 0.005
R23927 D.n8485 D.n8484 0.005
R23928 D.n8196 D.n8195 0.005
R23929 D.n7993 D.n7992 0.005
R23930 D.n7968 D.n7967 0.004
R23931 D.n7982 D.n7981 0.004
R23932 D.n13653 D.n13648 0.004
R23933 D.n13673 D.n13664 0.004
R23934 D.n13618 D.n13617 0.004
R23935 D.n13630 D.n13629 0.004
R23936 D.n12730 D.n12725 0.004
R23937 D.n12746 D.n12741 0.004
R23938 D.n12695 D.n12694 0.004
R23939 D.n12707 D.n12706 0.004
R23940 D.n11881 D.n11876 0.004
R23941 D.n11897 D.n11892 0.004
R23942 D.n11846 D.n11845 0.004
R23943 D.n11858 D.n11857 0.004
R23944 D.n11118 D.n11113 0.004
R23945 D.n11134 D.n11129 0.004
R23946 D.n11083 D.n11082 0.004
R23947 D.n11095 D.n11094 0.004
R23948 D.n10435 D.n10430 0.004
R23949 D.n10451 D.n10446 0.004
R23950 D.n10400 D.n10399 0.004
R23951 D.n10412 D.n10411 0.004
R23952 D.n9832 D.n9827 0.004
R23953 D.n9848 D.n9843 0.004
R23954 D.n9797 D.n9796 0.004
R23955 D.n9809 D.n9808 0.004
R23956 D.n9303 D.n9298 0.004
R23957 D.n9319 D.n9314 0.004
R23958 D.n9268 D.n9267 0.004
R23959 D.n9280 D.n9279 0.004
R23960 D.n8860 D.n8855 0.004
R23961 D.n8876 D.n8871 0.004
R23962 D.n8825 D.n8824 0.004
R23963 D.n8837 D.n8836 0.004
R23964 D.n8497 D.n8492 0.004
R23965 D.n8513 D.n8508 0.004
R23966 D.n8462 D.n8461 0.004
R23967 D.n8474 D.n8473 0.004
R23968 D.n8208 D.n8203 0.004
R23969 D.n8224 D.n8219 0.004
R23970 D.n8173 D.n8172 0.004
R23971 D.n8185 D.n8184 0.004
R23972 D.n8005 D.n8000 0.004
R23973 D.n8021 D.n8016 0.004
R23974 D.n13644 D.n13170 0.004
R23975 D.n12721 D.n12287 0.004
R23976 D.n11872 D.n11484 0.004
R23977 D.n11109 D.n10761 0.004
R23978 D.n10426 D.n10112 0.004
R23979 D.n9823 D.n9549 0.004
R23980 D.n9294 D.n9066 0.004
R23981 D.n8851 D.n8657 0.004
R23982 D.n8488 D.n8334 0.004
R23983 D.n8199 D.n8091 0.004
R23984 D.n7996 D.n7922 0.004
R23985 D.n13640 D.n13639 0.004
R23986 D.n12717 D.n12716 0.004
R23987 D.n11868 D.n11867 0.004
R23988 D.n11105 D.n11104 0.004
R23989 D.n10422 D.n10421 0.004
R23990 D.n9819 D.n9818 0.004
R23991 D.n9290 D.n9289 0.004
R23992 D.n8847 D.n8846 0.004
R23993 D.n8484 D.n8483 0.004
R23994 D.n8195 D.n8194 0.004
R23995 D.n7920 D.n7903 0.004
R23996 D.n7917 D.n7906 0.004
R23997 D.n7992 D.n7991 0.004
R23998 D.n13636 D.n13172 0.004
R23999 D.n12713 D.n12289 0.004
R24000 D.n11864 D.n11486 0.004
R24001 D.n11101 D.n10763 0.004
R24002 D.n10418 D.n10114 0.004
R24003 D.n9815 D.n9551 0.004
R24004 D.n9286 D.n9068 0.004
R24005 D.n8843 D.n8659 0.004
R24006 D.n8480 D.n8336 0.004
R24007 D.n8191 D.n8093 0.004
R24008 D.n7988 D.n7975 0.004
R24009 D.n531 D.n530 0.003
R24010 D.n1158 D.n1157 0.003
R24011 D.n1757 D.n1756 0.003
R24012 D.n2328 D.n2327 0.003
R24013 D.n2871 D.n2870 0.003
R24014 D.n3387 D.n3386 0.003
R24015 D.n3875 D.n3874 0.003
R24016 D.n4335 D.n4334 0.003
R24017 D.n4767 D.n4766 0.003
R24018 D.n5171 D.n5170 0.003
R24019 D.n5547 D.n5546 0.003
R24020 D.n5895 D.n5894 0.003
R24021 D.n6215 D.n6214 0.003
R24022 D.n6507 D.n6506 0.003
R24023 D.n6771 D.n6770 0.003
R24024 D.n7007 D.n7006 0.003
R24025 D.n7215 D.n7214 0.003
R24026 D.n7395 D.n7394 0.003
R24027 D.n7547 D.n7546 0.003
R24028 D.n7671 D.n7670 0.003
R24029 D.n7766 D.n7765 0.003
R24030 D.n7858 D.n7857 0.003
R24031 D.n7821 D.n7820 0.003
R24032 D.n7893 D.n7892 0.003
R24033 D.n7977 D.n7976 0.003
R24034 D.n13660 D.n13659 0.003
R24035 D.n13625 D.n13624 0.003
R24036 D.n12737 D.n12736 0.003
R24037 D.n12702 D.n12701 0.003
R24038 D.n11888 D.n11887 0.003
R24039 D.n11853 D.n11852 0.003
R24040 D.n11125 D.n11124 0.003
R24041 D.n11090 D.n11089 0.003
R24042 D.n10442 D.n10441 0.003
R24043 D.n10407 D.n10406 0.003
R24044 D.n9839 D.n9838 0.003
R24045 D.n9804 D.n9803 0.003
R24046 D.n9310 D.n9309 0.003
R24047 D.n9275 D.n9274 0.003
R24048 D.n8867 D.n8866 0.003
R24049 D.n8832 D.n8831 0.003
R24050 D.n8504 D.n8503 0.003
R24051 D.n8469 D.n8468 0.003
R24052 D.n8215 D.n8214 0.003
R24053 D.n8180 D.n8179 0.003
R24054 D.n8012 D.n8011 0.003
R24055 D.n7837 D.n7835 0.003
R24056 D.n7827 D.n7825 0.003
R24057 D.n448 D.n447 0.003
R24058 D.n439 D.n438 0.003
R24059 D.n30 D.n28 0.003
R24060 D.n7957 D.n7955 0.003
R24061 D.n7942 D.n7940 0.003
R24062 D.n14062 D.n14061 0.003
R24063 D.n14044 D.n14043 0.003
R24064 D.n14026 D.n14025 0.003
R24065 D.n14008 D.n14007 0.003
R24066 D.n13990 D.n13989 0.003
R24067 D.n13972 D.n13971 0.003
R24068 D.n13954 D.n13953 0.003
R24069 D.n13936 D.n13935 0.003
R24070 D.n13918 D.n13917 0.003
R24071 D.n13900 D.n13899 0.003
R24072 D.n13882 D.n13881 0.003
R24073 D.n13864 D.n13863 0.003
R24074 D.n13846 D.n13845 0.003
R24075 D.n13828 D.n13827 0.003
R24076 D.n13810 D.n13809 0.003
R24077 D.n13792 D.n13791 0.003
R24078 D.n13774 D.n13773 0.003
R24079 D.n13756 D.n13755 0.003
R24080 D.n13738 D.n13737 0.003
R24081 D.n13720 D.n13719 0.003
R24082 D.n13702 D.n13701 0.003
R24083 D.n13683 D.n13682 0.003
R24084 D.n13693 D.n13691 0.003
R24085 D.n13711 D.n13709 0.003
R24086 D.n13729 D.n13727 0.003
R24087 D.n13747 D.n13745 0.003
R24088 D.n13765 D.n13763 0.003
R24089 D.n13783 D.n13781 0.003
R24090 D.n13801 D.n13799 0.003
R24091 D.n13819 D.n13817 0.003
R24092 D.n13837 D.n13835 0.003
R24093 D.n13855 D.n13853 0.003
R24094 D.n13873 D.n13871 0.003
R24095 D.n13891 D.n13889 0.003
R24096 D.n13909 D.n13907 0.003
R24097 D.n13927 D.n13925 0.003
R24098 D.n13945 D.n13943 0.003
R24099 D.n13963 D.n13961 0.003
R24100 D.n13981 D.n13979 0.003
R24101 D.n13999 D.n13997 0.003
R24102 D.n14017 D.n14015 0.003
R24103 D.n14035 D.n14033 0.003
R24104 D.n14053 D.n14051 0.003
R24105 D.n14075 D.n14073 0.003
R24106 D.n13208 D.n13207 0.003
R24107 D.n13228 D.n13227 0.003
R24108 D.n13248 D.n13247 0.003
R24109 D.n13268 D.n13267 0.003
R24110 D.n13288 D.n13287 0.003
R24111 D.n13308 D.n13307 0.003
R24112 D.n13328 D.n13327 0.003
R24113 D.n13348 D.n13347 0.003
R24114 D.n13368 D.n13367 0.003
R24115 D.n13388 D.n13387 0.003
R24116 D.n13408 D.n13407 0.003
R24117 D.n13428 D.n13427 0.003
R24118 D.n13448 D.n13447 0.003
R24119 D.n13468 D.n13467 0.003
R24120 D.n13488 D.n13487 0.003
R24121 D.n13508 D.n13507 0.003
R24122 D.n13528 D.n13527 0.003
R24123 D.n13548 D.n13547 0.003
R24124 D.n13568 D.n13567 0.003
R24125 D.n13588 D.n13587 0.003
R24126 D.n13608 D.n13607 0.003
R24127 D.n13597 D.n13595 0.003
R24128 D.n13577 D.n13575 0.003
R24129 D.n13557 D.n13555 0.003
R24130 D.n13537 D.n13535 0.003
R24131 D.n13517 D.n13515 0.003
R24132 D.n13497 D.n13495 0.003
R24133 D.n13477 D.n13475 0.003
R24134 D.n13457 D.n13455 0.003
R24135 D.n13437 D.n13435 0.003
R24136 D.n13417 D.n13415 0.003
R24137 D.n13397 D.n13395 0.003
R24138 D.n13377 D.n13375 0.003
R24139 D.n13357 D.n13355 0.003
R24140 D.n13337 D.n13335 0.003
R24141 D.n13317 D.n13315 0.003
R24142 D.n13297 D.n13295 0.003
R24143 D.n13277 D.n13275 0.003
R24144 D.n13257 D.n13255 0.003
R24145 D.n13237 D.n13235 0.003
R24146 D.n13217 D.n13215 0.003
R24147 D.n13192 D.n13190 0.003
R24148 D.n13099 D.n13098 0.003
R24149 D.n13081 D.n13080 0.003
R24150 D.n13063 D.n13062 0.003
R24151 D.n13045 D.n13044 0.003
R24152 D.n13027 D.n13026 0.003
R24153 D.n13009 D.n13008 0.003
R24154 D.n12991 D.n12990 0.003
R24155 D.n12973 D.n12972 0.003
R24156 D.n12955 D.n12954 0.003
R24157 D.n12937 D.n12936 0.003
R24158 D.n12919 D.n12918 0.003
R24159 D.n12901 D.n12900 0.003
R24160 D.n12883 D.n12882 0.003
R24161 D.n12865 D.n12864 0.003
R24162 D.n12847 D.n12846 0.003
R24163 D.n12829 D.n12828 0.003
R24164 D.n12811 D.n12810 0.003
R24165 D.n12793 D.n12792 0.003
R24166 D.n12775 D.n12774 0.003
R24167 D.n12756 D.n12755 0.003
R24168 D.n12766 D.n12764 0.003
R24169 D.n12784 D.n12782 0.003
R24170 D.n12802 D.n12800 0.003
R24171 D.n12820 D.n12818 0.003
R24172 D.n12838 D.n12836 0.003
R24173 D.n12856 D.n12854 0.003
R24174 D.n12874 D.n12872 0.003
R24175 D.n12892 D.n12890 0.003
R24176 D.n12910 D.n12908 0.003
R24177 D.n12928 D.n12926 0.003
R24178 D.n12946 D.n12944 0.003
R24179 D.n12964 D.n12962 0.003
R24180 D.n12982 D.n12980 0.003
R24181 D.n13000 D.n12998 0.003
R24182 D.n13018 D.n13016 0.003
R24183 D.n13036 D.n13034 0.003
R24184 D.n13054 D.n13052 0.003
R24185 D.n13072 D.n13070 0.003
R24186 D.n13090 D.n13088 0.003
R24187 D.n13111 D.n13109 0.003
R24188 D.n12325 D.n12324 0.003
R24189 D.n12345 D.n12344 0.003
R24190 D.n12365 D.n12364 0.003
R24191 D.n12385 D.n12384 0.003
R24192 D.n12405 D.n12404 0.003
R24193 D.n12425 D.n12424 0.003
R24194 D.n12445 D.n12444 0.003
R24195 D.n12465 D.n12464 0.003
R24196 D.n12485 D.n12484 0.003
R24197 D.n12505 D.n12504 0.003
R24198 D.n12525 D.n12524 0.003
R24199 D.n12545 D.n12544 0.003
R24200 D.n12565 D.n12564 0.003
R24201 D.n12585 D.n12584 0.003
R24202 D.n12605 D.n12604 0.003
R24203 D.n12625 D.n12624 0.003
R24204 D.n12645 D.n12644 0.003
R24205 D.n12665 D.n12664 0.003
R24206 D.n12685 D.n12684 0.003
R24207 D.n12674 D.n12672 0.003
R24208 D.n12654 D.n12652 0.003
R24209 D.n12634 D.n12632 0.003
R24210 D.n12614 D.n12612 0.003
R24211 D.n12594 D.n12592 0.003
R24212 D.n12574 D.n12572 0.003
R24213 D.n12554 D.n12552 0.003
R24214 D.n12534 D.n12532 0.003
R24215 D.n12514 D.n12512 0.003
R24216 D.n12494 D.n12492 0.003
R24217 D.n12474 D.n12472 0.003
R24218 D.n12454 D.n12452 0.003
R24219 D.n12434 D.n12432 0.003
R24220 D.n12414 D.n12412 0.003
R24221 D.n12394 D.n12392 0.003
R24222 D.n12374 D.n12372 0.003
R24223 D.n12354 D.n12352 0.003
R24224 D.n12334 D.n12332 0.003
R24225 D.n12309 D.n12307 0.003
R24226 D.n12214 D.n12213 0.003
R24227 D.n12196 D.n12195 0.003
R24228 D.n12178 D.n12177 0.003
R24229 D.n12160 D.n12159 0.003
R24230 D.n12142 D.n12141 0.003
R24231 D.n12124 D.n12123 0.003
R24232 D.n12106 D.n12105 0.003
R24233 D.n12088 D.n12087 0.003
R24234 D.n12070 D.n12069 0.003
R24235 D.n12052 D.n12051 0.003
R24236 D.n12034 D.n12033 0.003
R24237 D.n12016 D.n12015 0.003
R24238 D.n11998 D.n11997 0.003
R24239 D.n11980 D.n11979 0.003
R24240 D.n11962 D.n11961 0.003
R24241 D.n11944 D.n11943 0.003
R24242 D.n11926 D.n11925 0.003
R24243 D.n11907 D.n11906 0.003
R24244 D.n11917 D.n11915 0.003
R24245 D.n11935 D.n11933 0.003
R24246 D.n11953 D.n11951 0.003
R24247 D.n11971 D.n11969 0.003
R24248 D.n11989 D.n11987 0.003
R24249 D.n12007 D.n12005 0.003
R24250 D.n12025 D.n12023 0.003
R24251 D.n12043 D.n12041 0.003
R24252 D.n12061 D.n12059 0.003
R24253 D.n12079 D.n12077 0.003
R24254 D.n12097 D.n12095 0.003
R24255 D.n12115 D.n12113 0.003
R24256 D.n12133 D.n12131 0.003
R24257 D.n12151 D.n12149 0.003
R24258 D.n12169 D.n12167 0.003
R24259 D.n12187 D.n12185 0.003
R24260 D.n12205 D.n12203 0.003
R24261 D.n12227 D.n12225 0.003
R24262 D.n11516 D.n11515 0.003
R24263 D.n11536 D.n11535 0.003
R24264 D.n11556 D.n11555 0.003
R24265 D.n11576 D.n11575 0.003
R24266 D.n11596 D.n11595 0.003
R24267 D.n11616 D.n11615 0.003
R24268 D.n11636 D.n11635 0.003
R24269 D.n11656 D.n11655 0.003
R24270 D.n11676 D.n11675 0.003
R24271 D.n11696 D.n11695 0.003
R24272 D.n11716 D.n11715 0.003
R24273 D.n11736 D.n11735 0.003
R24274 D.n11756 D.n11755 0.003
R24275 D.n11776 D.n11775 0.003
R24276 D.n11796 D.n11795 0.003
R24277 D.n11816 D.n11815 0.003
R24278 D.n11836 D.n11835 0.003
R24279 D.n11825 D.n11823 0.003
R24280 D.n11805 D.n11803 0.003
R24281 D.n11785 D.n11783 0.003
R24282 D.n11765 D.n11763 0.003
R24283 D.n11745 D.n11743 0.003
R24284 D.n11725 D.n11723 0.003
R24285 D.n11705 D.n11703 0.003
R24286 D.n11685 D.n11683 0.003
R24287 D.n11665 D.n11663 0.003
R24288 D.n11645 D.n11643 0.003
R24289 D.n11625 D.n11623 0.003
R24290 D.n11605 D.n11603 0.003
R24291 D.n11585 D.n11583 0.003
R24292 D.n11565 D.n11563 0.003
R24293 D.n11545 D.n11543 0.003
R24294 D.n11525 D.n11523 0.003
R24295 D.n11502 D.n11500 0.003
R24296 D.n11415 D.n11414 0.003
R24297 D.n11397 D.n11396 0.003
R24298 D.n11379 D.n11378 0.003
R24299 D.n11361 D.n11360 0.003
R24300 D.n11343 D.n11342 0.003
R24301 D.n11325 D.n11324 0.003
R24302 D.n11307 D.n11306 0.003
R24303 D.n11289 D.n11288 0.003
R24304 D.n11271 D.n11270 0.003
R24305 D.n11253 D.n11252 0.003
R24306 D.n11235 D.n11234 0.003
R24307 D.n11217 D.n11216 0.003
R24308 D.n11199 D.n11198 0.003
R24309 D.n11181 D.n11180 0.003
R24310 D.n11163 D.n11162 0.003
R24311 D.n11144 D.n11143 0.003
R24312 D.n11154 D.n11152 0.003
R24313 D.n11172 D.n11170 0.003
R24314 D.n11190 D.n11188 0.003
R24315 D.n11208 D.n11206 0.003
R24316 D.n11226 D.n11224 0.003
R24317 D.n11244 D.n11242 0.003
R24318 D.n11262 D.n11260 0.003
R24319 D.n11280 D.n11278 0.003
R24320 D.n11298 D.n11296 0.003
R24321 D.n11316 D.n11314 0.003
R24322 D.n11334 D.n11332 0.003
R24323 D.n11352 D.n11350 0.003
R24324 D.n11370 D.n11368 0.003
R24325 D.n11388 D.n11386 0.003
R24326 D.n11406 D.n11404 0.003
R24327 D.n11428 D.n11426 0.003
R24328 D.n10793 D.n10792 0.003
R24329 D.n10813 D.n10812 0.003
R24330 D.n10833 D.n10832 0.003
R24331 D.n10853 D.n10852 0.003
R24332 D.n10873 D.n10872 0.003
R24333 D.n10893 D.n10892 0.003
R24334 D.n10913 D.n10912 0.003
R24335 D.n10933 D.n10932 0.003
R24336 D.n10953 D.n10952 0.003
R24337 D.n10973 D.n10972 0.003
R24338 D.n10993 D.n10992 0.003
R24339 D.n11013 D.n11012 0.003
R24340 D.n11033 D.n11032 0.003
R24341 D.n11053 D.n11052 0.003
R24342 D.n11073 D.n11072 0.003
R24343 D.n11062 D.n11060 0.003
R24344 D.n11042 D.n11040 0.003
R24345 D.n11022 D.n11020 0.003
R24346 D.n11002 D.n11000 0.003
R24347 D.n10982 D.n10980 0.003
R24348 D.n10962 D.n10960 0.003
R24349 D.n10942 D.n10940 0.003
R24350 D.n10922 D.n10920 0.003
R24351 D.n10902 D.n10900 0.003
R24352 D.n10882 D.n10880 0.003
R24353 D.n10862 D.n10860 0.003
R24354 D.n10842 D.n10840 0.003
R24355 D.n10822 D.n10820 0.003
R24356 D.n10802 D.n10800 0.003
R24357 D.n10779 D.n10777 0.003
R24358 D.n10696 D.n10695 0.003
R24359 D.n10678 D.n10677 0.003
R24360 D.n10660 D.n10659 0.003
R24361 D.n10642 D.n10641 0.003
R24362 D.n10624 D.n10623 0.003
R24363 D.n10606 D.n10605 0.003
R24364 D.n10588 D.n10587 0.003
R24365 D.n10570 D.n10569 0.003
R24366 D.n10552 D.n10551 0.003
R24367 D.n10534 D.n10533 0.003
R24368 D.n10516 D.n10515 0.003
R24369 D.n10498 D.n10497 0.003
R24370 D.n10480 D.n10479 0.003
R24371 D.n10461 D.n10460 0.003
R24372 D.n10471 D.n10469 0.003
R24373 D.n10489 D.n10487 0.003
R24374 D.n10507 D.n10505 0.003
R24375 D.n10525 D.n10523 0.003
R24376 D.n10543 D.n10541 0.003
R24377 D.n10561 D.n10559 0.003
R24378 D.n10579 D.n10577 0.003
R24379 D.n10597 D.n10595 0.003
R24380 D.n10615 D.n10613 0.003
R24381 D.n10633 D.n10631 0.003
R24382 D.n10651 D.n10649 0.003
R24383 D.n10669 D.n10667 0.003
R24384 D.n10687 D.n10685 0.003
R24385 D.n10709 D.n10707 0.003
R24386 D.n10150 D.n10149 0.003
R24387 D.n10170 D.n10169 0.003
R24388 D.n10190 D.n10189 0.003
R24389 D.n10210 D.n10209 0.003
R24390 D.n10230 D.n10229 0.003
R24391 D.n10250 D.n10249 0.003
R24392 D.n10270 D.n10269 0.003
R24393 D.n10290 D.n10289 0.003
R24394 D.n10310 D.n10309 0.003
R24395 D.n10330 D.n10329 0.003
R24396 D.n10350 D.n10349 0.003
R24397 D.n10370 D.n10369 0.003
R24398 D.n10390 D.n10389 0.003
R24399 D.n10379 D.n10377 0.003
R24400 D.n10359 D.n10357 0.003
R24401 D.n10339 D.n10337 0.003
R24402 D.n10319 D.n10317 0.003
R24403 D.n10299 D.n10297 0.003
R24404 D.n10279 D.n10277 0.003
R24405 D.n10259 D.n10257 0.003
R24406 D.n10239 D.n10237 0.003
R24407 D.n10219 D.n10217 0.003
R24408 D.n10199 D.n10197 0.003
R24409 D.n10179 D.n10177 0.003
R24410 D.n10159 D.n10157 0.003
R24411 D.n10134 D.n10132 0.003
R24412 D.n10057 D.n10056 0.003
R24413 D.n10039 D.n10038 0.003
R24414 D.n10021 D.n10020 0.003
R24415 D.n10003 D.n10002 0.003
R24416 D.n9985 D.n9984 0.003
R24417 D.n9967 D.n9966 0.003
R24418 D.n9949 D.n9948 0.003
R24419 D.n9931 D.n9930 0.003
R24420 D.n9913 D.n9912 0.003
R24421 D.n9895 D.n9894 0.003
R24422 D.n9877 D.n9876 0.003
R24423 D.n9858 D.n9857 0.003
R24424 D.n9868 D.n9866 0.003
R24425 D.n9886 D.n9884 0.003
R24426 D.n9904 D.n9902 0.003
R24427 D.n9922 D.n9920 0.003
R24428 D.n9940 D.n9938 0.003
R24429 D.n9958 D.n9956 0.003
R24430 D.n9976 D.n9974 0.003
R24431 D.n9994 D.n9992 0.003
R24432 D.n10012 D.n10010 0.003
R24433 D.n10030 D.n10028 0.003
R24434 D.n10048 D.n10046 0.003
R24435 D.n10069 D.n10067 0.003
R24436 D.n9587 D.n9586 0.003
R24437 D.n9607 D.n9606 0.003
R24438 D.n9627 D.n9626 0.003
R24439 D.n9647 D.n9646 0.003
R24440 D.n9667 D.n9666 0.003
R24441 D.n9687 D.n9686 0.003
R24442 D.n9707 D.n9706 0.003
R24443 D.n9727 D.n9726 0.003
R24444 D.n9747 D.n9746 0.003
R24445 D.n9767 D.n9766 0.003
R24446 D.n9787 D.n9786 0.003
R24447 D.n9776 D.n9774 0.003
R24448 D.n9756 D.n9754 0.003
R24449 D.n9736 D.n9734 0.003
R24450 D.n9716 D.n9714 0.003
R24451 D.n9696 D.n9694 0.003
R24452 D.n9676 D.n9674 0.003
R24453 D.n9656 D.n9654 0.003
R24454 D.n9636 D.n9634 0.003
R24455 D.n9616 D.n9614 0.003
R24456 D.n9596 D.n9594 0.003
R24457 D.n9571 D.n9569 0.003
R24458 D.n9492 D.n9491 0.003
R24459 D.n9474 D.n9473 0.003
R24460 D.n9456 D.n9455 0.003
R24461 D.n9438 D.n9437 0.003
R24462 D.n9420 D.n9419 0.003
R24463 D.n9402 D.n9401 0.003
R24464 D.n9384 D.n9383 0.003
R24465 D.n9366 D.n9365 0.003
R24466 D.n9348 D.n9347 0.003
R24467 D.n9329 D.n9328 0.003
R24468 D.n9339 D.n9337 0.003
R24469 D.n9357 D.n9355 0.003
R24470 D.n9375 D.n9373 0.003
R24471 D.n9393 D.n9391 0.003
R24472 D.n9411 D.n9409 0.003
R24473 D.n9429 D.n9427 0.003
R24474 D.n9447 D.n9445 0.003
R24475 D.n9465 D.n9463 0.003
R24476 D.n9483 D.n9481 0.003
R24477 D.n9505 D.n9503 0.003
R24478 D.n9098 D.n9097 0.003
R24479 D.n9118 D.n9117 0.003
R24480 D.n9138 D.n9137 0.003
R24481 D.n9158 D.n9157 0.003
R24482 D.n9178 D.n9177 0.003
R24483 D.n9198 D.n9197 0.003
R24484 D.n9218 D.n9217 0.003
R24485 D.n9238 D.n9237 0.003
R24486 D.n9258 D.n9257 0.003
R24487 D.n9247 D.n9245 0.003
R24488 D.n9227 D.n9225 0.003
R24489 D.n9207 D.n9205 0.003
R24490 D.n9187 D.n9185 0.003
R24491 D.n9167 D.n9165 0.003
R24492 D.n9147 D.n9145 0.003
R24493 D.n9127 D.n9125 0.003
R24494 D.n9107 D.n9105 0.003
R24495 D.n9084 D.n9082 0.003
R24496 D.n9013 D.n9012 0.003
R24497 D.n8995 D.n8994 0.003
R24498 D.n8977 D.n8976 0.003
R24499 D.n8959 D.n8958 0.003
R24500 D.n8941 D.n8940 0.003
R24501 D.n8923 D.n8922 0.003
R24502 D.n8905 D.n8904 0.003
R24503 D.n8886 D.n8885 0.003
R24504 D.n8896 D.n8894 0.003
R24505 D.n8914 D.n8912 0.003
R24506 D.n8932 D.n8930 0.003
R24507 D.n8950 D.n8948 0.003
R24508 D.n8968 D.n8966 0.003
R24509 D.n8986 D.n8984 0.003
R24510 D.n9004 D.n9002 0.003
R24511 D.n9026 D.n9024 0.003
R24512 D.n8695 D.n8694 0.003
R24513 D.n8715 D.n8714 0.003
R24514 D.n8735 D.n8734 0.003
R24515 D.n8755 D.n8754 0.003
R24516 D.n8775 D.n8774 0.003
R24517 D.n8795 D.n8794 0.003
R24518 D.n8815 D.n8814 0.003
R24519 D.n8804 D.n8802 0.003
R24520 D.n8784 D.n8782 0.003
R24521 D.n8764 D.n8762 0.003
R24522 D.n8744 D.n8742 0.003
R24523 D.n8724 D.n8722 0.003
R24524 D.n8704 D.n8702 0.003
R24525 D.n8679 D.n8677 0.003
R24526 D.n8614 D.n8613 0.003
R24527 D.n8596 D.n8595 0.003
R24528 D.n8578 D.n8577 0.003
R24529 D.n8560 D.n8559 0.003
R24530 D.n8542 D.n8541 0.003
R24531 D.n8523 D.n8522 0.003
R24532 D.n8533 D.n8531 0.003
R24533 D.n8551 D.n8549 0.003
R24534 D.n8569 D.n8567 0.003
R24535 D.n8587 D.n8585 0.003
R24536 D.n8605 D.n8603 0.003
R24537 D.n8626 D.n8624 0.003
R24538 D.n8372 D.n8371 0.003
R24539 D.n8392 D.n8391 0.003
R24540 D.n8412 D.n8411 0.003
R24541 D.n8432 D.n8431 0.003
R24542 D.n8452 D.n8451 0.003
R24543 D.n8441 D.n8439 0.003
R24544 D.n8421 D.n8419 0.003
R24545 D.n8401 D.n8399 0.003
R24546 D.n8381 D.n8379 0.003
R24547 D.n8356 D.n8354 0.003
R24548 D.n8289 D.n8288 0.003
R24549 D.n8271 D.n8270 0.003
R24550 D.n8253 D.n8252 0.003
R24551 D.n8234 D.n8233 0.003
R24552 D.n8244 D.n8242 0.003
R24553 D.n8262 D.n8260 0.003
R24554 D.n8280 D.n8278 0.003
R24555 D.n8302 D.n8300 0.003
R24556 D.n8123 D.n8122 0.003
R24557 D.n8143 D.n8142 0.003
R24558 D.n8163 D.n8162 0.003
R24559 D.n8152 D.n8150 0.003
R24560 D.n8132 D.n8130 0.003
R24561 D.n8109 D.n8107 0.003
R24562 D.n8050 D.n8049 0.003
R24563 D.n8031 D.n8030 0.003
R24564 D.n8041 D.n8039 0.003
R24565 D.n8063 D.n8061 0.003
R24566 D.n52 D.n50 0.003
R24567 D.n61 D.n59 0.003
R24568 D.n70 D.n68 0.003
R24569 D.n79 D.n77 0.003
R24570 D.n88 D.n86 0.003
R24571 D.n97 D.n95 0.003
R24572 D.n106 D.n104 0.003
R24573 D.n115 D.n113 0.003
R24574 D.n124 D.n122 0.003
R24575 D.n133 D.n131 0.003
R24576 D.n142 D.n140 0.003
R24577 D.n151 D.n149 0.003
R24578 D.n160 D.n158 0.003
R24579 D.n169 D.n167 0.003
R24580 D.n178 D.n176 0.003
R24581 D.n187 D.n185 0.003
R24582 D.n196 D.n194 0.003
R24583 D.n205 D.n203 0.003
R24584 D.n214 D.n212 0.003
R24585 D.n223 D.n221 0.003
R24586 D.n232 D.n230 0.003
R24587 D.n241 D.n239 0.003
R24588 D.n250 D.n248 0.003
R24589 D.n259 D.n257 0.003
R24590 D.n268 D.n266 0.003
R24591 D.n277 D.n275 0.003
R24592 D.n286 D.n284 0.003
R24593 D.n295 D.n293 0.003
R24594 D.n304 D.n302 0.003
R24595 D.n313 D.n311 0.003
R24596 D.n322 D.n320 0.003
R24597 D.n331 D.n329 0.003
R24598 D.n340 D.n338 0.003
R24599 D.n349 D.n347 0.003
R24600 D.n358 D.n356 0.003
R24601 D.n367 D.n365 0.003
R24602 D.n376 D.n374 0.003
R24603 D.n385 D.n383 0.003
R24604 D.n394 D.n392 0.003
R24605 D.n403 D.n401 0.003
R24606 D.n412 D.n410 0.003
R24607 D.n421 D.n419 0.003
R24608 D.n430 D.n428 0.003
R24609 D.n524 D.n523 0.003
R24610 D.n540 D.n539 0.003
R24611 D.n1128 D.n1127 0.003
R24612 D.n1114 D.n1113 0.003
R24613 D.n1100 D.n1099 0.003
R24614 D.n1086 D.n1085 0.003
R24615 D.n1072 D.n1071 0.003
R24616 D.n1058 D.n1057 0.003
R24617 D.n1044 D.n1043 0.003
R24618 D.n1030 D.n1029 0.003
R24619 D.n1016 D.n1015 0.003
R24620 D.n1002 D.n1001 0.003
R24621 D.n988 D.n987 0.003
R24622 D.n974 D.n973 0.003
R24623 D.n960 D.n959 0.003
R24624 D.n946 D.n945 0.003
R24625 D.n932 D.n931 0.003
R24626 D.n918 D.n917 0.003
R24627 D.n904 D.n903 0.003
R24628 D.n890 D.n889 0.003
R24629 D.n876 D.n875 0.003
R24630 D.n862 D.n861 0.003
R24631 D.n848 D.n847 0.003
R24632 D.n834 D.n833 0.003
R24633 D.n820 D.n819 0.003
R24634 D.n806 D.n805 0.003
R24635 D.n792 D.n791 0.003
R24636 D.n778 D.n777 0.003
R24637 D.n764 D.n763 0.003
R24638 D.n750 D.n749 0.003
R24639 D.n736 D.n735 0.003
R24640 D.n722 D.n721 0.003
R24641 D.n708 D.n707 0.003
R24642 D.n694 D.n693 0.003
R24643 D.n680 D.n679 0.003
R24644 D.n666 D.n665 0.003
R24645 D.n652 D.n651 0.003
R24646 D.n638 D.n637 0.003
R24647 D.n624 D.n623 0.003
R24648 D.n610 D.n609 0.003
R24649 D.n596 D.n595 0.003
R24650 D.n582 D.n581 0.003
R24651 D.n568 D.n567 0.003
R24652 D.n554 D.n553 0.003
R24653 D.n1151 D.n1150 0.003
R24654 D.n1167 D.n1166 0.003
R24655 D.n1727 D.n1726 0.003
R24656 D.n1713 D.n1712 0.003
R24657 D.n1699 D.n1698 0.003
R24658 D.n1685 D.n1684 0.003
R24659 D.n1671 D.n1670 0.003
R24660 D.n1657 D.n1656 0.003
R24661 D.n1643 D.n1642 0.003
R24662 D.n1629 D.n1628 0.003
R24663 D.n1615 D.n1614 0.003
R24664 D.n1601 D.n1600 0.003
R24665 D.n1587 D.n1586 0.003
R24666 D.n1573 D.n1572 0.003
R24667 D.n1559 D.n1558 0.003
R24668 D.n1545 D.n1544 0.003
R24669 D.n1531 D.n1530 0.003
R24670 D.n1517 D.n1516 0.003
R24671 D.n1503 D.n1502 0.003
R24672 D.n1489 D.n1488 0.003
R24673 D.n1475 D.n1474 0.003
R24674 D.n1461 D.n1460 0.003
R24675 D.n1447 D.n1446 0.003
R24676 D.n1433 D.n1432 0.003
R24677 D.n1419 D.n1418 0.003
R24678 D.n1405 D.n1404 0.003
R24679 D.n1391 D.n1390 0.003
R24680 D.n1377 D.n1376 0.003
R24681 D.n1363 D.n1362 0.003
R24682 D.n1349 D.n1348 0.003
R24683 D.n1335 D.n1334 0.003
R24684 D.n1321 D.n1320 0.003
R24685 D.n1307 D.n1306 0.003
R24686 D.n1293 D.n1292 0.003
R24687 D.n1279 D.n1278 0.003
R24688 D.n1265 D.n1264 0.003
R24689 D.n1251 D.n1250 0.003
R24690 D.n1237 D.n1236 0.003
R24691 D.n1223 D.n1222 0.003
R24692 D.n1209 D.n1208 0.003
R24693 D.n1195 D.n1194 0.003
R24694 D.n1181 D.n1180 0.003
R24695 D.n1750 D.n1749 0.003
R24696 D.n1766 D.n1765 0.003
R24697 D.n2298 D.n2297 0.003
R24698 D.n2284 D.n2283 0.003
R24699 D.n2270 D.n2269 0.003
R24700 D.n2256 D.n2255 0.003
R24701 D.n2242 D.n2241 0.003
R24702 D.n2228 D.n2227 0.003
R24703 D.n2214 D.n2213 0.003
R24704 D.n2200 D.n2199 0.003
R24705 D.n2186 D.n2185 0.003
R24706 D.n2172 D.n2171 0.003
R24707 D.n2158 D.n2157 0.003
R24708 D.n2144 D.n2143 0.003
R24709 D.n2130 D.n2129 0.003
R24710 D.n2116 D.n2115 0.003
R24711 D.n2102 D.n2101 0.003
R24712 D.n2088 D.n2087 0.003
R24713 D.n2074 D.n2073 0.003
R24714 D.n2060 D.n2059 0.003
R24715 D.n2046 D.n2045 0.003
R24716 D.n2032 D.n2031 0.003
R24717 D.n2018 D.n2017 0.003
R24718 D.n2004 D.n2003 0.003
R24719 D.n1990 D.n1989 0.003
R24720 D.n1976 D.n1975 0.003
R24721 D.n1962 D.n1961 0.003
R24722 D.n1948 D.n1947 0.003
R24723 D.n1934 D.n1933 0.003
R24724 D.n1920 D.n1919 0.003
R24725 D.n1906 D.n1905 0.003
R24726 D.n1892 D.n1891 0.003
R24727 D.n1878 D.n1877 0.003
R24728 D.n1864 D.n1863 0.003
R24729 D.n1850 D.n1849 0.003
R24730 D.n1836 D.n1835 0.003
R24731 D.n1822 D.n1821 0.003
R24732 D.n1808 D.n1807 0.003
R24733 D.n1794 D.n1793 0.003
R24734 D.n1780 D.n1779 0.003
R24735 D.n2321 D.n2320 0.003
R24736 D.n2337 D.n2336 0.003
R24737 D.n2841 D.n2840 0.003
R24738 D.n2827 D.n2826 0.003
R24739 D.n2813 D.n2812 0.003
R24740 D.n2799 D.n2798 0.003
R24741 D.n2785 D.n2784 0.003
R24742 D.n2771 D.n2770 0.003
R24743 D.n2757 D.n2756 0.003
R24744 D.n2743 D.n2742 0.003
R24745 D.n2729 D.n2728 0.003
R24746 D.n2715 D.n2714 0.003
R24747 D.n2701 D.n2700 0.003
R24748 D.n2687 D.n2686 0.003
R24749 D.n2673 D.n2672 0.003
R24750 D.n2659 D.n2658 0.003
R24751 D.n2645 D.n2644 0.003
R24752 D.n2631 D.n2630 0.003
R24753 D.n2617 D.n2616 0.003
R24754 D.n2603 D.n2602 0.003
R24755 D.n2589 D.n2588 0.003
R24756 D.n2575 D.n2574 0.003
R24757 D.n2561 D.n2560 0.003
R24758 D.n2547 D.n2546 0.003
R24759 D.n2533 D.n2532 0.003
R24760 D.n2519 D.n2518 0.003
R24761 D.n2505 D.n2504 0.003
R24762 D.n2491 D.n2490 0.003
R24763 D.n2477 D.n2476 0.003
R24764 D.n2463 D.n2462 0.003
R24765 D.n2449 D.n2448 0.003
R24766 D.n2435 D.n2434 0.003
R24767 D.n2421 D.n2420 0.003
R24768 D.n2407 D.n2406 0.003
R24769 D.n2393 D.n2392 0.003
R24770 D.n2379 D.n2378 0.003
R24771 D.n2365 D.n2364 0.003
R24772 D.n2351 D.n2350 0.003
R24773 D.n2864 D.n2863 0.003
R24774 D.n2880 D.n2879 0.003
R24775 D.n3356 D.n3355 0.003
R24776 D.n3342 D.n3341 0.003
R24777 D.n3328 D.n3327 0.003
R24778 D.n3314 D.n3313 0.003
R24779 D.n3300 D.n3299 0.003
R24780 D.n3286 D.n3285 0.003
R24781 D.n3272 D.n3271 0.003
R24782 D.n3258 D.n3257 0.003
R24783 D.n3244 D.n3243 0.003
R24784 D.n3230 D.n3229 0.003
R24785 D.n3216 D.n3215 0.003
R24786 D.n3202 D.n3201 0.003
R24787 D.n3188 D.n3187 0.003
R24788 D.n3174 D.n3173 0.003
R24789 D.n3160 D.n3159 0.003
R24790 D.n3146 D.n3145 0.003
R24791 D.n3132 D.n3131 0.003
R24792 D.n3118 D.n3117 0.003
R24793 D.n3104 D.n3103 0.003
R24794 D.n3090 D.n3089 0.003
R24795 D.n3076 D.n3075 0.003
R24796 D.n3062 D.n3061 0.003
R24797 D.n3048 D.n3047 0.003
R24798 D.n3034 D.n3033 0.003
R24799 D.n3020 D.n3019 0.003
R24800 D.n3006 D.n3005 0.003
R24801 D.n2992 D.n2991 0.003
R24802 D.n2978 D.n2977 0.003
R24803 D.n2964 D.n2963 0.003
R24804 D.n2950 D.n2949 0.003
R24805 D.n2936 D.n2935 0.003
R24806 D.n2922 D.n2921 0.003
R24807 D.n2908 D.n2907 0.003
R24808 D.n2894 D.n2893 0.003
R24809 D.n3380 D.n3379 0.003
R24810 D.n3396 D.n3395 0.003
R24811 D.n3844 D.n3843 0.003
R24812 D.n3830 D.n3829 0.003
R24813 D.n3816 D.n3815 0.003
R24814 D.n3802 D.n3801 0.003
R24815 D.n3788 D.n3787 0.003
R24816 D.n3774 D.n3773 0.003
R24817 D.n3760 D.n3759 0.003
R24818 D.n3746 D.n3745 0.003
R24819 D.n3732 D.n3731 0.003
R24820 D.n3718 D.n3717 0.003
R24821 D.n3704 D.n3703 0.003
R24822 D.n3690 D.n3689 0.003
R24823 D.n3676 D.n3675 0.003
R24824 D.n3662 D.n3661 0.003
R24825 D.n3648 D.n3647 0.003
R24826 D.n3634 D.n3633 0.003
R24827 D.n3620 D.n3619 0.003
R24828 D.n3606 D.n3605 0.003
R24829 D.n3592 D.n3591 0.003
R24830 D.n3578 D.n3577 0.003
R24831 D.n3564 D.n3563 0.003
R24832 D.n3550 D.n3549 0.003
R24833 D.n3536 D.n3535 0.003
R24834 D.n3522 D.n3521 0.003
R24835 D.n3508 D.n3507 0.003
R24836 D.n3494 D.n3493 0.003
R24837 D.n3480 D.n3479 0.003
R24838 D.n3466 D.n3465 0.003
R24839 D.n3452 D.n3451 0.003
R24840 D.n3438 D.n3437 0.003
R24841 D.n3424 D.n3423 0.003
R24842 D.n3410 D.n3409 0.003
R24843 D.n3868 D.n3867 0.003
R24844 D.n3884 D.n3883 0.003
R24845 D.n4304 D.n4303 0.003
R24846 D.n4290 D.n4289 0.003
R24847 D.n4276 D.n4275 0.003
R24848 D.n4262 D.n4261 0.003
R24849 D.n4248 D.n4247 0.003
R24850 D.n4234 D.n4233 0.003
R24851 D.n4220 D.n4219 0.003
R24852 D.n4206 D.n4205 0.003
R24853 D.n4192 D.n4191 0.003
R24854 D.n4178 D.n4177 0.003
R24855 D.n4164 D.n4163 0.003
R24856 D.n4150 D.n4149 0.003
R24857 D.n4136 D.n4135 0.003
R24858 D.n4122 D.n4121 0.003
R24859 D.n4108 D.n4107 0.003
R24860 D.n4094 D.n4093 0.003
R24861 D.n4080 D.n4079 0.003
R24862 D.n4066 D.n4065 0.003
R24863 D.n4052 D.n4051 0.003
R24864 D.n4038 D.n4037 0.003
R24865 D.n4024 D.n4023 0.003
R24866 D.n4010 D.n4009 0.003
R24867 D.n3996 D.n3995 0.003
R24868 D.n3982 D.n3981 0.003
R24869 D.n3968 D.n3967 0.003
R24870 D.n3954 D.n3953 0.003
R24871 D.n3940 D.n3939 0.003
R24872 D.n3926 D.n3925 0.003
R24873 D.n3912 D.n3911 0.003
R24874 D.n3898 D.n3897 0.003
R24875 D.n4328 D.n4327 0.003
R24876 D.n4344 D.n4343 0.003
R24877 D.n4736 D.n4735 0.003
R24878 D.n4722 D.n4721 0.003
R24879 D.n4708 D.n4707 0.003
R24880 D.n4694 D.n4693 0.003
R24881 D.n4680 D.n4679 0.003
R24882 D.n4666 D.n4665 0.003
R24883 D.n4652 D.n4651 0.003
R24884 D.n4638 D.n4637 0.003
R24885 D.n4624 D.n4623 0.003
R24886 D.n4610 D.n4609 0.003
R24887 D.n4596 D.n4595 0.003
R24888 D.n4582 D.n4581 0.003
R24889 D.n4568 D.n4567 0.003
R24890 D.n4554 D.n4553 0.003
R24891 D.n4540 D.n4539 0.003
R24892 D.n4526 D.n4525 0.003
R24893 D.n4512 D.n4511 0.003
R24894 D.n4498 D.n4497 0.003
R24895 D.n4484 D.n4483 0.003
R24896 D.n4470 D.n4469 0.003
R24897 D.n4456 D.n4455 0.003
R24898 D.n4442 D.n4441 0.003
R24899 D.n4428 D.n4427 0.003
R24900 D.n4414 D.n4413 0.003
R24901 D.n4400 D.n4399 0.003
R24902 D.n4386 D.n4385 0.003
R24903 D.n4372 D.n4371 0.003
R24904 D.n4358 D.n4357 0.003
R24905 D.n4760 D.n4759 0.003
R24906 D.n4776 D.n4775 0.003
R24907 D.n5140 D.n5139 0.003
R24908 D.n5126 D.n5125 0.003
R24909 D.n5112 D.n5111 0.003
R24910 D.n5098 D.n5097 0.003
R24911 D.n5084 D.n5083 0.003
R24912 D.n5070 D.n5069 0.003
R24913 D.n5056 D.n5055 0.003
R24914 D.n5042 D.n5041 0.003
R24915 D.n5028 D.n5027 0.003
R24916 D.n5014 D.n5013 0.003
R24917 D.n5000 D.n4999 0.003
R24918 D.n4986 D.n4985 0.003
R24919 D.n4972 D.n4971 0.003
R24920 D.n4958 D.n4957 0.003
R24921 D.n4944 D.n4943 0.003
R24922 D.n4930 D.n4929 0.003
R24923 D.n4916 D.n4915 0.003
R24924 D.n4902 D.n4901 0.003
R24925 D.n4888 D.n4887 0.003
R24926 D.n4874 D.n4873 0.003
R24927 D.n4860 D.n4859 0.003
R24928 D.n4846 D.n4845 0.003
R24929 D.n4832 D.n4831 0.003
R24930 D.n4818 D.n4817 0.003
R24931 D.n4804 D.n4803 0.003
R24932 D.n4790 D.n4789 0.003
R24933 D.n5164 D.n5163 0.003
R24934 D.n5180 D.n5179 0.003
R24935 D.n5516 D.n5515 0.003
R24936 D.n5502 D.n5501 0.003
R24937 D.n5488 D.n5487 0.003
R24938 D.n5474 D.n5473 0.003
R24939 D.n5460 D.n5459 0.003
R24940 D.n5446 D.n5445 0.003
R24941 D.n5432 D.n5431 0.003
R24942 D.n5418 D.n5417 0.003
R24943 D.n5404 D.n5403 0.003
R24944 D.n5390 D.n5389 0.003
R24945 D.n5376 D.n5375 0.003
R24946 D.n5362 D.n5361 0.003
R24947 D.n5348 D.n5347 0.003
R24948 D.n5334 D.n5333 0.003
R24949 D.n5320 D.n5319 0.003
R24950 D.n5306 D.n5305 0.003
R24951 D.n5292 D.n5291 0.003
R24952 D.n5278 D.n5277 0.003
R24953 D.n5264 D.n5263 0.003
R24954 D.n5250 D.n5249 0.003
R24955 D.n5236 D.n5235 0.003
R24956 D.n5222 D.n5221 0.003
R24957 D.n5208 D.n5207 0.003
R24958 D.n5194 D.n5193 0.003
R24959 D.n5540 D.n5539 0.003
R24960 D.n5556 D.n5555 0.003
R24961 D.n5864 D.n5863 0.003
R24962 D.n5850 D.n5849 0.003
R24963 D.n5836 D.n5835 0.003
R24964 D.n5822 D.n5821 0.003
R24965 D.n5808 D.n5807 0.003
R24966 D.n5794 D.n5793 0.003
R24967 D.n5780 D.n5779 0.003
R24968 D.n5766 D.n5765 0.003
R24969 D.n5752 D.n5751 0.003
R24970 D.n5738 D.n5737 0.003
R24971 D.n5724 D.n5723 0.003
R24972 D.n5710 D.n5709 0.003
R24973 D.n5696 D.n5695 0.003
R24974 D.n5682 D.n5681 0.003
R24975 D.n5668 D.n5667 0.003
R24976 D.n5654 D.n5653 0.003
R24977 D.n5640 D.n5639 0.003
R24978 D.n5626 D.n5625 0.003
R24979 D.n5612 D.n5611 0.003
R24980 D.n5598 D.n5597 0.003
R24981 D.n5584 D.n5583 0.003
R24982 D.n5570 D.n5569 0.003
R24983 D.n5888 D.n5887 0.003
R24984 D.n5904 D.n5903 0.003
R24985 D.n6184 D.n6183 0.003
R24986 D.n6170 D.n6169 0.003
R24987 D.n6156 D.n6155 0.003
R24988 D.n6142 D.n6141 0.003
R24989 D.n6128 D.n6127 0.003
R24990 D.n6114 D.n6113 0.003
R24991 D.n6100 D.n6099 0.003
R24992 D.n6086 D.n6085 0.003
R24993 D.n6072 D.n6071 0.003
R24994 D.n6058 D.n6057 0.003
R24995 D.n6044 D.n6043 0.003
R24996 D.n6030 D.n6029 0.003
R24997 D.n6016 D.n6015 0.003
R24998 D.n6002 D.n6001 0.003
R24999 D.n5988 D.n5987 0.003
R25000 D.n5974 D.n5973 0.003
R25001 D.n5960 D.n5959 0.003
R25002 D.n5946 D.n5945 0.003
R25003 D.n5932 D.n5931 0.003
R25004 D.n5918 D.n5917 0.003
R25005 D.n6208 D.n6207 0.003
R25006 D.n6224 D.n6223 0.003
R25007 D.n6476 D.n6475 0.003
R25008 D.n6462 D.n6461 0.003
R25009 D.n6448 D.n6447 0.003
R25010 D.n6434 D.n6433 0.003
R25011 D.n6420 D.n6419 0.003
R25012 D.n6406 D.n6405 0.003
R25013 D.n6392 D.n6391 0.003
R25014 D.n6378 D.n6377 0.003
R25015 D.n6364 D.n6363 0.003
R25016 D.n6350 D.n6349 0.003
R25017 D.n6336 D.n6335 0.003
R25018 D.n6322 D.n6321 0.003
R25019 D.n6308 D.n6307 0.003
R25020 D.n6294 D.n6293 0.003
R25021 D.n6280 D.n6279 0.003
R25022 D.n6266 D.n6265 0.003
R25023 D.n6252 D.n6251 0.003
R25024 D.n6238 D.n6237 0.003
R25025 D.n6500 D.n6499 0.003
R25026 D.n6516 D.n6515 0.003
R25027 D.n6740 D.n6739 0.003
R25028 D.n6726 D.n6725 0.003
R25029 D.n6712 D.n6711 0.003
R25030 D.n6698 D.n6697 0.003
R25031 D.n6684 D.n6683 0.003
R25032 D.n6670 D.n6669 0.003
R25033 D.n6656 D.n6655 0.003
R25034 D.n6642 D.n6641 0.003
R25035 D.n6628 D.n6627 0.003
R25036 D.n6614 D.n6613 0.003
R25037 D.n6600 D.n6599 0.003
R25038 D.n6586 D.n6585 0.003
R25039 D.n6572 D.n6571 0.003
R25040 D.n6558 D.n6557 0.003
R25041 D.n6544 D.n6543 0.003
R25042 D.n6530 D.n6529 0.003
R25043 D.n6764 D.n6763 0.003
R25044 D.n6780 D.n6779 0.003
R25045 D.n6976 D.n6975 0.003
R25046 D.n6962 D.n6961 0.003
R25047 D.n6948 D.n6947 0.003
R25048 D.n6934 D.n6933 0.003
R25049 D.n6920 D.n6919 0.003
R25050 D.n6906 D.n6905 0.003
R25051 D.n6892 D.n6891 0.003
R25052 D.n6878 D.n6877 0.003
R25053 D.n6864 D.n6863 0.003
R25054 D.n6850 D.n6849 0.003
R25055 D.n6836 D.n6835 0.003
R25056 D.n6822 D.n6821 0.003
R25057 D.n6808 D.n6807 0.003
R25058 D.n6794 D.n6793 0.003
R25059 D.n7000 D.n6999 0.003
R25060 D.n7016 D.n7015 0.003
R25061 D.n7184 D.n7183 0.003
R25062 D.n7170 D.n7169 0.003
R25063 D.n7156 D.n7155 0.003
R25064 D.n7142 D.n7141 0.003
R25065 D.n7128 D.n7127 0.003
R25066 D.n7114 D.n7113 0.003
R25067 D.n7100 D.n7099 0.003
R25068 D.n7086 D.n7085 0.003
R25069 D.n7072 D.n7071 0.003
R25070 D.n7058 D.n7057 0.003
R25071 D.n7044 D.n7043 0.003
R25072 D.n7030 D.n7029 0.003
R25073 D.n7208 D.n7207 0.003
R25074 D.n7224 D.n7223 0.003
R25075 D.n7364 D.n7363 0.003
R25076 D.n7350 D.n7349 0.003
R25077 D.n7336 D.n7335 0.003
R25078 D.n7322 D.n7321 0.003
R25079 D.n7308 D.n7307 0.003
R25080 D.n7294 D.n7293 0.003
R25081 D.n7280 D.n7279 0.003
R25082 D.n7266 D.n7265 0.003
R25083 D.n7252 D.n7251 0.003
R25084 D.n7238 D.n7237 0.003
R25085 D.n7388 D.n7387 0.003
R25086 D.n7404 D.n7403 0.003
R25087 D.n7516 D.n7515 0.003
R25088 D.n7502 D.n7501 0.003
R25089 D.n7488 D.n7487 0.003
R25090 D.n7474 D.n7473 0.003
R25091 D.n7460 D.n7459 0.003
R25092 D.n7446 D.n7445 0.003
R25093 D.n7432 D.n7431 0.003
R25094 D.n7418 D.n7417 0.003
R25095 D.n7540 D.n7539 0.003
R25096 D.n7556 D.n7555 0.003
R25097 D.n7640 D.n7639 0.003
R25098 D.n7626 D.n7625 0.003
R25099 D.n7612 D.n7611 0.003
R25100 D.n7598 D.n7597 0.003
R25101 D.n7584 D.n7583 0.003
R25102 D.n7570 D.n7569 0.003
R25103 D.n7664 D.n7663 0.003
R25104 D.n7680 D.n7679 0.003
R25105 D.n7736 D.n7735 0.003
R25106 D.n7722 D.n7721 0.003
R25107 D.n7708 D.n7707 0.003
R25108 D.n7694 D.n7693 0.003
R25109 D.n7759 D.n7758 0.003
R25110 D.n7775 D.n7774 0.003
R25111 D.n7803 D.n7802 0.003
R25112 D.n7789 D.n7788 0.003
R25113 D.n7854 D.n7853 0.003
R25114 D.n7818 D.n7817 0.003
R25115 D.n7840 D.n7838 0.003
R25116 D.n7830 D.n7828 0.003
R25117 D.n451 D.n449 0.003
R25118 D.n442 D.n440 0.003
R25119 D.n33 D.n31 0.003
R25120 D.n7931 D.n7930 0.003
R25121 D.n7960 D.n7958 0.003
R25122 D.n7945 D.n7943 0.003
R25123 D.n14065 D.n14063 0.003
R25124 D.n14047 D.n14045 0.003
R25125 D.n14029 D.n14027 0.003
R25126 D.n14011 D.n14009 0.003
R25127 D.n13993 D.n13991 0.003
R25128 D.n13975 D.n13973 0.003
R25129 D.n13957 D.n13955 0.003
R25130 D.n13939 D.n13937 0.003
R25131 D.n13921 D.n13919 0.003
R25132 D.n13903 D.n13901 0.003
R25133 D.n13885 D.n13883 0.003
R25134 D.n13867 D.n13865 0.003
R25135 D.n13849 D.n13847 0.003
R25136 D.n13831 D.n13829 0.003
R25137 D.n13813 D.n13811 0.003
R25138 D.n13795 D.n13793 0.003
R25139 D.n13777 D.n13775 0.003
R25140 D.n13759 D.n13757 0.003
R25141 D.n13741 D.n13739 0.003
R25142 D.n13723 D.n13721 0.003
R25143 D.n13705 D.n13703 0.003
R25144 D.n13686 D.n13684 0.003
R25145 D.n13696 D.n13694 0.003
R25146 D.n13714 D.n13712 0.003
R25147 D.n13732 D.n13730 0.003
R25148 D.n13750 D.n13748 0.003
R25149 D.n13768 D.n13766 0.003
R25150 D.n13786 D.n13784 0.003
R25151 D.n13804 D.n13802 0.003
R25152 D.n13822 D.n13820 0.003
R25153 D.n13840 D.n13838 0.003
R25154 D.n13858 D.n13856 0.003
R25155 D.n13876 D.n13874 0.003
R25156 D.n13894 D.n13892 0.003
R25157 D.n13912 D.n13910 0.003
R25158 D.n13930 D.n13928 0.003
R25159 D.n13948 D.n13946 0.003
R25160 D.n13966 D.n13964 0.003
R25161 D.n13984 D.n13982 0.003
R25162 D.n14002 D.n14000 0.003
R25163 D.n14020 D.n14018 0.003
R25164 D.n14038 D.n14036 0.003
R25165 D.n14056 D.n14054 0.003
R25166 D.n14078 D.n14076 0.003
R25167 D.n14091 D.n14090 0.003
R25168 D.n13211 D.n13209 0.003
R25169 D.n13231 D.n13229 0.003
R25170 D.n13251 D.n13249 0.003
R25171 D.n13271 D.n13269 0.003
R25172 D.n13291 D.n13289 0.003
R25173 D.n13311 D.n13309 0.003
R25174 D.n13331 D.n13329 0.003
R25175 D.n13351 D.n13349 0.003
R25176 D.n13371 D.n13369 0.003
R25177 D.n13391 D.n13389 0.003
R25178 D.n13411 D.n13409 0.003
R25179 D.n13431 D.n13429 0.003
R25180 D.n13451 D.n13449 0.003
R25181 D.n13471 D.n13469 0.003
R25182 D.n13491 D.n13489 0.003
R25183 D.n13511 D.n13509 0.003
R25184 D.n13531 D.n13529 0.003
R25185 D.n13551 D.n13549 0.003
R25186 D.n13571 D.n13569 0.003
R25187 D.n13591 D.n13589 0.003
R25188 D.n13611 D.n13609 0.003
R25189 D.n13600 D.n13598 0.003
R25190 D.n13580 D.n13578 0.003
R25191 D.n13560 D.n13558 0.003
R25192 D.n13540 D.n13538 0.003
R25193 D.n13520 D.n13518 0.003
R25194 D.n13500 D.n13498 0.003
R25195 D.n13480 D.n13478 0.003
R25196 D.n13460 D.n13458 0.003
R25197 D.n13440 D.n13438 0.003
R25198 D.n13420 D.n13418 0.003
R25199 D.n13400 D.n13398 0.003
R25200 D.n13380 D.n13378 0.003
R25201 D.n13360 D.n13358 0.003
R25202 D.n13340 D.n13338 0.003
R25203 D.n13320 D.n13318 0.003
R25204 D.n13300 D.n13298 0.003
R25205 D.n13280 D.n13278 0.003
R25206 D.n13260 D.n13258 0.003
R25207 D.n13240 D.n13238 0.003
R25208 D.n13220 D.n13218 0.003
R25209 D.n13195 D.n13193 0.003
R25210 D.n13178 D.n13177 0.003
R25211 D.n13102 D.n13100 0.003
R25212 D.n13084 D.n13082 0.003
R25213 D.n13066 D.n13064 0.003
R25214 D.n13048 D.n13046 0.003
R25215 D.n13030 D.n13028 0.003
R25216 D.n13012 D.n13010 0.003
R25217 D.n12994 D.n12992 0.003
R25218 D.n12976 D.n12974 0.003
R25219 D.n12958 D.n12956 0.003
R25220 D.n12940 D.n12938 0.003
R25221 D.n12922 D.n12920 0.003
R25222 D.n12904 D.n12902 0.003
R25223 D.n12886 D.n12884 0.003
R25224 D.n12868 D.n12866 0.003
R25225 D.n12850 D.n12848 0.003
R25226 D.n12832 D.n12830 0.003
R25227 D.n12814 D.n12812 0.003
R25228 D.n12796 D.n12794 0.003
R25229 D.n12778 D.n12776 0.003
R25230 D.n12759 D.n12757 0.003
R25231 D.n12769 D.n12767 0.003
R25232 D.n12787 D.n12785 0.003
R25233 D.n12805 D.n12803 0.003
R25234 D.n12823 D.n12821 0.003
R25235 D.n12841 D.n12839 0.003
R25236 D.n12859 D.n12857 0.003
R25237 D.n12877 D.n12875 0.003
R25238 D.n12895 D.n12893 0.003
R25239 D.n12913 D.n12911 0.003
R25240 D.n12931 D.n12929 0.003
R25241 D.n12949 D.n12947 0.003
R25242 D.n12967 D.n12965 0.003
R25243 D.n12985 D.n12983 0.003
R25244 D.n13003 D.n13001 0.003
R25245 D.n13021 D.n13019 0.003
R25246 D.n13039 D.n13037 0.003
R25247 D.n13057 D.n13055 0.003
R25248 D.n13075 D.n13073 0.003
R25249 D.n13093 D.n13091 0.003
R25250 D.n13114 D.n13112 0.003
R25251 D.n13121 D.n13120 0.003
R25252 D.n12328 D.n12326 0.003
R25253 D.n12348 D.n12346 0.003
R25254 D.n12368 D.n12366 0.003
R25255 D.n12388 D.n12386 0.003
R25256 D.n12408 D.n12406 0.003
R25257 D.n12428 D.n12426 0.003
R25258 D.n12448 D.n12446 0.003
R25259 D.n12468 D.n12466 0.003
R25260 D.n12488 D.n12486 0.003
R25261 D.n12508 D.n12506 0.003
R25262 D.n12528 D.n12526 0.003
R25263 D.n12548 D.n12546 0.003
R25264 D.n12568 D.n12566 0.003
R25265 D.n12588 D.n12586 0.003
R25266 D.n12608 D.n12606 0.003
R25267 D.n12628 D.n12626 0.003
R25268 D.n12648 D.n12646 0.003
R25269 D.n12668 D.n12666 0.003
R25270 D.n12688 D.n12686 0.003
R25271 D.n12677 D.n12675 0.003
R25272 D.n12657 D.n12655 0.003
R25273 D.n12637 D.n12635 0.003
R25274 D.n12617 D.n12615 0.003
R25275 D.n12597 D.n12595 0.003
R25276 D.n12577 D.n12575 0.003
R25277 D.n12557 D.n12555 0.003
R25278 D.n12537 D.n12535 0.003
R25279 D.n12517 D.n12515 0.003
R25280 D.n12497 D.n12495 0.003
R25281 D.n12477 D.n12475 0.003
R25282 D.n12457 D.n12455 0.003
R25283 D.n12437 D.n12435 0.003
R25284 D.n12417 D.n12415 0.003
R25285 D.n12397 D.n12395 0.003
R25286 D.n12377 D.n12375 0.003
R25287 D.n12357 D.n12355 0.003
R25288 D.n12337 D.n12335 0.003
R25289 D.n12312 D.n12310 0.003
R25290 D.n12295 D.n12294 0.003
R25291 D.n12217 D.n12215 0.003
R25292 D.n12199 D.n12197 0.003
R25293 D.n12181 D.n12179 0.003
R25294 D.n12163 D.n12161 0.003
R25295 D.n12145 D.n12143 0.003
R25296 D.n12127 D.n12125 0.003
R25297 D.n12109 D.n12107 0.003
R25298 D.n12091 D.n12089 0.003
R25299 D.n12073 D.n12071 0.003
R25300 D.n12055 D.n12053 0.003
R25301 D.n12037 D.n12035 0.003
R25302 D.n12019 D.n12017 0.003
R25303 D.n12001 D.n11999 0.003
R25304 D.n11983 D.n11981 0.003
R25305 D.n11965 D.n11963 0.003
R25306 D.n11947 D.n11945 0.003
R25307 D.n11929 D.n11927 0.003
R25308 D.n11910 D.n11908 0.003
R25309 D.n11920 D.n11918 0.003
R25310 D.n11938 D.n11936 0.003
R25311 D.n11956 D.n11954 0.003
R25312 D.n11974 D.n11972 0.003
R25313 D.n11992 D.n11990 0.003
R25314 D.n12010 D.n12008 0.003
R25315 D.n12028 D.n12026 0.003
R25316 D.n12046 D.n12044 0.003
R25317 D.n12064 D.n12062 0.003
R25318 D.n12082 D.n12080 0.003
R25319 D.n12100 D.n12098 0.003
R25320 D.n12118 D.n12116 0.003
R25321 D.n12136 D.n12134 0.003
R25322 D.n12154 D.n12152 0.003
R25323 D.n12172 D.n12170 0.003
R25324 D.n12190 D.n12188 0.003
R25325 D.n12208 D.n12206 0.003
R25326 D.n12230 D.n12228 0.003
R25327 D.n12243 D.n12242 0.003
R25328 D.n11519 D.n11517 0.003
R25329 D.n11539 D.n11537 0.003
R25330 D.n11559 D.n11557 0.003
R25331 D.n11579 D.n11577 0.003
R25332 D.n11599 D.n11597 0.003
R25333 D.n11619 D.n11617 0.003
R25334 D.n11639 D.n11637 0.003
R25335 D.n11659 D.n11657 0.003
R25336 D.n11679 D.n11677 0.003
R25337 D.n11699 D.n11697 0.003
R25338 D.n11719 D.n11717 0.003
R25339 D.n11739 D.n11737 0.003
R25340 D.n11759 D.n11757 0.003
R25341 D.n11779 D.n11777 0.003
R25342 D.n11799 D.n11797 0.003
R25343 D.n11819 D.n11817 0.003
R25344 D.n11839 D.n11837 0.003
R25345 D.n11828 D.n11826 0.003
R25346 D.n11808 D.n11806 0.003
R25347 D.n11788 D.n11786 0.003
R25348 D.n11768 D.n11766 0.003
R25349 D.n11748 D.n11746 0.003
R25350 D.n11728 D.n11726 0.003
R25351 D.n11708 D.n11706 0.003
R25352 D.n11688 D.n11686 0.003
R25353 D.n11668 D.n11666 0.003
R25354 D.n11648 D.n11646 0.003
R25355 D.n11628 D.n11626 0.003
R25356 D.n11608 D.n11606 0.003
R25357 D.n11588 D.n11586 0.003
R25358 D.n11568 D.n11566 0.003
R25359 D.n11548 D.n11546 0.003
R25360 D.n11528 D.n11526 0.003
R25361 D.n11505 D.n11503 0.003
R25362 D.n11491 D.n11490 0.003
R25363 D.n11418 D.n11416 0.003
R25364 D.n11400 D.n11398 0.003
R25365 D.n11382 D.n11380 0.003
R25366 D.n11364 D.n11362 0.003
R25367 D.n11346 D.n11344 0.003
R25368 D.n11328 D.n11326 0.003
R25369 D.n11310 D.n11308 0.003
R25370 D.n11292 D.n11290 0.003
R25371 D.n11274 D.n11272 0.003
R25372 D.n11256 D.n11254 0.003
R25373 D.n11238 D.n11236 0.003
R25374 D.n11220 D.n11218 0.003
R25375 D.n11202 D.n11200 0.003
R25376 D.n11184 D.n11182 0.003
R25377 D.n11166 D.n11164 0.003
R25378 D.n11147 D.n11145 0.003
R25379 D.n11157 D.n11155 0.003
R25380 D.n11175 D.n11173 0.003
R25381 D.n11193 D.n11191 0.003
R25382 D.n11211 D.n11209 0.003
R25383 D.n11229 D.n11227 0.003
R25384 D.n11247 D.n11245 0.003
R25385 D.n11265 D.n11263 0.003
R25386 D.n11283 D.n11281 0.003
R25387 D.n11301 D.n11299 0.003
R25388 D.n11319 D.n11317 0.003
R25389 D.n11337 D.n11335 0.003
R25390 D.n11355 D.n11353 0.003
R25391 D.n11373 D.n11371 0.003
R25392 D.n11391 D.n11389 0.003
R25393 D.n11409 D.n11407 0.003
R25394 D.n11431 D.n11429 0.003
R25395 D.n11444 D.n11443 0.003
R25396 D.n10796 D.n10794 0.003
R25397 D.n10816 D.n10814 0.003
R25398 D.n10836 D.n10834 0.003
R25399 D.n10856 D.n10854 0.003
R25400 D.n10876 D.n10874 0.003
R25401 D.n10896 D.n10894 0.003
R25402 D.n10916 D.n10914 0.003
R25403 D.n10936 D.n10934 0.003
R25404 D.n10956 D.n10954 0.003
R25405 D.n10976 D.n10974 0.003
R25406 D.n10996 D.n10994 0.003
R25407 D.n11016 D.n11014 0.003
R25408 D.n11036 D.n11034 0.003
R25409 D.n11056 D.n11054 0.003
R25410 D.n11076 D.n11074 0.003
R25411 D.n11065 D.n11063 0.003
R25412 D.n11045 D.n11043 0.003
R25413 D.n11025 D.n11023 0.003
R25414 D.n11005 D.n11003 0.003
R25415 D.n10985 D.n10983 0.003
R25416 D.n10965 D.n10963 0.003
R25417 D.n10945 D.n10943 0.003
R25418 D.n10925 D.n10923 0.003
R25419 D.n10905 D.n10903 0.003
R25420 D.n10885 D.n10883 0.003
R25421 D.n10865 D.n10863 0.003
R25422 D.n10845 D.n10843 0.003
R25423 D.n10825 D.n10823 0.003
R25424 D.n10805 D.n10803 0.003
R25425 D.n10782 D.n10780 0.003
R25426 D.n10768 D.n10767 0.003
R25427 D.n10699 D.n10697 0.003
R25428 D.n10681 D.n10679 0.003
R25429 D.n10663 D.n10661 0.003
R25430 D.n10645 D.n10643 0.003
R25431 D.n10627 D.n10625 0.003
R25432 D.n10609 D.n10607 0.003
R25433 D.n10591 D.n10589 0.003
R25434 D.n10573 D.n10571 0.003
R25435 D.n10555 D.n10553 0.003
R25436 D.n10537 D.n10535 0.003
R25437 D.n10519 D.n10517 0.003
R25438 D.n10501 D.n10499 0.003
R25439 D.n10483 D.n10481 0.003
R25440 D.n10464 D.n10462 0.003
R25441 D.n10474 D.n10472 0.003
R25442 D.n10492 D.n10490 0.003
R25443 D.n10510 D.n10508 0.003
R25444 D.n10528 D.n10526 0.003
R25445 D.n10546 D.n10544 0.003
R25446 D.n10564 D.n10562 0.003
R25447 D.n10582 D.n10580 0.003
R25448 D.n10600 D.n10598 0.003
R25449 D.n10618 D.n10616 0.003
R25450 D.n10636 D.n10634 0.003
R25451 D.n10654 D.n10652 0.003
R25452 D.n10672 D.n10670 0.003
R25453 D.n10690 D.n10688 0.003
R25454 D.n10712 D.n10710 0.003
R25455 D.n10725 D.n10724 0.003
R25456 D.n10153 D.n10151 0.003
R25457 D.n10173 D.n10171 0.003
R25458 D.n10193 D.n10191 0.003
R25459 D.n10213 D.n10211 0.003
R25460 D.n10233 D.n10231 0.003
R25461 D.n10253 D.n10251 0.003
R25462 D.n10273 D.n10271 0.003
R25463 D.n10293 D.n10291 0.003
R25464 D.n10313 D.n10311 0.003
R25465 D.n10333 D.n10331 0.003
R25466 D.n10353 D.n10351 0.003
R25467 D.n10373 D.n10371 0.003
R25468 D.n10393 D.n10391 0.003
R25469 D.n10382 D.n10380 0.003
R25470 D.n10362 D.n10360 0.003
R25471 D.n10342 D.n10340 0.003
R25472 D.n10322 D.n10320 0.003
R25473 D.n10302 D.n10300 0.003
R25474 D.n10282 D.n10280 0.003
R25475 D.n10262 D.n10260 0.003
R25476 D.n10242 D.n10240 0.003
R25477 D.n10222 D.n10220 0.003
R25478 D.n10202 D.n10200 0.003
R25479 D.n10182 D.n10180 0.003
R25480 D.n10162 D.n10160 0.003
R25481 D.n10137 D.n10135 0.003
R25482 D.n10120 D.n10119 0.003
R25483 D.n10060 D.n10058 0.003
R25484 D.n10042 D.n10040 0.003
R25485 D.n10024 D.n10022 0.003
R25486 D.n10006 D.n10004 0.003
R25487 D.n9988 D.n9986 0.003
R25488 D.n9970 D.n9968 0.003
R25489 D.n9952 D.n9950 0.003
R25490 D.n9934 D.n9932 0.003
R25491 D.n9916 D.n9914 0.003
R25492 D.n9898 D.n9896 0.003
R25493 D.n9880 D.n9878 0.003
R25494 D.n9861 D.n9859 0.003
R25495 D.n9871 D.n9869 0.003
R25496 D.n9889 D.n9887 0.003
R25497 D.n9907 D.n9905 0.003
R25498 D.n9925 D.n9923 0.003
R25499 D.n9943 D.n9941 0.003
R25500 D.n9961 D.n9959 0.003
R25501 D.n9979 D.n9977 0.003
R25502 D.n9997 D.n9995 0.003
R25503 D.n10015 D.n10013 0.003
R25504 D.n10033 D.n10031 0.003
R25505 D.n10051 D.n10049 0.003
R25506 D.n10072 D.n10070 0.003
R25507 D.n10079 D.n10078 0.003
R25508 D.n9590 D.n9588 0.003
R25509 D.n9610 D.n9608 0.003
R25510 D.n9630 D.n9628 0.003
R25511 D.n9650 D.n9648 0.003
R25512 D.n9670 D.n9668 0.003
R25513 D.n9690 D.n9688 0.003
R25514 D.n9710 D.n9708 0.003
R25515 D.n9730 D.n9728 0.003
R25516 D.n9750 D.n9748 0.003
R25517 D.n9770 D.n9768 0.003
R25518 D.n9790 D.n9788 0.003
R25519 D.n9779 D.n9777 0.003
R25520 D.n9759 D.n9757 0.003
R25521 D.n9739 D.n9737 0.003
R25522 D.n9719 D.n9717 0.003
R25523 D.n9699 D.n9697 0.003
R25524 D.n9679 D.n9677 0.003
R25525 D.n9659 D.n9657 0.003
R25526 D.n9639 D.n9637 0.003
R25527 D.n9619 D.n9617 0.003
R25528 D.n9599 D.n9597 0.003
R25529 D.n9574 D.n9572 0.003
R25530 D.n9557 D.n9556 0.003
R25531 D.n9495 D.n9493 0.003
R25532 D.n9477 D.n9475 0.003
R25533 D.n9459 D.n9457 0.003
R25534 D.n9441 D.n9439 0.003
R25535 D.n9423 D.n9421 0.003
R25536 D.n9405 D.n9403 0.003
R25537 D.n9387 D.n9385 0.003
R25538 D.n9369 D.n9367 0.003
R25539 D.n9351 D.n9349 0.003
R25540 D.n9332 D.n9330 0.003
R25541 D.n9342 D.n9340 0.003
R25542 D.n9360 D.n9358 0.003
R25543 D.n9378 D.n9376 0.003
R25544 D.n9396 D.n9394 0.003
R25545 D.n9414 D.n9412 0.003
R25546 D.n9432 D.n9430 0.003
R25547 D.n9450 D.n9448 0.003
R25548 D.n9468 D.n9466 0.003
R25549 D.n9486 D.n9484 0.003
R25550 D.n9508 D.n9506 0.003
R25551 D.n9521 D.n9520 0.003
R25552 D.n9101 D.n9099 0.003
R25553 D.n9121 D.n9119 0.003
R25554 D.n9141 D.n9139 0.003
R25555 D.n9161 D.n9159 0.003
R25556 D.n9181 D.n9179 0.003
R25557 D.n9201 D.n9199 0.003
R25558 D.n9221 D.n9219 0.003
R25559 D.n9241 D.n9239 0.003
R25560 D.n9261 D.n9259 0.003
R25561 D.n9250 D.n9248 0.003
R25562 D.n9230 D.n9228 0.003
R25563 D.n9210 D.n9208 0.003
R25564 D.n9190 D.n9188 0.003
R25565 D.n9170 D.n9168 0.003
R25566 D.n9150 D.n9148 0.003
R25567 D.n9130 D.n9128 0.003
R25568 D.n9110 D.n9108 0.003
R25569 D.n9087 D.n9085 0.003
R25570 D.n9073 D.n9072 0.003
R25571 D.n9016 D.n9014 0.003
R25572 D.n8998 D.n8996 0.003
R25573 D.n8980 D.n8978 0.003
R25574 D.n8962 D.n8960 0.003
R25575 D.n8944 D.n8942 0.003
R25576 D.n8926 D.n8924 0.003
R25577 D.n8908 D.n8906 0.003
R25578 D.n8889 D.n8887 0.003
R25579 D.n8899 D.n8897 0.003
R25580 D.n8917 D.n8915 0.003
R25581 D.n8935 D.n8933 0.003
R25582 D.n8953 D.n8951 0.003
R25583 D.n8971 D.n8969 0.003
R25584 D.n8989 D.n8987 0.003
R25585 D.n9007 D.n9005 0.003
R25586 D.n9029 D.n9027 0.003
R25587 D.n9042 D.n9041 0.003
R25588 D.n8698 D.n8696 0.003
R25589 D.n8718 D.n8716 0.003
R25590 D.n8738 D.n8736 0.003
R25591 D.n8758 D.n8756 0.003
R25592 D.n8778 D.n8776 0.003
R25593 D.n8798 D.n8796 0.003
R25594 D.n8818 D.n8816 0.003
R25595 D.n8807 D.n8805 0.003
R25596 D.n8787 D.n8785 0.003
R25597 D.n8767 D.n8765 0.003
R25598 D.n8747 D.n8745 0.003
R25599 D.n8727 D.n8725 0.003
R25600 D.n8707 D.n8705 0.003
R25601 D.n8682 D.n8680 0.003
R25602 D.n8665 D.n8664 0.003
R25603 D.n8617 D.n8615 0.003
R25604 D.n8599 D.n8597 0.003
R25605 D.n8581 D.n8579 0.003
R25606 D.n8563 D.n8561 0.003
R25607 D.n8545 D.n8543 0.003
R25608 D.n8526 D.n8524 0.003
R25609 D.n8536 D.n8534 0.003
R25610 D.n8554 D.n8552 0.003
R25611 D.n8572 D.n8570 0.003
R25612 D.n8590 D.n8588 0.003
R25613 D.n8608 D.n8606 0.003
R25614 D.n8629 D.n8627 0.003
R25615 D.n8636 D.n8635 0.003
R25616 D.n8375 D.n8373 0.003
R25617 D.n8395 D.n8393 0.003
R25618 D.n8415 D.n8413 0.003
R25619 D.n8435 D.n8433 0.003
R25620 D.n8455 D.n8453 0.003
R25621 D.n8444 D.n8442 0.003
R25622 D.n8424 D.n8422 0.003
R25623 D.n8404 D.n8402 0.003
R25624 D.n8384 D.n8382 0.003
R25625 D.n8359 D.n8357 0.003
R25626 D.n8342 D.n8341 0.003
R25627 D.n8292 D.n8290 0.003
R25628 D.n8274 D.n8272 0.003
R25629 D.n8256 D.n8254 0.003
R25630 D.n8237 D.n8235 0.003
R25631 D.n8247 D.n8245 0.003
R25632 D.n8265 D.n8263 0.003
R25633 D.n8283 D.n8281 0.003
R25634 D.n8305 D.n8303 0.003
R25635 D.n8318 D.n8317 0.003
R25636 D.n8126 D.n8124 0.003
R25637 D.n8146 D.n8144 0.003
R25638 D.n8166 D.n8164 0.003
R25639 D.n8155 D.n8153 0.003
R25640 D.n8135 D.n8133 0.003
R25641 D.n8112 D.n8110 0.003
R25642 D.n8098 D.n8097 0.003
R25643 D.n8053 D.n8051 0.003
R25644 D.n8034 D.n8032 0.003
R25645 D.n8044 D.n8042 0.003
R25646 D.n8066 D.n8064 0.003
R25647 D.n8079 D.n8078 0.003
R25648 D.n7910 D.n7909 0.003
R25649 D.n55 D.n53 0.003
R25650 D.n64 D.n62 0.003
R25651 D.n73 D.n71 0.003
R25652 D.n82 D.n80 0.003
R25653 D.n91 D.n89 0.003
R25654 D.n100 D.n98 0.003
R25655 D.n109 D.n107 0.003
R25656 D.n118 D.n116 0.003
R25657 D.n127 D.n125 0.003
R25658 D.n136 D.n134 0.003
R25659 D.n145 D.n143 0.003
R25660 D.n154 D.n152 0.003
R25661 D.n163 D.n161 0.003
R25662 D.n172 D.n170 0.003
R25663 D.n181 D.n179 0.003
R25664 D.n190 D.n188 0.003
R25665 D.n199 D.n197 0.003
R25666 D.n208 D.n206 0.003
R25667 D.n217 D.n215 0.003
R25668 D.n226 D.n224 0.003
R25669 D.n235 D.n233 0.003
R25670 D.n244 D.n242 0.003
R25671 D.n253 D.n251 0.003
R25672 D.n262 D.n260 0.003
R25673 D.n271 D.n269 0.003
R25674 D.n280 D.n278 0.003
R25675 D.n289 D.n287 0.003
R25676 D.n298 D.n296 0.003
R25677 D.n307 D.n305 0.003
R25678 D.n316 D.n314 0.003
R25679 D.n325 D.n323 0.003
R25680 D.n334 D.n332 0.003
R25681 D.n343 D.n341 0.003
R25682 D.n352 D.n350 0.003
R25683 D.n361 D.n359 0.003
R25684 D.n370 D.n368 0.003
R25685 D.n379 D.n377 0.003
R25686 D.n388 D.n386 0.003
R25687 D.n397 D.n395 0.003
R25688 D.n406 D.n404 0.003
R25689 D.n415 D.n413 0.003
R25690 D.n424 D.n422 0.003
R25691 D.n433 D.n431 0.003
R25692 D.n527 D.n525 0.003
R25693 D.n543 D.n541 0.003
R25694 D.n514 D.n513 0.003
R25695 D.n1131 D.n1129 0.003
R25696 D.n1117 D.n1115 0.003
R25697 D.n1103 D.n1101 0.003
R25698 D.n1089 D.n1087 0.003
R25699 D.n1075 D.n1073 0.003
R25700 D.n1061 D.n1059 0.003
R25701 D.n1047 D.n1045 0.003
R25702 D.n1033 D.n1031 0.003
R25703 D.n1019 D.n1017 0.003
R25704 D.n1005 D.n1003 0.003
R25705 D.n991 D.n989 0.003
R25706 D.n977 D.n975 0.003
R25707 D.n963 D.n961 0.003
R25708 D.n949 D.n947 0.003
R25709 D.n935 D.n933 0.003
R25710 D.n921 D.n919 0.003
R25711 D.n907 D.n905 0.003
R25712 D.n893 D.n891 0.003
R25713 D.n879 D.n877 0.003
R25714 D.n865 D.n863 0.003
R25715 D.n851 D.n849 0.003
R25716 D.n837 D.n835 0.003
R25717 D.n823 D.n821 0.003
R25718 D.n809 D.n807 0.003
R25719 D.n795 D.n793 0.003
R25720 D.n781 D.n779 0.003
R25721 D.n767 D.n765 0.003
R25722 D.n753 D.n751 0.003
R25723 D.n739 D.n737 0.003
R25724 D.n725 D.n723 0.003
R25725 D.n711 D.n709 0.003
R25726 D.n697 D.n695 0.003
R25727 D.n683 D.n681 0.003
R25728 D.n669 D.n667 0.003
R25729 D.n655 D.n653 0.003
R25730 D.n641 D.n639 0.003
R25731 D.n627 D.n625 0.003
R25732 D.n613 D.n611 0.003
R25733 D.n599 D.n597 0.003
R25734 D.n585 D.n583 0.003
R25735 D.n571 D.n569 0.003
R25736 D.n557 D.n555 0.003
R25737 D.n1154 D.n1152 0.003
R25738 D.n1170 D.n1168 0.003
R25739 D.n1144 D.n1143 0.003
R25740 D.n1730 D.n1728 0.003
R25741 D.n1716 D.n1714 0.003
R25742 D.n1702 D.n1700 0.003
R25743 D.n1688 D.n1686 0.003
R25744 D.n1674 D.n1672 0.003
R25745 D.n1660 D.n1658 0.003
R25746 D.n1646 D.n1644 0.003
R25747 D.n1632 D.n1630 0.003
R25748 D.n1618 D.n1616 0.003
R25749 D.n1604 D.n1602 0.003
R25750 D.n1590 D.n1588 0.003
R25751 D.n1576 D.n1574 0.003
R25752 D.n1562 D.n1560 0.003
R25753 D.n1548 D.n1546 0.003
R25754 D.n1534 D.n1532 0.003
R25755 D.n1520 D.n1518 0.003
R25756 D.n1506 D.n1504 0.003
R25757 D.n1492 D.n1490 0.003
R25758 D.n1478 D.n1476 0.003
R25759 D.n1464 D.n1462 0.003
R25760 D.n1450 D.n1448 0.003
R25761 D.n1436 D.n1434 0.003
R25762 D.n1422 D.n1420 0.003
R25763 D.n1408 D.n1406 0.003
R25764 D.n1394 D.n1392 0.003
R25765 D.n1380 D.n1378 0.003
R25766 D.n1366 D.n1364 0.003
R25767 D.n1352 D.n1350 0.003
R25768 D.n1338 D.n1336 0.003
R25769 D.n1324 D.n1322 0.003
R25770 D.n1310 D.n1308 0.003
R25771 D.n1296 D.n1294 0.003
R25772 D.n1282 D.n1280 0.003
R25773 D.n1268 D.n1266 0.003
R25774 D.n1254 D.n1252 0.003
R25775 D.n1240 D.n1238 0.003
R25776 D.n1226 D.n1224 0.003
R25777 D.n1212 D.n1210 0.003
R25778 D.n1198 D.n1196 0.003
R25779 D.n1184 D.n1182 0.003
R25780 D.n1753 D.n1751 0.003
R25781 D.n1769 D.n1767 0.003
R25782 D.n1743 D.n1742 0.003
R25783 D.n2301 D.n2299 0.003
R25784 D.n2287 D.n2285 0.003
R25785 D.n2273 D.n2271 0.003
R25786 D.n2259 D.n2257 0.003
R25787 D.n2245 D.n2243 0.003
R25788 D.n2231 D.n2229 0.003
R25789 D.n2217 D.n2215 0.003
R25790 D.n2203 D.n2201 0.003
R25791 D.n2189 D.n2187 0.003
R25792 D.n2175 D.n2173 0.003
R25793 D.n2161 D.n2159 0.003
R25794 D.n2147 D.n2145 0.003
R25795 D.n2133 D.n2131 0.003
R25796 D.n2119 D.n2117 0.003
R25797 D.n2105 D.n2103 0.003
R25798 D.n2091 D.n2089 0.003
R25799 D.n2077 D.n2075 0.003
R25800 D.n2063 D.n2061 0.003
R25801 D.n2049 D.n2047 0.003
R25802 D.n2035 D.n2033 0.003
R25803 D.n2021 D.n2019 0.003
R25804 D.n2007 D.n2005 0.003
R25805 D.n1993 D.n1991 0.003
R25806 D.n1979 D.n1977 0.003
R25807 D.n1965 D.n1963 0.003
R25808 D.n1951 D.n1949 0.003
R25809 D.n1937 D.n1935 0.003
R25810 D.n1923 D.n1921 0.003
R25811 D.n1909 D.n1907 0.003
R25812 D.n1895 D.n1893 0.003
R25813 D.n1881 D.n1879 0.003
R25814 D.n1867 D.n1865 0.003
R25815 D.n1853 D.n1851 0.003
R25816 D.n1839 D.n1837 0.003
R25817 D.n1825 D.n1823 0.003
R25818 D.n1811 D.n1809 0.003
R25819 D.n1797 D.n1795 0.003
R25820 D.n1783 D.n1781 0.003
R25821 D.n2324 D.n2322 0.003
R25822 D.n2340 D.n2338 0.003
R25823 D.n2314 D.n2313 0.003
R25824 D.n2844 D.n2842 0.003
R25825 D.n2830 D.n2828 0.003
R25826 D.n2816 D.n2814 0.003
R25827 D.n2802 D.n2800 0.003
R25828 D.n2788 D.n2786 0.003
R25829 D.n2774 D.n2772 0.003
R25830 D.n2760 D.n2758 0.003
R25831 D.n2746 D.n2744 0.003
R25832 D.n2732 D.n2730 0.003
R25833 D.n2718 D.n2716 0.003
R25834 D.n2704 D.n2702 0.003
R25835 D.n2690 D.n2688 0.003
R25836 D.n2676 D.n2674 0.003
R25837 D.n2662 D.n2660 0.003
R25838 D.n2648 D.n2646 0.003
R25839 D.n2634 D.n2632 0.003
R25840 D.n2620 D.n2618 0.003
R25841 D.n2606 D.n2604 0.003
R25842 D.n2592 D.n2590 0.003
R25843 D.n2578 D.n2576 0.003
R25844 D.n2564 D.n2562 0.003
R25845 D.n2550 D.n2548 0.003
R25846 D.n2536 D.n2534 0.003
R25847 D.n2522 D.n2520 0.003
R25848 D.n2508 D.n2506 0.003
R25849 D.n2494 D.n2492 0.003
R25850 D.n2480 D.n2478 0.003
R25851 D.n2466 D.n2464 0.003
R25852 D.n2452 D.n2450 0.003
R25853 D.n2438 D.n2436 0.003
R25854 D.n2424 D.n2422 0.003
R25855 D.n2410 D.n2408 0.003
R25856 D.n2396 D.n2394 0.003
R25857 D.n2382 D.n2380 0.003
R25858 D.n2368 D.n2366 0.003
R25859 D.n2354 D.n2352 0.003
R25860 D.n2867 D.n2865 0.003
R25861 D.n2883 D.n2881 0.003
R25862 D.n2857 D.n2856 0.003
R25863 D.n3359 D.n3357 0.003
R25864 D.n3345 D.n3343 0.003
R25865 D.n3331 D.n3329 0.003
R25866 D.n3317 D.n3315 0.003
R25867 D.n3303 D.n3301 0.003
R25868 D.n3289 D.n3287 0.003
R25869 D.n3275 D.n3273 0.003
R25870 D.n3261 D.n3259 0.003
R25871 D.n3247 D.n3245 0.003
R25872 D.n3233 D.n3231 0.003
R25873 D.n3219 D.n3217 0.003
R25874 D.n3205 D.n3203 0.003
R25875 D.n3191 D.n3189 0.003
R25876 D.n3177 D.n3175 0.003
R25877 D.n3163 D.n3161 0.003
R25878 D.n3149 D.n3147 0.003
R25879 D.n3135 D.n3133 0.003
R25880 D.n3121 D.n3119 0.003
R25881 D.n3107 D.n3105 0.003
R25882 D.n3093 D.n3091 0.003
R25883 D.n3079 D.n3077 0.003
R25884 D.n3065 D.n3063 0.003
R25885 D.n3051 D.n3049 0.003
R25886 D.n3037 D.n3035 0.003
R25887 D.n3023 D.n3021 0.003
R25888 D.n3009 D.n3007 0.003
R25889 D.n2995 D.n2993 0.003
R25890 D.n2981 D.n2979 0.003
R25891 D.n2967 D.n2965 0.003
R25892 D.n2953 D.n2951 0.003
R25893 D.n2939 D.n2937 0.003
R25894 D.n2925 D.n2923 0.003
R25895 D.n2911 D.n2909 0.003
R25896 D.n2897 D.n2895 0.003
R25897 D.n3383 D.n3381 0.003
R25898 D.n3399 D.n3397 0.003
R25899 D.n3373 D.n3372 0.003
R25900 D.n3847 D.n3845 0.003
R25901 D.n3833 D.n3831 0.003
R25902 D.n3819 D.n3817 0.003
R25903 D.n3805 D.n3803 0.003
R25904 D.n3791 D.n3789 0.003
R25905 D.n3777 D.n3775 0.003
R25906 D.n3763 D.n3761 0.003
R25907 D.n3749 D.n3747 0.003
R25908 D.n3735 D.n3733 0.003
R25909 D.n3721 D.n3719 0.003
R25910 D.n3707 D.n3705 0.003
R25911 D.n3693 D.n3691 0.003
R25912 D.n3679 D.n3677 0.003
R25913 D.n3665 D.n3663 0.003
R25914 D.n3651 D.n3649 0.003
R25915 D.n3637 D.n3635 0.003
R25916 D.n3623 D.n3621 0.003
R25917 D.n3609 D.n3607 0.003
R25918 D.n3595 D.n3593 0.003
R25919 D.n3581 D.n3579 0.003
R25920 D.n3567 D.n3565 0.003
R25921 D.n3553 D.n3551 0.003
R25922 D.n3539 D.n3537 0.003
R25923 D.n3525 D.n3523 0.003
R25924 D.n3511 D.n3509 0.003
R25925 D.n3497 D.n3495 0.003
R25926 D.n3483 D.n3481 0.003
R25927 D.n3469 D.n3467 0.003
R25928 D.n3455 D.n3453 0.003
R25929 D.n3441 D.n3439 0.003
R25930 D.n3427 D.n3425 0.003
R25931 D.n3413 D.n3411 0.003
R25932 D.n3871 D.n3869 0.003
R25933 D.n3887 D.n3885 0.003
R25934 D.n3861 D.n3860 0.003
R25935 D.n4307 D.n4305 0.003
R25936 D.n4293 D.n4291 0.003
R25937 D.n4279 D.n4277 0.003
R25938 D.n4265 D.n4263 0.003
R25939 D.n4251 D.n4249 0.003
R25940 D.n4237 D.n4235 0.003
R25941 D.n4223 D.n4221 0.003
R25942 D.n4209 D.n4207 0.003
R25943 D.n4195 D.n4193 0.003
R25944 D.n4181 D.n4179 0.003
R25945 D.n4167 D.n4165 0.003
R25946 D.n4153 D.n4151 0.003
R25947 D.n4139 D.n4137 0.003
R25948 D.n4125 D.n4123 0.003
R25949 D.n4111 D.n4109 0.003
R25950 D.n4097 D.n4095 0.003
R25951 D.n4083 D.n4081 0.003
R25952 D.n4069 D.n4067 0.003
R25953 D.n4055 D.n4053 0.003
R25954 D.n4041 D.n4039 0.003
R25955 D.n4027 D.n4025 0.003
R25956 D.n4013 D.n4011 0.003
R25957 D.n3999 D.n3997 0.003
R25958 D.n3985 D.n3983 0.003
R25959 D.n3971 D.n3969 0.003
R25960 D.n3957 D.n3955 0.003
R25961 D.n3943 D.n3941 0.003
R25962 D.n3929 D.n3927 0.003
R25963 D.n3915 D.n3913 0.003
R25964 D.n3901 D.n3899 0.003
R25965 D.n4331 D.n4329 0.003
R25966 D.n4347 D.n4345 0.003
R25967 D.n4321 D.n4320 0.003
R25968 D.n4739 D.n4737 0.003
R25969 D.n4725 D.n4723 0.003
R25970 D.n4711 D.n4709 0.003
R25971 D.n4697 D.n4695 0.003
R25972 D.n4683 D.n4681 0.003
R25973 D.n4669 D.n4667 0.003
R25974 D.n4655 D.n4653 0.003
R25975 D.n4641 D.n4639 0.003
R25976 D.n4627 D.n4625 0.003
R25977 D.n4613 D.n4611 0.003
R25978 D.n4599 D.n4597 0.003
R25979 D.n4585 D.n4583 0.003
R25980 D.n4571 D.n4569 0.003
R25981 D.n4557 D.n4555 0.003
R25982 D.n4543 D.n4541 0.003
R25983 D.n4529 D.n4527 0.003
R25984 D.n4515 D.n4513 0.003
R25985 D.n4501 D.n4499 0.003
R25986 D.n4487 D.n4485 0.003
R25987 D.n4473 D.n4471 0.003
R25988 D.n4459 D.n4457 0.003
R25989 D.n4445 D.n4443 0.003
R25990 D.n4431 D.n4429 0.003
R25991 D.n4417 D.n4415 0.003
R25992 D.n4403 D.n4401 0.003
R25993 D.n4389 D.n4387 0.003
R25994 D.n4375 D.n4373 0.003
R25995 D.n4361 D.n4359 0.003
R25996 D.n4763 D.n4761 0.003
R25997 D.n4779 D.n4777 0.003
R25998 D.n4753 D.n4752 0.003
R25999 D.n5143 D.n5141 0.003
R26000 D.n5129 D.n5127 0.003
R26001 D.n5115 D.n5113 0.003
R26002 D.n5101 D.n5099 0.003
R26003 D.n5087 D.n5085 0.003
R26004 D.n5073 D.n5071 0.003
R26005 D.n5059 D.n5057 0.003
R26006 D.n5045 D.n5043 0.003
R26007 D.n5031 D.n5029 0.003
R26008 D.n5017 D.n5015 0.003
R26009 D.n5003 D.n5001 0.003
R26010 D.n4989 D.n4987 0.003
R26011 D.n4975 D.n4973 0.003
R26012 D.n4961 D.n4959 0.003
R26013 D.n4947 D.n4945 0.003
R26014 D.n4933 D.n4931 0.003
R26015 D.n4919 D.n4917 0.003
R26016 D.n4905 D.n4903 0.003
R26017 D.n4891 D.n4889 0.003
R26018 D.n4877 D.n4875 0.003
R26019 D.n4863 D.n4861 0.003
R26020 D.n4849 D.n4847 0.003
R26021 D.n4835 D.n4833 0.003
R26022 D.n4821 D.n4819 0.003
R26023 D.n4807 D.n4805 0.003
R26024 D.n4793 D.n4791 0.003
R26025 D.n5167 D.n5165 0.003
R26026 D.n5183 D.n5181 0.003
R26027 D.n5157 D.n5156 0.003
R26028 D.n5519 D.n5517 0.003
R26029 D.n5505 D.n5503 0.003
R26030 D.n5491 D.n5489 0.003
R26031 D.n5477 D.n5475 0.003
R26032 D.n5463 D.n5461 0.003
R26033 D.n5449 D.n5447 0.003
R26034 D.n5435 D.n5433 0.003
R26035 D.n5421 D.n5419 0.003
R26036 D.n5407 D.n5405 0.003
R26037 D.n5393 D.n5391 0.003
R26038 D.n5379 D.n5377 0.003
R26039 D.n5365 D.n5363 0.003
R26040 D.n5351 D.n5349 0.003
R26041 D.n5337 D.n5335 0.003
R26042 D.n5323 D.n5321 0.003
R26043 D.n5309 D.n5307 0.003
R26044 D.n5295 D.n5293 0.003
R26045 D.n5281 D.n5279 0.003
R26046 D.n5267 D.n5265 0.003
R26047 D.n5253 D.n5251 0.003
R26048 D.n5239 D.n5237 0.003
R26049 D.n5225 D.n5223 0.003
R26050 D.n5211 D.n5209 0.003
R26051 D.n5197 D.n5195 0.003
R26052 D.n5543 D.n5541 0.003
R26053 D.n5559 D.n5557 0.003
R26054 D.n5533 D.n5532 0.003
R26055 D.n5867 D.n5865 0.003
R26056 D.n5853 D.n5851 0.003
R26057 D.n5839 D.n5837 0.003
R26058 D.n5825 D.n5823 0.003
R26059 D.n5811 D.n5809 0.003
R26060 D.n5797 D.n5795 0.003
R26061 D.n5783 D.n5781 0.003
R26062 D.n5769 D.n5767 0.003
R26063 D.n5755 D.n5753 0.003
R26064 D.n5741 D.n5739 0.003
R26065 D.n5727 D.n5725 0.003
R26066 D.n5713 D.n5711 0.003
R26067 D.n5699 D.n5697 0.003
R26068 D.n5685 D.n5683 0.003
R26069 D.n5671 D.n5669 0.003
R26070 D.n5657 D.n5655 0.003
R26071 D.n5643 D.n5641 0.003
R26072 D.n5629 D.n5627 0.003
R26073 D.n5615 D.n5613 0.003
R26074 D.n5601 D.n5599 0.003
R26075 D.n5587 D.n5585 0.003
R26076 D.n5573 D.n5571 0.003
R26077 D.n5891 D.n5889 0.003
R26078 D.n5907 D.n5905 0.003
R26079 D.n5881 D.n5880 0.003
R26080 D.n6187 D.n6185 0.003
R26081 D.n6173 D.n6171 0.003
R26082 D.n6159 D.n6157 0.003
R26083 D.n6145 D.n6143 0.003
R26084 D.n6131 D.n6129 0.003
R26085 D.n6117 D.n6115 0.003
R26086 D.n6103 D.n6101 0.003
R26087 D.n6089 D.n6087 0.003
R26088 D.n6075 D.n6073 0.003
R26089 D.n6061 D.n6059 0.003
R26090 D.n6047 D.n6045 0.003
R26091 D.n6033 D.n6031 0.003
R26092 D.n6019 D.n6017 0.003
R26093 D.n6005 D.n6003 0.003
R26094 D.n5991 D.n5989 0.003
R26095 D.n5977 D.n5975 0.003
R26096 D.n5963 D.n5961 0.003
R26097 D.n5949 D.n5947 0.003
R26098 D.n5935 D.n5933 0.003
R26099 D.n5921 D.n5919 0.003
R26100 D.n6211 D.n6209 0.003
R26101 D.n6227 D.n6225 0.003
R26102 D.n6201 D.n6200 0.003
R26103 D.n6479 D.n6477 0.003
R26104 D.n6465 D.n6463 0.003
R26105 D.n6451 D.n6449 0.003
R26106 D.n6437 D.n6435 0.003
R26107 D.n6423 D.n6421 0.003
R26108 D.n6409 D.n6407 0.003
R26109 D.n6395 D.n6393 0.003
R26110 D.n6381 D.n6379 0.003
R26111 D.n6367 D.n6365 0.003
R26112 D.n6353 D.n6351 0.003
R26113 D.n6339 D.n6337 0.003
R26114 D.n6325 D.n6323 0.003
R26115 D.n6311 D.n6309 0.003
R26116 D.n6297 D.n6295 0.003
R26117 D.n6283 D.n6281 0.003
R26118 D.n6269 D.n6267 0.003
R26119 D.n6255 D.n6253 0.003
R26120 D.n6241 D.n6239 0.003
R26121 D.n6503 D.n6501 0.003
R26122 D.n6519 D.n6517 0.003
R26123 D.n6493 D.n6492 0.003
R26124 D.n6743 D.n6741 0.003
R26125 D.n6729 D.n6727 0.003
R26126 D.n6715 D.n6713 0.003
R26127 D.n6701 D.n6699 0.003
R26128 D.n6687 D.n6685 0.003
R26129 D.n6673 D.n6671 0.003
R26130 D.n6659 D.n6657 0.003
R26131 D.n6645 D.n6643 0.003
R26132 D.n6631 D.n6629 0.003
R26133 D.n6617 D.n6615 0.003
R26134 D.n6603 D.n6601 0.003
R26135 D.n6589 D.n6587 0.003
R26136 D.n6575 D.n6573 0.003
R26137 D.n6561 D.n6559 0.003
R26138 D.n6547 D.n6545 0.003
R26139 D.n6533 D.n6531 0.003
R26140 D.n6767 D.n6765 0.003
R26141 D.n6783 D.n6781 0.003
R26142 D.n6757 D.n6756 0.003
R26143 D.n6979 D.n6977 0.003
R26144 D.n6965 D.n6963 0.003
R26145 D.n6951 D.n6949 0.003
R26146 D.n6937 D.n6935 0.003
R26147 D.n6923 D.n6921 0.003
R26148 D.n6909 D.n6907 0.003
R26149 D.n6895 D.n6893 0.003
R26150 D.n6881 D.n6879 0.003
R26151 D.n6867 D.n6865 0.003
R26152 D.n6853 D.n6851 0.003
R26153 D.n6839 D.n6837 0.003
R26154 D.n6825 D.n6823 0.003
R26155 D.n6811 D.n6809 0.003
R26156 D.n6797 D.n6795 0.003
R26157 D.n7003 D.n7001 0.003
R26158 D.n7019 D.n7017 0.003
R26159 D.n6993 D.n6992 0.003
R26160 D.n7187 D.n7185 0.003
R26161 D.n7173 D.n7171 0.003
R26162 D.n7159 D.n7157 0.003
R26163 D.n7145 D.n7143 0.003
R26164 D.n7131 D.n7129 0.003
R26165 D.n7117 D.n7115 0.003
R26166 D.n7103 D.n7101 0.003
R26167 D.n7089 D.n7087 0.003
R26168 D.n7075 D.n7073 0.003
R26169 D.n7061 D.n7059 0.003
R26170 D.n7047 D.n7045 0.003
R26171 D.n7033 D.n7031 0.003
R26172 D.n7211 D.n7209 0.003
R26173 D.n7227 D.n7225 0.003
R26174 D.n7201 D.n7200 0.003
R26175 D.n7367 D.n7365 0.003
R26176 D.n7353 D.n7351 0.003
R26177 D.n7339 D.n7337 0.003
R26178 D.n7325 D.n7323 0.003
R26179 D.n7311 D.n7309 0.003
R26180 D.n7297 D.n7295 0.003
R26181 D.n7283 D.n7281 0.003
R26182 D.n7269 D.n7267 0.003
R26183 D.n7255 D.n7253 0.003
R26184 D.n7241 D.n7239 0.003
R26185 D.n7391 D.n7389 0.003
R26186 D.n7407 D.n7405 0.003
R26187 D.n7381 D.n7380 0.003
R26188 D.n7519 D.n7517 0.003
R26189 D.n7505 D.n7503 0.003
R26190 D.n7491 D.n7489 0.003
R26191 D.n7477 D.n7475 0.003
R26192 D.n7463 D.n7461 0.003
R26193 D.n7449 D.n7447 0.003
R26194 D.n7435 D.n7433 0.003
R26195 D.n7421 D.n7419 0.003
R26196 D.n7543 D.n7541 0.003
R26197 D.n7559 D.n7557 0.003
R26198 D.n7533 D.n7532 0.003
R26199 D.n7643 D.n7641 0.003
R26200 D.n7629 D.n7627 0.003
R26201 D.n7615 D.n7613 0.003
R26202 D.n7601 D.n7599 0.003
R26203 D.n7587 D.n7585 0.003
R26204 D.n7573 D.n7571 0.003
R26205 D.n7667 D.n7665 0.003
R26206 D.n7683 D.n7681 0.003
R26207 D.n7657 D.n7656 0.003
R26208 D.n7739 D.n7737 0.003
R26209 D.n7725 D.n7723 0.003
R26210 D.n7711 D.n7709 0.003
R26211 D.n7697 D.n7695 0.003
R26212 D.n7762 D.n7760 0.003
R26213 D.n7778 D.n7776 0.003
R26214 D.n7752 D.n7751 0.003
R26215 D.n7806 D.n7804 0.003
R26216 D.n7792 D.n7790 0.003
R26217 D.n529 D.n528 0.003
R26218 D.n545 D.n544 0.003
R26219 D.n559 D.n558 0.003
R26220 D.n573 D.n572 0.003
R26221 D.n587 D.n586 0.003
R26222 D.n601 D.n600 0.003
R26223 D.n615 D.n614 0.003
R26224 D.n629 D.n628 0.003
R26225 D.n643 D.n642 0.003
R26226 D.n657 D.n656 0.003
R26227 D.n671 D.n670 0.003
R26228 D.n685 D.n684 0.003
R26229 D.n699 D.n698 0.003
R26230 D.n713 D.n712 0.003
R26231 D.n727 D.n726 0.003
R26232 D.n741 D.n740 0.003
R26233 D.n755 D.n754 0.003
R26234 D.n769 D.n768 0.003
R26235 D.n783 D.n782 0.003
R26236 D.n797 D.n796 0.003
R26237 D.n811 D.n810 0.003
R26238 D.n825 D.n824 0.003
R26239 D.n839 D.n838 0.003
R26240 D.n853 D.n852 0.003
R26241 D.n867 D.n866 0.003
R26242 D.n881 D.n880 0.003
R26243 D.n895 D.n894 0.003
R26244 D.n909 D.n908 0.003
R26245 D.n923 D.n922 0.003
R26246 D.n937 D.n936 0.003
R26247 D.n951 D.n950 0.003
R26248 D.n965 D.n964 0.003
R26249 D.n979 D.n978 0.003
R26250 D.n993 D.n992 0.003
R26251 D.n1007 D.n1006 0.003
R26252 D.n1021 D.n1020 0.003
R26253 D.n1035 D.n1034 0.003
R26254 D.n1049 D.n1048 0.003
R26255 D.n1063 D.n1062 0.003
R26256 D.n1077 D.n1076 0.003
R26257 D.n1091 D.n1090 0.003
R26258 D.n1105 D.n1104 0.003
R26259 D.n1119 D.n1118 0.003
R26260 D.n1133 D.n1132 0.003
R26261 D.n1156 D.n1155 0.003
R26262 D.n1172 D.n1171 0.003
R26263 D.n1186 D.n1185 0.003
R26264 D.n1200 D.n1199 0.003
R26265 D.n1214 D.n1213 0.003
R26266 D.n1228 D.n1227 0.003
R26267 D.n1242 D.n1241 0.003
R26268 D.n1256 D.n1255 0.003
R26269 D.n1270 D.n1269 0.003
R26270 D.n1284 D.n1283 0.003
R26271 D.n1298 D.n1297 0.003
R26272 D.n1312 D.n1311 0.003
R26273 D.n1326 D.n1325 0.003
R26274 D.n1340 D.n1339 0.003
R26275 D.n1354 D.n1353 0.003
R26276 D.n1368 D.n1367 0.003
R26277 D.n1382 D.n1381 0.003
R26278 D.n1396 D.n1395 0.003
R26279 D.n1410 D.n1409 0.003
R26280 D.n1424 D.n1423 0.003
R26281 D.n1438 D.n1437 0.003
R26282 D.n1452 D.n1451 0.003
R26283 D.n1466 D.n1465 0.003
R26284 D.n1480 D.n1479 0.003
R26285 D.n1494 D.n1493 0.003
R26286 D.n1508 D.n1507 0.003
R26287 D.n1522 D.n1521 0.003
R26288 D.n1536 D.n1535 0.003
R26289 D.n1550 D.n1549 0.003
R26290 D.n1564 D.n1563 0.003
R26291 D.n1578 D.n1577 0.003
R26292 D.n1592 D.n1591 0.003
R26293 D.n1606 D.n1605 0.003
R26294 D.n1620 D.n1619 0.003
R26295 D.n1634 D.n1633 0.003
R26296 D.n1648 D.n1647 0.003
R26297 D.n1662 D.n1661 0.003
R26298 D.n1676 D.n1675 0.003
R26299 D.n1690 D.n1689 0.003
R26300 D.n1704 D.n1703 0.003
R26301 D.n1718 D.n1717 0.003
R26302 D.n1732 D.n1731 0.003
R26303 D.n1755 D.n1754 0.003
R26304 D.n1771 D.n1770 0.003
R26305 D.n1785 D.n1784 0.003
R26306 D.n1799 D.n1798 0.003
R26307 D.n1813 D.n1812 0.003
R26308 D.n1827 D.n1826 0.003
R26309 D.n1841 D.n1840 0.003
R26310 D.n1855 D.n1854 0.003
R26311 D.n1869 D.n1868 0.003
R26312 D.n1883 D.n1882 0.003
R26313 D.n1897 D.n1896 0.003
R26314 D.n1911 D.n1910 0.003
R26315 D.n1925 D.n1924 0.003
R26316 D.n1939 D.n1938 0.003
R26317 D.n1953 D.n1952 0.003
R26318 D.n1967 D.n1966 0.003
R26319 D.n1981 D.n1980 0.003
R26320 D.n1995 D.n1994 0.003
R26321 D.n2009 D.n2008 0.003
R26322 D.n2023 D.n2022 0.003
R26323 D.n2037 D.n2036 0.003
R26324 D.n2051 D.n2050 0.003
R26325 D.n2065 D.n2064 0.003
R26326 D.n2079 D.n2078 0.003
R26327 D.n2093 D.n2092 0.003
R26328 D.n2107 D.n2106 0.003
R26329 D.n2121 D.n2120 0.003
R26330 D.n2135 D.n2134 0.003
R26331 D.n2149 D.n2148 0.003
R26332 D.n2163 D.n2162 0.003
R26333 D.n2177 D.n2176 0.003
R26334 D.n2191 D.n2190 0.003
R26335 D.n2205 D.n2204 0.003
R26336 D.n2219 D.n2218 0.003
R26337 D.n2233 D.n2232 0.003
R26338 D.n2247 D.n2246 0.003
R26339 D.n2261 D.n2260 0.003
R26340 D.n2275 D.n2274 0.003
R26341 D.n2289 D.n2288 0.003
R26342 D.n2303 D.n2302 0.003
R26343 D.n2326 D.n2325 0.003
R26344 D.n2342 D.n2341 0.003
R26345 D.n2356 D.n2355 0.003
R26346 D.n2370 D.n2369 0.003
R26347 D.n2384 D.n2383 0.003
R26348 D.n2398 D.n2397 0.003
R26349 D.n2412 D.n2411 0.003
R26350 D.n2426 D.n2425 0.003
R26351 D.n2440 D.n2439 0.003
R26352 D.n2454 D.n2453 0.003
R26353 D.n2468 D.n2467 0.003
R26354 D.n2482 D.n2481 0.003
R26355 D.n2496 D.n2495 0.003
R26356 D.n2510 D.n2509 0.003
R26357 D.n2524 D.n2523 0.003
R26358 D.n2538 D.n2537 0.003
R26359 D.n2552 D.n2551 0.003
R26360 D.n2566 D.n2565 0.003
R26361 D.n2580 D.n2579 0.003
R26362 D.n2594 D.n2593 0.003
R26363 D.n2608 D.n2607 0.003
R26364 D.n2622 D.n2621 0.003
R26365 D.n2636 D.n2635 0.003
R26366 D.n2650 D.n2649 0.003
R26367 D.n2664 D.n2663 0.003
R26368 D.n2678 D.n2677 0.003
R26369 D.n2692 D.n2691 0.003
R26370 D.n2706 D.n2705 0.003
R26371 D.n2720 D.n2719 0.003
R26372 D.n2734 D.n2733 0.003
R26373 D.n2748 D.n2747 0.003
R26374 D.n2762 D.n2761 0.003
R26375 D.n2776 D.n2775 0.003
R26376 D.n2790 D.n2789 0.003
R26377 D.n2804 D.n2803 0.003
R26378 D.n2818 D.n2817 0.003
R26379 D.n2832 D.n2831 0.003
R26380 D.n2846 D.n2845 0.003
R26381 D.n2869 D.n2868 0.003
R26382 D.n2885 D.n2884 0.003
R26383 D.n2899 D.n2898 0.003
R26384 D.n2913 D.n2912 0.003
R26385 D.n2927 D.n2926 0.003
R26386 D.n2941 D.n2940 0.003
R26387 D.n2955 D.n2954 0.003
R26388 D.n2969 D.n2968 0.003
R26389 D.n2983 D.n2982 0.003
R26390 D.n2997 D.n2996 0.003
R26391 D.n3011 D.n3010 0.003
R26392 D.n3025 D.n3024 0.003
R26393 D.n3039 D.n3038 0.003
R26394 D.n3053 D.n3052 0.003
R26395 D.n3067 D.n3066 0.003
R26396 D.n3081 D.n3080 0.003
R26397 D.n3095 D.n3094 0.003
R26398 D.n3109 D.n3108 0.003
R26399 D.n3123 D.n3122 0.003
R26400 D.n3137 D.n3136 0.003
R26401 D.n3151 D.n3150 0.003
R26402 D.n3165 D.n3164 0.003
R26403 D.n3179 D.n3178 0.003
R26404 D.n3193 D.n3192 0.003
R26405 D.n3207 D.n3206 0.003
R26406 D.n3221 D.n3220 0.003
R26407 D.n3235 D.n3234 0.003
R26408 D.n3249 D.n3248 0.003
R26409 D.n3263 D.n3262 0.003
R26410 D.n3277 D.n3276 0.003
R26411 D.n3291 D.n3290 0.003
R26412 D.n3305 D.n3304 0.003
R26413 D.n3319 D.n3318 0.003
R26414 D.n3333 D.n3332 0.003
R26415 D.n3347 D.n3346 0.003
R26416 D.n3361 D.n3360 0.003
R26417 D.n3385 D.n3384 0.003
R26418 D.n3401 D.n3400 0.003
R26419 D.n3415 D.n3414 0.003
R26420 D.n3429 D.n3428 0.003
R26421 D.n3443 D.n3442 0.003
R26422 D.n3457 D.n3456 0.003
R26423 D.n3471 D.n3470 0.003
R26424 D.n3485 D.n3484 0.003
R26425 D.n3499 D.n3498 0.003
R26426 D.n3513 D.n3512 0.003
R26427 D.n3527 D.n3526 0.003
R26428 D.n3541 D.n3540 0.003
R26429 D.n3555 D.n3554 0.003
R26430 D.n3569 D.n3568 0.003
R26431 D.n3583 D.n3582 0.003
R26432 D.n3597 D.n3596 0.003
R26433 D.n3611 D.n3610 0.003
R26434 D.n3625 D.n3624 0.003
R26435 D.n3639 D.n3638 0.003
R26436 D.n3653 D.n3652 0.003
R26437 D.n3667 D.n3666 0.003
R26438 D.n3681 D.n3680 0.003
R26439 D.n3695 D.n3694 0.003
R26440 D.n3709 D.n3708 0.003
R26441 D.n3723 D.n3722 0.003
R26442 D.n3737 D.n3736 0.003
R26443 D.n3751 D.n3750 0.003
R26444 D.n3765 D.n3764 0.003
R26445 D.n3779 D.n3778 0.003
R26446 D.n3793 D.n3792 0.003
R26447 D.n3807 D.n3806 0.003
R26448 D.n3821 D.n3820 0.003
R26449 D.n3835 D.n3834 0.003
R26450 D.n3849 D.n3848 0.003
R26451 D.n3873 D.n3872 0.003
R26452 D.n3889 D.n3888 0.003
R26453 D.n3903 D.n3902 0.003
R26454 D.n3917 D.n3916 0.003
R26455 D.n3931 D.n3930 0.003
R26456 D.n3945 D.n3944 0.003
R26457 D.n3959 D.n3958 0.003
R26458 D.n3973 D.n3972 0.003
R26459 D.n3987 D.n3986 0.003
R26460 D.n4001 D.n4000 0.003
R26461 D.n4015 D.n4014 0.003
R26462 D.n4029 D.n4028 0.003
R26463 D.n4043 D.n4042 0.003
R26464 D.n4057 D.n4056 0.003
R26465 D.n4071 D.n4070 0.003
R26466 D.n4085 D.n4084 0.003
R26467 D.n4099 D.n4098 0.003
R26468 D.n4113 D.n4112 0.003
R26469 D.n4127 D.n4126 0.003
R26470 D.n4141 D.n4140 0.003
R26471 D.n4155 D.n4154 0.003
R26472 D.n4169 D.n4168 0.003
R26473 D.n4183 D.n4182 0.003
R26474 D.n4197 D.n4196 0.003
R26475 D.n4211 D.n4210 0.003
R26476 D.n4225 D.n4224 0.003
R26477 D.n4239 D.n4238 0.003
R26478 D.n4253 D.n4252 0.003
R26479 D.n4267 D.n4266 0.003
R26480 D.n4281 D.n4280 0.003
R26481 D.n4295 D.n4294 0.003
R26482 D.n4309 D.n4308 0.003
R26483 D.n4333 D.n4332 0.003
R26484 D.n4349 D.n4348 0.003
R26485 D.n4363 D.n4362 0.003
R26486 D.n4377 D.n4376 0.003
R26487 D.n4391 D.n4390 0.003
R26488 D.n4405 D.n4404 0.003
R26489 D.n4419 D.n4418 0.003
R26490 D.n4433 D.n4432 0.003
R26491 D.n4447 D.n4446 0.003
R26492 D.n4461 D.n4460 0.003
R26493 D.n4475 D.n4474 0.003
R26494 D.n4489 D.n4488 0.003
R26495 D.n4503 D.n4502 0.003
R26496 D.n4517 D.n4516 0.003
R26497 D.n4531 D.n4530 0.003
R26498 D.n4545 D.n4544 0.003
R26499 D.n4559 D.n4558 0.003
R26500 D.n4573 D.n4572 0.003
R26501 D.n4587 D.n4586 0.003
R26502 D.n4601 D.n4600 0.003
R26503 D.n4615 D.n4614 0.003
R26504 D.n4629 D.n4628 0.003
R26505 D.n4643 D.n4642 0.003
R26506 D.n4657 D.n4656 0.003
R26507 D.n4671 D.n4670 0.003
R26508 D.n4685 D.n4684 0.003
R26509 D.n4699 D.n4698 0.003
R26510 D.n4713 D.n4712 0.003
R26511 D.n4727 D.n4726 0.003
R26512 D.n4741 D.n4740 0.003
R26513 D.n4765 D.n4764 0.003
R26514 D.n4781 D.n4780 0.003
R26515 D.n4795 D.n4794 0.003
R26516 D.n4809 D.n4808 0.003
R26517 D.n4823 D.n4822 0.003
R26518 D.n4837 D.n4836 0.003
R26519 D.n4851 D.n4850 0.003
R26520 D.n4865 D.n4864 0.003
R26521 D.n4879 D.n4878 0.003
R26522 D.n4893 D.n4892 0.003
R26523 D.n4907 D.n4906 0.003
R26524 D.n4921 D.n4920 0.003
R26525 D.n4935 D.n4934 0.003
R26526 D.n4949 D.n4948 0.003
R26527 D.n4963 D.n4962 0.003
R26528 D.n4977 D.n4976 0.003
R26529 D.n4991 D.n4990 0.003
R26530 D.n5005 D.n5004 0.003
R26531 D.n5019 D.n5018 0.003
R26532 D.n5033 D.n5032 0.003
R26533 D.n5047 D.n5046 0.003
R26534 D.n5061 D.n5060 0.003
R26535 D.n5075 D.n5074 0.003
R26536 D.n5089 D.n5088 0.003
R26537 D.n5103 D.n5102 0.003
R26538 D.n5117 D.n5116 0.003
R26539 D.n5131 D.n5130 0.003
R26540 D.n5145 D.n5144 0.003
R26541 D.n5169 D.n5168 0.003
R26542 D.n5185 D.n5184 0.003
R26543 D.n5199 D.n5198 0.003
R26544 D.n5213 D.n5212 0.003
R26545 D.n5227 D.n5226 0.003
R26546 D.n5241 D.n5240 0.003
R26547 D.n5255 D.n5254 0.003
R26548 D.n5269 D.n5268 0.003
R26549 D.n5283 D.n5282 0.003
R26550 D.n5297 D.n5296 0.003
R26551 D.n5311 D.n5310 0.003
R26552 D.n5325 D.n5324 0.003
R26553 D.n5339 D.n5338 0.003
R26554 D.n5353 D.n5352 0.003
R26555 D.n5367 D.n5366 0.003
R26556 D.n5381 D.n5380 0.003
R26557 D.n5395 D.n5394 0.003
R26558 D.n5409 D.n5408 0.003
R26559 D.n5423 D.n5422 0.003
R26560 D.n5437 D.n5436 0.003
R26561 D.n5451 D.n5450 0.003
R26562 D.n5465 D.n5464 0.003
R26563 D.n5479 D.n5478 0.003
R26564 D.n5493 D.n5492 0.003
R26565 D.n5507 D.n5506 0.003
R26566 D.n5521 D.n5520 0.003
R26567 D.n5545 D.n5544 0.003
R26568 D.n5561 D.n5560 0.003
R26569 D.n5575 D.n5574 0.003
R26570 D.n5589 D.n5588 0.003
R26571 D.n5603 D.n5602 0.003
R26572 D.n5617 D.n5616 0.003
R26573 D.n5631 D.n5630 0.003
R26574 D.n5645 D.n5644 0.003
R26575 D.n5659 D.n5658 0.003
R26576 D.n5673 D.n5672 0.003
R26577 D.n5687 D.n5686 0.003
R26578 D.n5701 D.n5700 0.003
R26579 D.n5715 D.n5714 0.003
R26580 D.n5729 D.n5728 0.003
R26581 D.n5743 D.n5742 0.003
R26582 D.n5757 D.n5756 0.003
R26583 D.n5771 D.n5770 0.003
R26584 D.n5785 D.n5784 0.003
R26585 D.n5799 D.n5798 0.003
R26586 D.n5813 D.n5812 0.003
R26587 D.n5827 D.n5826 0.003
R26588 D.n5841 D.n5840 0.003
R26589 D.n5855 D.n5854 0.003
R26590 D.n5869 D.n5868 0.003
R26591 D.n5893 D.n5892 0.003
R26592 D.n5909 D.n5908 0.003
R26593 D.n5923 D.n5922 0.003
R26594 D.n5937 D.n5936 0.003
R26595 D.n5951 D.n5950 0.003
R26596 D.n5965 D.n5964 0.003
R26597 D.n5979 D.n5978 0.003
R26598 D.n5993 D.n5992 0.003
R26599 D.n6007 D.n6006 0.003
R26600 D.n6021 D.n6020 0.003
R26601 D.n6035 D.n6034 0.003
R26602 D.n6049 D.n6048 0.003
R26603 D.n6063 D.n6062 0.003
R26604 D.n6077 D.n6076 0.003
R26605 D.n6091 D.n6090 0.003
R26606 D.n6105 D.n6104 0.003
R26607 D.n6119 D.n6118 0.003
R26608 D.n6133 D.n6132 0.003
R26609 D.n6147 D.n6146 0.003
R26610 D.n6161 D.n6160 0.003
R26611 D.n6175 D.n6174 0.003
R26612 D.n6189 D.n6188 0.003
R26613 D.n6213 D.n6212 0.003
R26614 D.n6229 D.n6228 0.003
R26615 D.n6243 D.n6242 0.003
R26616 D.n6257 D.n6256 0.003
R26617 D.n6271 D.n6270 0.003
R26618 D.n6285 D.n6284 0.003
R26619 D.n6299 D.n6298 0.003
R26620 D.n6313 D.n6312 0.003
R26621 D.n6327 D.n6326 0.003
R26622 D.n6341 D.n6340 0.003
R26623 D.n6355 D.n6354 0.003
R26624 D.n6369 D.n6368 0.003
R26625 D.n6383 D.n6382 0.003
R26626 D.n6397 D.n6396 0.003
R26627 D.n6411 D.n6410 0.003
R26628 D.n6425 D.n6424 0.003
R26629 D.n6439 D.n6438 0.003
R26630 D.n6453 D.n6452 0.003
R26631 D.n6467 D.n6466 0.003
R26632 D.n6481 D.n6480 0.003
R26633 D.n6505 D.n6504 0.003
R26634 D.n6521 D.n6520 0.003
R26635 D.n6535 D.n6534 0.003
R26636 D.n6549 D.n6548 0.003
R26637 D.n6563 D.n6562 0.003
R26638 D.n6577 D.n6576 0.003
R26639 D.n6591 D.n6590 0.003
R26640 D.n6605 D.n6604 0.003
R26641 D.n6619 D.n6618 0.003
R26642 D.n6633 D.n6632 0.003
R26643 D.n6647 D.n6646 0.003
R26644 D.n6661 D.n6660 0.003
R26645 D.n6675 D.n6674 0.003
R26646 D.n6689 D.n6688 0.003
R26647 D.n6703 D.n6702 0.003
R26648 D.n6717 D.n6716 0.003
R26649 D.n6731 D.n6730 0.003
R26650 D.n6745 D.n6744 0.003
R26651 D.n6769 D.n6768 0.003
R26652 D.n6785 D.n6784 0.003
R26653 D.n6799 D.n6798 0.003
R26654 D.n6813 D.n6812 0.003
R26655 D.n6827 D.n6826 0.003
R26656 D.n6841 D.n6840 0.003
R26657 D.n6855 D.n6854 0.003
R26658 D.n6869 D.n6868 0.003
R26659 D.n6883 D.n6882 0.003
R26660 D.n6897 D.n6896 0.003
R26661 D.n6911 D.n6910 0.003
R26662 D.n6925 D.n6924 0.003
R26663 D.n6939 D.n6938 0.003
R26664 D.n6953 D.n6952 0.003
R26665 D.n6967 D.n6966 0.003
R26666 D.n6981 D.n6980 0.003
R26667 D.n7005 D.n7004 0.003
R26668 D.n7021 D.n7020 0.003
R26669 D.n7035 D.n7034 0.003
R26670 D.n7049 D.n7048 0.003
R26671 D.n7063 D.n7062 0.003
R26672 D.n7077 D.n7076 0.003
R26673 D.n7091 D.n7090 0.003
R26674 D.n7105 D.n7104 0.003
R26675 D.n7119 D.n7118 0.003
R26676 D.n7133 D.n7132 0.003
R26677 D.n7147 D.n7146 0.003
R26678 D.n7161 D.n7160 0.003
R26679 D.n7175 D.n7174 0.003
R26680 D.n7189 D.n7188 0.003
R26681 D.n7213 D.n7212 0.003
R26682 D.n7229 D.n7228 0.003
R26683 D.n7243 D.n7242 0.003
R26684 D.n7257 D.n7256 0.003
R26685 D.n7271 D.n7270 0.003
R26686 D.n7285 D.n7284 0.003
R26687 D.n7299 D.n7298 0.003
R26688 D.n7313 D.n7312 0.003
R26689 D.n7327 D.n7326 0.003
R26690 D.n7341 D.n7340 0.003
R26691 D.n7355 D.n7354 0.003
R26692 D.n7369 D.n7368 0.003
R26693 D.n7393 D.n7392 0.003
R26694 D.n7409 D.n7408 0.003
R26695 D.n7423 D.n7422 0.003
R26696 D.n7437 D.n7436 0.003
R26697 D.n7451 D.n7450 0.003
R26698 D.n7465 D.n7464 0.003
R26699 D.n7479 D.n7478 0.003
R26700 D.n7493 D.n7492 0.003
R26701 D.n7507 D.n7506 0.003
R26702 D.n7521 D.n7520 0.003
R26703 D.n7545 D.n7544 0.003
R26704 D.n7561 D.n7560 0.003
R26705 D.n7575 D.n7574 0.003
R26706 D.n7589 D.n7588 0.003
R26707 D.n7603 D.n7602 0.003
R26708 D.n7617 D.n7616 0.003
R26709 D.n7631 D.n7630 0.003
R26710 D.n7645 D.n7644 0.003
R26711 D.n7669 D.n7668 0.003
R26712 D.n7685 D.n7684 0.003
R26713 D.n7699 D.n7698 0.003
R26714 D.n7713 D.n7712 0.003
R26715 D.n7727 D.n7726 0.003
R26716 D.n7741 D.n7740 0.003
R26717 D.n7764 D.n7763 0.003
R26718 D.n7780 D.n7779 0.003
R26719 D.n7794 D.n7793 0.003
R26720 D.n7810 D.n7808 0.003
R26721 D.n39 D.n38 0.003
R26722 D.n37 D.n36 0.003
R26723 D.n13643 D.n13642 0.003
R26724 D.n12720 D.n12719 0.003
R26725 D.n11871 D.n11870 0.003
R26726 D.n11108 D.n11107 0.003
R26727 D.n10425 D.n10424 0.003
R26728 D.n9822 D.n9821 0.003
R26729 D.n9293 D.n9292 0.003
R26730 D.n8850 D.n8849 0.003
R26731 D.n8487 D.n8486 0.003
R26732 D.n8198 D.n8197 0.003
R26733 D.n7995 D.n7994 0.003
R26734 D.n7832 D.n7824 0.003
R26735 D.n7962 D.n7954 0.003
R26736 D.n7842 D.n7834 0.003
R26737 D.n7952 D.n7939 0.003
R26738 D.n13212 D.n13204 0.003
R26739 D.n13222 D.n13214 0.003
R26740 D.n13232 D.n13224 0.003
R26741 D.n13242 D.n13234 0.003
R26742 D.n13252 D.n13244 0.003
R26743 D.n13262 D.n13254 0.003
R26744 D.n13272 D.n13264 0.003
R26745 D.n13282 D.n13274 0.003
R26746 D.n13292 D.n13284 0.003
R26747 D.n13302 D.n13294 0.003
R26748 D.n13312 D.n13304 0.003
R26749 D.n13322 D.n13314 0.003
R26750 D.n13332 D.n13324 0.003
R26751 D.n13342 D.n13334 0.003
R26752 D.n13352 D.n13344 0.003
R26753 D.n13362 D.n13354 0.003
R26754 D.n13372 D.n13364 0.003
R26755 D.n13382 D.n13374 0.003
R26756 D.n13392 D.n13384 0.003
R26757 D.n13402 D.n13394 0.003
R26758 D.n13412 D.n13404 0.003
R26759 D.n13422 D.n13414 0.003
R26760 D.n13432 D.n13424 0.003
R26761 D.n13442 D.n13434 0.003
R26762 D.n13452 D.n13444 0.003
R26763 D.n13462 D.n13454 0.003
R26764 D.n13472 D.n13464 0.003
R26765 D.n13482 D.n13474 0.003
R26766 D.n13492 D.n13484 0.003
R26767 D.n13502 D.n13494 0.003
R26768 D.n13512 D.n13504 0.003
R26769 D.n13522 D.n13514 0.003
R26770 D.n13532 D.n13524 0.003
R26771 D.n13542 D.n13534 0.003
R26772 D.n13552 D.n13544 0.003
R26773 D.n13562 D.n13554 0.003
R26774 D.n13572 D.n13564 0.003
R26775 D.n13582 D.n13574 0.003
R26776 D.n13592 D.n13584 0.003
R26777 D.n13602 D.n13594 0.003
R26778 D.n13612 D.n13604 0.003
R26779 D.n12329 D.n12321 0.003
R26780 D.n12339 D.n12331 0.003
R26781 D.n12349 D.n12341 0.003
R26782 D.n12359 D.n12351 0.003
R26783 D.n12369 D.n12361 0.003
R26784 D.n12379 D.n12371 0.003
R26785 D.n12389 D.n12381 0.003
R26786 D.n12399 D.n12391 0.003
R26787 D.n12409 D.n12401 0.003
R26788 D.n12419 D.n12411 0.003
R26789 D.n12429 D.n12421 0.003
R26790 D.n12439 D.n12431 0.003
R26791 D.n12449 D.n12441 0.003
R26792 D.n12459 D.n12451 0.003
R26793 D.n12469 D.n12461 0.003
R26794 D.n12479 D.n12471 0.003
R26795 D.n12489 D.n12481 0.003
R26796 D.n12499 D.n12491 0.003
R26797 D.n12509 D.n12501 0.003
R26798 D.n12519 D.n12511 0.003
R26799 D.n12529 D.n12521 0.003
R26800 D.n12539 D.n12531 0.003
R26801 D.n12549 D.n12541 0.003
R26802 D.n12559 D.n12551 0.003
R26803 D.n12569 D.n12561 0.003
R26804 D.n12579 D.n12571 0.003
R26805 D.n12589 D.n12581 0.003
R26806 D.n12599 D.n12591 0.003
R26807 D.n12609 D.n12601 0.003
R26808 D.n12619 D.n12611 0.003
R26809 D.n12629 D.n12621 0.003
R26810 D.n12639 D.n12631 0.003
R26811 D.n12649 D.n12641 0.003
R26812 D.n12659 D.n12651 0.003
R26813 D.n12669 D.n12661 0.003
R26814 D.n12679 D.n12671 0.003
R26815 D.n12689 D.n12681 0.003
R26816 D.n11520 D.n11512 0.003
R26817 D.n11530 D.n11522 0.003
R26818 D.n11540 D.n11532 0.003
R26819 D.n11550 D.n11542 0.003
R26820 D.n11560 D.n11552 0.003
R26821 D.n11570 D.n11562 0.003
R26822 D.n11580 D.n11572 0.003
R26823 D.n11590 D.n11582 0.003
R26824 D.n11600 D.n11592 0.003
R26825 D.n11610 D.n11602 0.003
R26826 D.n11620 D.n11612 0.003
R26827 D.n11630 D.n11622 0.003
R26828 D.n11640 D.n11632 0.003
R26829 D.n11650 D.n11642 0.003
R26830 D.n11660 D.n11652 0.003
R26831 D.n11670 D.n11662 0.003
R26832 D.n11680 D.n11672 0.003
R26833 D.n11690 D.n11682 0.003
R26834 D.n11700 D.n11692 0.003
R26835 D.n11710 D.n11702 0.003
R26836 D.n11720 D.n11712 0.003
R26837 D.n11730 D.n11722 0.003
R26838 D.n11740 D.n11732 0.003
R26839 D.n11750 D.n11742 0.003
R26840 D.n11760 D.n11752 0.003
R26841 D.n11770 D.n11762 0.003
R26842 D.n11780 D.n11772 0.003
R26843 D.n11790 D.n11782 0.003
R26844 D.n11800 D.n11792 0.003
R26845 D.n11810 D.n11802 0.003
R26846 D.n11820 D.n11812 0.003
R26847 D.n11830 D.n11822 0.003
R26848 D.n11840 D.n11832 0.003
R26849 D.n10797 D.n10789 0.003
R26850 D.n10807 D.n10799 0.003
R26851 D.n10817 D.n10809 0.003
R26852 D.n10827 D.n10819 0.003
R26853 D.n10837 D.n10829 0.003
R26854 D.n10847 D.n10839 0.003
R26855 D.n10857 D.n10849 0.003
R26856 D.n10867 D.n10859 0.003
R26857 D.n10877 D.n10869 0.003
R26858 D.n10887 D.n10879 0.003
R26859 D.n10897 D.n10889 0.003
R26860 D.n10907 D.n10899 0.003
R26861 D.n10917 D.n10909 0.003
R26862 D.n10927 D.n10919 0.003
R26863 D.n10937 D.n10929 0.003
R26864 D.n10947 D.n10939 0.003
R26865 D.n10957 D.n10949 0.003
R26866 D.n10967 D.n10959 0.003
R26867 D.n10977 D.n10969 0.003
R26868 D.n10987 D.n10979 0.003
R26869 D.n10997 D.n10989 0.003
R26870 D.n11007 D.n10999 0.003
R26871 D.n11017 D.n11009 0.003
R26872 D.n11027 D.n11019 0.003
R26873 D.n11037 D.n11029 0.003
R26874 D.n11047 D.n11039 0.003
R26875 D.n11057 D.n11049 0.003
R26876 D.n11067 D.n11059 0.003
R26877 D.n11077 D.n11069 0.003
R26878 D.n10154 D.n10146 0.003
R26879 D.n10164 D.n10156 0.003
R26880 D.n10174 D.n10166 0.003
R26881 D.n10184 D.n10176 0.003
R26882 D.n10194 D.n10186 0.003
R26883 D.n10204 D.n10196 0.003
R26884 D.n10214 D.n10206 0.003
R26885 D.n10224 D.n10216 0.003
R26886 D.n10234 D.n10226 0.003
R26887 D.n10244 D.n10236 0.003
R26888 D.n10254 D.n10246 0.003
R26889 D.n10264 D.n10256 0.003
R26890 D.n10274 D.n10266 0.003
R26891 D.n10284 D.n10276 0.003
R26892 D.n10294 D.n10286 0.003
R26893 D.n10304 D.n10296 0.003
R26894 D.n10314 D.n10306 0.003
R26895 D.n10324 D.n10316 0.003
R26896 D.n10334 D.n10326 0.003
R26897 D.n10344 D.n10336 0.003
R26898 D.n10354 D.n10346 0.003
R26899 D.n10364 D.n10356 0.003
R26900 D.n10374 D.n10366 0.003
R26901 D.n10384 D.n10376 0.003
R26902 D.n10394 D.n10386 0.003
R26903 D.n9591 D.n9583 0.003
R26904 D.n9601 D.n9593 0.003
R26905 D.n9611 D.n9603 0.003
R26906 D.n9621 D.n9613 0.003
R26907 D.n9631 D.n9623 0.003
R26908 D.n9641 D.n9633 0.003
R26909 D.n9651 D.n9643 0.003
R26910 D.n9661 D.n9653 0.003
R26911 D.n9671 D.n9663 0.003
R26912 D.n9681 D.n9673 0.003
R26913 D.n9691 D.n9683 0.003
R26914 D.n9701 D.n9693 0.003
R26915 D.n9711 D.n9703 0.003
R26916 D.n9721 D.n9713 0.003
R26917 D.n9731 D.n9723 0.003
R26918 D.n9741 D.n9733 0.003
R26919 D.n9751 D.n9743 0.003
R26920 D.n9761 D.n9753 0.003
R26921 D.n9771 D.n9763 0.003
R26922 D.n9781 D.n9773 0.003
R26923 D.n9791 D.n9783 0.003
R26924 D.n9102 D.n9094 0.003
R26925 D.n9112 D.n9104 0.003
R26926 D.n9122 D.n9114 0.003
R26927 D.n9132 D.n9124 0.003
R26928 D.n9142 D.n9134 0.003
R26929 D.n9152 D.n9144 0.003
R26930 D.n9162 D.n9154 0.003
R26931 D.n9172 D.n9164 0.003
R26932 D.n9182 D.n9174 0.003
R26933 D.n9192 D.n9184 0.003
R26934 D.n9202 D.n9194 0.003
R26935 D.n9212 D.n9204 0.003
R26936 D.n9222 D.n9214 0.003
R26937 D.n9232 D.n9224 0.003
R26938 D.n9242 D.n9234 0.003
R26939 D.n9252 D.n9244 0.003
R26940 D.n9262 D.n9254 0.003
R26941 D.n8699 D.n8691 0.003
R26942 D.n8709 D.n8701 0.003
R26943 D.n8719 D.n8711 0.003
R26944 D.n8729 D.n8721 0.003
R26945 D.n8739 D.n8731 0.003
R26946 D.n8749 D.n8741 0.003
R26947 D.n8759 D.n8751 0.003
R26948 D.n8769 D.n8761 0.003
R26949 D.n8779 D.n8771 0.003
R26950 D.n8789 D.n8781 0.003
R26951 D.n8799 D.n8791 0.003
R26952 D.n8809 D.n8801 0.003
R26953 D.n8819 D.n8811 0.003
R26954 D.n8376 D.n8368 0.003
R26955 D.n8386 D.n8378 0.003
R26956 D.n8396 D.n8388 0.003
R26957 D.n8406 D.n8398 0.003
R26958 D.n8416 D.n8408 0.003
R26959 D.n8426 D.n8418 0.003
R26960 D.n8436 D.n8428 0.003
R26961 D.n8446 D.n8438 0.003
R26962 D.n8456 D.n8448 0.003
R26963 D.n8127 D.n8119 0.003
R26964 D.n8137 D.n8129 0.003
R26965 D.n8147 D.n8139 0.003
R26966 D.n8157 D.n8149 0.003
R26967 D.n8167 D.n8159 0.003
R26968 D.n13202 D.n13189 0.003
R26969 D.n12319 D.n12306 0.003
R26970 D.n11510 D.n11499 0.003
R26971 D.n10787 D.n10776 0.003
R26972 D.n10144 D.n10131 0.003
R26973 D.n9581 D.n9568 0.003
R26974 D.n9092 D.n9081 0.003
R26975 D.n8689 D.n8676 0.003
R26976 D.n8366 D.n8353 0.003
R26977 D.n8117 D.n8106 0.003
R26978 D.n13668 D.n13667 0.002
R26979 D.n21 D.n20 0.002
R26980 D.n19 D.n18 0.002
R26981 D.n7984 D.n7983 0.001
R26982 D.n13655 D.n13654 0.001
R26983 D.n13675 D.n13674 0.001
R26984 D.n13620 D.n13619 0.001
R26985 D.n13632 D.n13631 0.001
R26986 D.n13638 D.n13637 0.001
R26987 D.n12732 D.n12731 0.001
R26988 D.n12748 D.n12747 0.001
R26989 D.n12697 D.n12696 0.001
R26990 D.n12709 D.n12708 0.001
R26991 D.n12715 D.n12714 0.001
R26992 D.n11883 D.n11882 0.001
R26993 D.n11899 D.n11898 0.001
R26994 D.n11848 D.n11847 0.001
R26995 D.n11860 D.n11859 0.001
R26996 D.n11866 D.n11865 0.001
R26997 D.n11120 D.n11119 0.001
R26998 D.n11136 D.n11135 0.001
R26999 D.n11085 D.n11084 0.001
R27000 D.n11097 D.n11096 0.001
R27001 D.n11103 D.n11102 0.001
R27002 D.n10437 D.n10436 0.001
R27003 D.n10453 D.n10452 0.001
R27004 D.n10402 D.n10401 0.001
R27005 D.n10414 D.n10413 0.001
R27006 D.n10420 D.n10419 0.001
R27007 D.n9834 D.n9833 0.001
R27008 D.n9850 D.n9849 0.001
R27009 D.n9799 D.n9798 0.001
R27010 D.n9811 D.n9810 0.001
R27011 D.n9817 D.n9816 0.001
R27012 D.n9305 D.n9304 0.001
R27013 D.n9321 D.n9320 0.001
R27014 D.n9270 D.n9269 0.001
R27015 D.n9282 D.n9281 0.001
R27016 D.n9288 D.n9287 0.001
R27017 D.n8862 D.n8861 0.001
R27018 D.n8878 D.n8877 0.001
R27019 D.n8827 D.n8826 0.001
R27020 D.n8839 D.n8838 0.001
R27021 D.n8845 D.n8844 0.001
R27022 D.n8499 D.n8498 0.001
R27023 D.n8515 D.n8514 0.001
R27024 D.n8464 D.n8463 0.001
R27025 D.n8476 D.n8475 0.001
R27026 D.n8482 D.n8481 0.001
R27027 D.n8210 D.n8209 0.001
R27028 D.n8226 D.n8225 0.001
R27029 D.n8175 D.n8174 0.001
R27030 D.n8187 D.n8186 0.001
R27031 D.n8193 D.n8192 0.001
R27032 D.n8007 D.n8006 0.001
R27033 D.n8023 D.n8022 0.001
R27034 D.n7990 D.n7989 0.001
R27035 D.n7970 D.n7969 0.001
R27036 D.n507 D.n506 0.001
R27037 D.n43 D.n42 0.001
R27038 D.n15 D.n14 0.001
R27039 D.n25 D.n24 0.001
R27040 D.n7850 D.n7849 0.001
R27041 D.n14141 D.n13679 0.001
R27042 D.n13168 D.n12752 0.001
R27043 D.n12285 D.n11903 0.001
R27044 D.n11482 D.n11140 0.001
R27045 D.n10759 D.n10457 0.001
R27046 D.n10110 D.n9854 0.001
R27047 D.n9547 D.n9325 0.001
R27048 D.n9064 D.n8882 0.001
R27049 D.n8655 D.n8519 0.001
R27050 D.n8332 D.n8230 0.001
R27051 D.n8089 D.n8027 0.001
R27052 D.n7921 D.n7902 0.001
R27053 D.n456 D.n453 0.001
R27054 D.n457 D.n444 0.001
R27055 D.n458 D.n435 0.001
R27056 D.n459 D.n426 0.001
R27057 D.n460 D.n417 0.001
R27058 D.n461 D.n408 0.001
R27059 D.n462 D.n399 0.001
R27060 D.n463 D.n390 0.001
R27061 D.n464 D.n381 0.001
R27062 D.n465 D.n372 0.001
R27063 D.n466 D.n363 0.001
R27064 D.n467 D.n354 0.001
R27065 D.n468 D.n345 0.001
R27066 D.n469 D.n336 0.001
R27067 D.n470 D.n327 0.001
R27068 D.n471 D.n318 0.001
R27069 D.n472 D.n309 0.001
R27070 D.n473 D.n300 0.001
R27071 D.n474 D.n291 0.001
R27072 D.n475 D.n282 0.001
R27073 D.n476 D.n273 0.001
R27074 D.n477 D.n264 0.001
R27075 D.n478 D.n255 0.001
R27076 D.n479 D.n246 0.001
R27077 D.n480 D.n237 0.001
R27078 D.n481 D.n228 0.001
R27079 D.n482 D.n219 0.001
R27080 D.n483 D.n210 0.001
R27081 D.n484 D.n201 0.001
R27082 D.n485 D.n192 0.001
R27083 D.n486 D.n183 0.001
R27084 D.n487 D.n174 0.001
R27085 D.n488 D.n165 0.001
R27086 D.n489 D.n156 0.001
R27087 D.n490 D.n147 0.001
R27088 D.n491 D.n138 0.001
R27089 D.n492 D.n129 0.001
R27090 D.n493 D.n120 0.001
R27091 D.n494 D.n111 0.001
R27092 D.n495 D.n102 0.001
R27093 D.n496 D.n93 0.001
R27094 D.n497 D.n84 0.001
R27095 D.n498 D.n75 0.001
R27096 D.n499 D.n66 0.001
R27097 D.n500 D.n57 0.001
R27098 D.n501 D.n47 0.001
R27099 D.n14097 D.n14081 0.001
R27100 D.n14098 D.n14067 0.001
R27101 D.n14099 D.n14058 0.001
R27102 D.n14100 D.n14049 0.001
R27103 D.n14101 D.n14040 0.001
R27104 D.n14102 D.n14031 0.001
R27105 D.n14103 D.n14022 0.001
R27106 D.n14104 D.n14013 0.001
R27107 D.n14105 D.n14004 0.001
R27108 D.n14106 D.n13995 0.001
R27109 D.n14107 D.n13986 0.001
R27110 D.n14108 D.n13977 0.001
R27111 D.n14109 D.n13968 0.001
R27112 D.n14110 D.n13959 0.001
R27113 D.n14111 D.n13950 0.001
R27114 D.n14112 D.n13941 0.001
R27115 D.n14113 D.n13932 0.001
R27116 D.n14114 D.n13923 0.001
R27117 D.n14115 D.n13914 0.001
R27118 D.n14116 D.n13905 0.001
R27119 D.n14117 D.n13896 0.001
R27120 D.n14118 D.n13887 0.001
R27121 D.n14119 D.n13878 0.001
R27122 D.n14120 D.n13869 0.001
R27123 D.n14121 D.n13860 0.001
R27124 D.n14122 D.n13851 0.001
R27125 D.n14123 D.n13842 0.001
R27126 D.n14124 D.n13833 0.001
R27127 D.n14125 D.n13824 0.001
R27128 D.n14126 D.n13815 0.001
R27129 D.n14127 D.n13806 0.001
R27130 D.n14128 D.n13797 0.001
R27131 D.n14129 D.n13788 0.001
R27132 D.n14130 D.n13779 0.001
R27133 D.n14131 D.n13770 0.001
R27134 D.n14132 D.n13761 0.001
R27135 D.n14133 D.n13752 0.001
R27136 D.n14134 D.n13743 0.001
R27137 D.n14135 D.n13734 0.001
R27138 D.n14136 D.n13725 0.001
R27139 D.n14137 D.n13716 0.001
R27140 D.n14138 D.n13707 0.001
R27141 D.n14139 D.n13698 0.001
R27142 D.n14140 D.n13689 0.001
R27143 D.n13128 D.n13117 0.001
R27144 D.n13129 D.n13104 0.001
R27145 D.n13130 D.n13095 0.001
R27146 D.n13131 D.n13086 0.001
R27147 D.n13132 D.n13077 0.001
R27148 D.n13133 D.n13068 0.001
R27149 D.n13134 D.n13059 0.001
R27150 D.n13135 D.n13050 0.001
R27151 D.n13136 D.n13041 0.001
R27152 D.n13137 D.n13032 0.001
R27153 D.n13138 D.n13023 0.001
R27154 D.n13139 D.n13014 0.001
R27155 D.n13140 D.n13005 0.001
R27156 D.n13141 D.n12996 0.001
R27157 D.n13142 D.n12987 0.001
R27158 D.n13143 D.n12978 0.001
R27159 D.n13144 D.n12969 0.001
R27160 D.n13145 D.n12960 0.001
R27161 D.n13146 D.n12951 0.001
R27162 D.n13147 D.n12942 0.001
R27163 D.n13148 D.n12933 0.001
R27164 D.n13149 D.n12924 0.001
R27165 D.n13150 D.n12915 0.001
R27166 D.n13151 D.n12906 0.001
R27167 D.n13152 D.n12897 0.001
R27168 D.n13153 D.n12888 0.001
R27169 D.n13154 D.n12879 0.001
R27170 D.n13155 D.n12870 0.001
R27171 D.n13156 D.n12861 0.001
R27172 D.n13157 D.n12852 0.001
R27173 D.n13158 D.n12843 0.001
R27174 D.n13159 D.n12834 0.001
R27175 D.n13160 D.n12825 0.001
R27176 D.n13161 D.n12816 0.001
R27177 D.n13162 D.n12807 0.001
R27178 D.n13163 D.n12798 0.001
R27179 D.n13164 D.n12789 0.001
R27180 D.n13165 D.n12780 0.001
R27181 D.n13166 D.n12771 0.001
R27182 D.n13167 D.n12762 0.001
R27183 D.n12249 D.n12232 0.001
R27184 D.n12250 D.n12219 0.001
R27185 D.n12251 D.n12210 0.001
R27186 D.n12252 D.n12201 0.001
R27187 D.n12253 D.n12192 0.001
R27188 D.n12254 D.n12183 0.001
R27189 D.n12255 D.n12174 0.001
R27190 D.n12256 D.n12165 0.001
R27191 D.n12257 D.n12156 0.001
R27192 D.n12258 D.n12147 0.001
R27193 D.n12259 D.n12138 0.001
R27194 D.n12260 D.n12129 0.001
R27195 D.n12261 D.n12120 0.001
R27196 D.n12262 D.n12111 0.001
R27197 D.n12263 D.n12102 0.001
R27198 D.n12264 D.n12093 0.001
R27199 D.n12265 D.n12084 0.001
R27200 D.n12266 D.n12075 0.001
R27201 D.n12267 D.n12066 0.001
R27202 D.n12268 D.n12057 0.001
R27203 D.n12269 D.n12048 0.001
R27204 D.n12270 D.n12039 0.001
R27205 D.n12271 D.n12030 0.001
R27206 D.n12272 D.n12021 0.001
R27207 D.n12273 D.n12012 0.001
R27208 D.n12274 D.n12003 0.001
R27209 D.n12275 D.n11994 0.001
R27210 D.n12276 D.n11985 0.001
R27211 D.n12277 D.n11976 0.001
R27212 D.n12278 D.n11967 0.001
R27213 D.n12279 D.n11958 0.001
R27214 D.n12280 D.n11949 0.001
R27215 D.n12281 D.n11940 0.001
R27216 D.n12282 D.n11931 0.001
R27217 D.n12283 D.n11922 0.001
R27218 D.n12284 D.n11913 0.001
R27219 D.n11450 D.n11433 0.001
R27220 D.n11451 D.n11420 0.001
R27221 D.n11452 D.n11411 0.001
R27222 D.n11453 D.n11402 0.001
R27223 D.n11454 D.n11393 0.001
R27224 D.n11455 D.n11384 0.001
R27225 D.n11456 D.n11375 0.001
R27226 D.n11457 D.n11366 0.001
R27227 D.n11458 D.n11357 0.001
R27228 D.n11459 D.n11348 0.001
R27229 D.n11460 D.n11339 0.001
R27230 D.n11461 D.n11330 0.001
R27231 D.n11462 D.n11321 0.001
R27232 D.n11463 D.n11312 0.001
R27233 D.n11464 D.n11303 0.001
R27234 D.n11465 D.n11294 0.001
R27235 D.n11466 D.n11285 0.001
R27236 D.n11467 D.n11276 0.001
R27237 D.n11468 D.n11267 0.001
R27238 D.n11469 D.n11258 0.001
R27239 D.n11470 D.n11249 0.001
R27240 D.n11471 D.n11240 0.001
R27241 D.n11472 D.n11231 0.001
R27242 D.n11473 D.n11222 0.001
R27243 D.n11474 D.n11213 0.001
R27244 D.n11475 D.n11204 0.001
R27245 D.n11476 D.n11195 0.001
R27246 D.n11477 D.n11186 0.001
R27247 D.n11478 D.n11177 0.001
R27248 D.n11479 D.n11168 0.001
R27249 D.n11480 D.n11159 0.001
R27250 D.n11481 D.n11150 0.001
R27251 D.n10731 D.n10714 0.001
R27252 D.n10732 D.n10701 0.001
R27253 D.n10733 D.n10692 0.001
R27254 D.n10734 D.n10683 0.001
R27255 D.n10735 D.n10674 0.001
R27256 D.n10736 D.n10665 0.001
R27257 D.n10737 D.n10656 0.001
R27258 D.n10738 D.n10647 0.001
R27259 D.n10739 D.n10638 0.001
R27260 D.n10740 D.n10629 0.001
R27261 D.n10741 D.n10620 0.001
R27262 D.n10742 D.n10611 0.001
R27263 D.n10743 D.n10602 0.001
R27264 D.n10744 D.n10593 0.001
R27265 D.n10745 D.n10584 0.001
R27266 D.n10746 D.n10575 0.001
R27267 D.n10747 D.n10566 0.001
R27268 D.n10748 D.n10557 0.001
R27269 D.n10749 D.n10548 0.001
R27270 D.n10750 D.n10539 0.001
R27271 D.n10751 D.n10530 0.001
R27272 D.n10752 D.n10521 0.001
R27273 D.n10753 D.n10512 0.001
R27274 D.n10754 D.n10503 0.001
R27275 D.n10755 D.n10494 0.001
R27276 D.n10756 D.n10485 0.001
R27277 D.n10757 D.n10476 0.001
R27278 D.n10758 D.n10467 0.001
R27279 D.n10086 D.n10075 0.001
R27280 D.n10087 D.n10062 0.001
R27281 D.n10088 D.n10053 0.001
R27282 D.n10089 D.n10044 0.001
R27283 D.n10090 D.n10035 0.001
R27284 D.n10091 D.n10026 0.001
R27285 D.n10092 D.n10017 0.001
R27286 D.n10093 D.n10008 0.001
R27287 D.n10094 D.n9999 0.001
R27288 D.n10095 D.n9990 0.001
R27289 D.n10096 D.n9981 0.001
R27290 D.n10097 D.n9972 0.001
R27291 D.n10098 D.n9963 0.001
R27292 D.n10099 D.n9954 0.001
R27293 D.n10100 D.n9945 0.001
R27294 D.n10101 D.n9936 0.001
R27295 D.n10102 D.n9927 0.001
R27296 D.n10103 D.n9918 0.001
R27297 D.n10104 D.n9909 0.001
R27298 D.n10105 D.n9900 0.001
R27299 D.n10106 D.n9891 0.001
R27300 D.n10107 D.n9882 0.001
R27301 D.n10108 D.n9873 0.001
R27302 D.n10109 D.n9864 0.001
R27303 D.n9527 D.n9510 0.001
R27304 D.n9528 D.n9497 0.001
R27305 D.n9529 D.n9488 0.001
R27306 D.n9530 D.n9479 0.001
R27307 D.n9531 D.n9470 0.001
R27308 D.n9532 D.n9461 0.001
R27309 D.n9533 D.n9452 0.001
R27310 D.n9534 D.n9443 0.001
R27311 D.n9535 D.n9434 0.001
R27312 D.n9536 D.n9425 0.001
R27313 D.n9537 D.n9416 0.001
R27314 D.n9538 D.n9407 0.001
R27315 D.n9539 D.n9398 0.001
R27316 D.n9540 D.n9389 0.001
R27317 D.n9541 D.n9380 0.001
R27318 D.n9542 D.n9371 0.001
R27319 D.n9543 D.n9362 0.001
R27320 D.n9544 D.n9353 0.001
R27321 D.n9545 D.n9344 0.001
R27322 D.n9546 D.n9335 0.001
R27323 D.n9048 D.n9031 0.001
R27324 D.n9049 D.n9018 0.001
R27325 D.n9050 D.n9009 0.001
R27326 D.n9051 D.n9000 0.001
R27327 D.n9052 D.n8991 0.001
R27328 D.n9053 D.n8982 0.001
R27329 D.n9054 D.n8973 0.001
R27330 D.n9055 D.n8964 0.001
R27331 D.n9056 D.n8955 0.001
R27332 D.n9057 D.n8946 0.001
R27333 D.n9058 D.n8937 0.001
R27334 D.n9059 D.n8928 0.001
R27335 D.n9060 D.n8919 0.001
R27336 D.n9061 D.n8910 0.001
R27337 D.n9062 D.n8901 0.001
R27338 D.n9063 D.n8892 0.001
R27339 D.n8643 D.n8632 0.001
R27340 D.n8644 D.n8619 0.001
R27341 D.n8645 D.n8610 0.001
R27342 D.n8646 D.n8601 0.001
R27343 D.n8647 D.n8592 0.001
R27344 D.n8648 D.n8583 0.001
R27345 D.n8649 D.n8574 0.001
R27346 D.n8650 D.n8565 0.001
R27347 D.n8651 D.n8556 0.001
R27348 D.n8652 D.n8547 0.001
R27349 D.n8653 D.n8538 0.001
R27350 D.n8654 D.n8529 0.001
R27351 D.n8324 D.n8307 0.001
R27352 D.n8325 D.n8294 0.001
R27353 D.n8326 D.n8285 0.001
R27354 D.n8327 D.n8276 0.001
R27355 D.n8328 D.n8267 0.001
R27356 D.n8329 D.n8258 0.001
R27357 D.n8330 D.n8249 0.001
R27358 D.n8331 D.n8240 0.001
R27359 D.n8085 D.n8068 0.001
R27360 D.n8086 D.n8055 0.001
R27361 D.n8087 D.n8046 0.001
R27362 D.n8088 D.n8037 0.001
R27363 D.n1138 D.n1137 0.001
R27364 D.n1124 D.n1123 0.001
R27365 D.n1110 D.n1109 0.001
R27366 D.n1096 D.n1095 0.001
R27367 D.n1082 D.n1081 0.001
R27368 D.n1068 D.n1067 0.001
R27369 D.n1054 D.n1053 0.001
R27370 D.n1040 D.n1039 0.001
R27371 D.n1026 D.n1025 0.001
R27372 D.n1012 D.n1011 0.001
R27373 D.n998 D.n997 0.001
R27374 D.n984 D.n983 0.001
R27375 D.n970 D.n969 0.001
R27376 D.n956 D.n955 0.001
R27377 D.n942 D.n941 0.001
R27378 D.n928 D.n927 0.001
R27379 D.n914 D.n913 0.001
R27380 D.n900 D.n899 0.001
R27381 D.n886 D.n885 0.001
R27382 D.n872 D.n871 0.001
R27383 D.n858 D.n857 0.001
R27384 D.n844 D.n843 0.001
R27385 D.n830 D.n829 0.001
R27386 D.n816 D.n815 0.001
R27387 D.n802 D.n801 0.001
R27388 D.n788 D.n787 0.001
R27389 D.n774 D.n773 0.001
R27390 D.n760 D.n759 0.001
R27391 D.n746 D.n745 0.001
R27392 D.n732 D.n731 0.001
R27393 D.n718 D.n717 0.001
R27394 D.n704 D.n703 0.001
R27395 D.n690 D.n689 0.001
R27396 D.n676 D.n675 0.001
R27397 D.n662 D.n661 0.001
R27398 D.n648 D.n647 0.001
R27399 D.n634 D.n633 0.001
R27400 D.n620 D.n619 0.001
R27401 D.n606 D.n605 0.001
R27402 D.n592 D.n591 0.001
R27403 D.n578 D.n577 0.001
R27404 D.n564 D.n563 0.001
R27405 D.n550 D.n549 0.001
R27406 D.n536 D.n535 0.001
R27407 D.n1737 D.n1736 0.001
R27408 D.n1723 D.n1722 0.001
R27409 D.n1709 D.n1708 0.001
R27410 D.n1695 D.n1694 0.001
R27411 D.n1681 D.n1680 0.001
R27412 D.n1667 D.n1666 0.001
R27413 D.n1653 D.n1652 0.001
R27414 D.n1639 D.n1638 0.001
R27415 D.n1625 D.n1624 0.001
R27416 D.n1611 D.n1610 0.001
R27417 D.n1597 D.n1596 0.001
R27418 D.n1583 D.n1582 0.001
R27419 D.n1569 D.n1568 0.001
R27420 D.n1555 D.n1554 0.001
R27421 D.n1541 D.n1540 0.001
R27422 D.n1527 D.n1526 0.001
R27423 D.n1513 D.n1512 0.001
R27424 D.n1499 D.n1498 0.001
R27425 D.n1485 D.n1484 0.001
R27426 D.n1471 D.n1470 0.001
R27427 D.n1457 D.n1456 0.001
R27428 D.n1443 D.n1442 0.001
R27429 D.n1429 D.n1428 0.001
R27430 D.n1415 D.n1414 0.001
R27431 D.n1401 D.n1400 0.001
R27432 D.n1387 D.n1386 0.001
R27433 D.n1373 D.n1372 0.001
R27434 D.n1359 D.n1358 0.001
R27435 D.n1345 D.n1344 0.001
R27436 D.n1331 D.n1330 0.001
R27437 D.n1317 D.n1316 0.001
R27438 D.n1303 D.n1302 0.001
R27439 D.n1289 D.n1288 0.001
R27440 D.n1275 D.n1274 0.001
R27441 D.n1261 D.n1260 0.001
R27442 D.n1247 D.n1246 0.001
R27443 D.n1233 D.n1232 0.001
R27444 D.n1219 D.n1218 0.001
R27445 D.n1205 D.n1204 0.001
R27446 D.n1191 D.n1190 0.001
R27447 D.n1177 D.n1176 0.001
R27448 D.n1163 D.n1162 0.001
R27449 D.n2308 D.n2307 0.001
R27450 D.n2294 D.n2293 0.001
R27451 D.n2280 D.n2279 0.001
R27452 D.n2266 D.n2265 0.001
R27453 D.n2252 D.n2251 0.001
R27454 D.n2238 D.n2237 0.001
R27455 D.n2224 D.n2223 0.001
R27456 D.n2210 D.n2209 0.001
R27457 D.n2196 D.n2195 0.001
R27458 D.n2182 D.n2181 0.001
R27459 D.n2168 D.n2167 0.001
R27460 D.n2154 D.n2153 0.001
R27461 D.n2140 D.n2139 0.001
R27462 D.n2126 D.n2125 0.001
R27463 D.n2112 D.n2111 0.001
R27464 D.n2098 D.n2097 0.001
R27465 D.n2084 D.n2083 0.001
R27466 D.n2070 D.n2069 0.001
R27467 D.n2056 D.n2055 0.001
R27468 D.n2042 D.n2041 0.001
R27469 D.n2028 D.n2027 0.001
R27470 D.n2014 D.n2013 0.001
R27471 D.n2000 D.n1999 0.001
R27472 D.n1986 D.n1985 0.001
R27473 D.n1972 D.n1971 0.001
R27474 D.n1958 D.n1957 0.001
R27475 D.n1944 D.n1943 0.001
R27476 D.n1930 D.n1929 0.001
R27477 D.n1916 D.n1915 0.001
R27478 D.n1902 D.n1901 0.001
R27479 D.n1888 D.n1887 0.001
R27480 D.n1874 D.n1873 0.001
R27481 D.n1860 D.n1859 0.001
R27482 D.n1846 D.n1845 0.001
R27483 D.n1832 D.n1831 0.001
R27484 D.n1818 D.n1817 0.001
R27485 D.n1804 D.n1803 0.001
R27486 D.n1790 D.n1789 0.001
R27487 D.n1776 D.n1775 0.001
R27488 D.n1762 D.n1761 0.001
R27489 D.n2851 D.n2850 0.001
R27490 D.n2837 D.n2836 0.001
R27491 D.n2823 D.n2822 0.001
R27492 D.n2809 D.n2808 0.001
R27493 D.n2795 D.n2794 0.001
R27494 D.n2781 D.n2780 0.001
R27495 D.n2767 D.n2766 0.001
R27496 D.n2753 D.n2752 0.001
R27497 D.n2739 D.n2738 0.001
R27498 D.n2725 D.n2724 0.001
R27499 D.n2711 D.n2710 0.001
R27500 D.n2697 D.n2696 0.001
R27501 D.n2683 D.n2682 0.001
R27502 D.n2669 D.n2668 0.001
R27503 D.n2655 D.n2654 0.001
R27504 D.n2641 D.n2640 0.001
R27505 D.n2627 D.n2626 0.001
R27506 D.n2613 D.n2612 0.001
R27507 D.n2599 D.n2598 0.001
R27508 D.n2585 D.n2584 0.001
R27509 D.n2571 D.n2570 0.001
R27510 D.n2557 D.n2556 0.001
R27511 D.n2543 D.n2542 0.001
R27512 D.n2529 D.n2528 0.001
R27513 D.n2515 D.n2514 0.001
R27514 D.n2501 D.n2500 0.001
R27515 D.n2487 D.n2486 0.001
R27516 D.n2473 D.n2472 0.001
R27517 D.n2459 D.n2458 0.001
R27518 D.n2445 D.n2444 0.001
R27519 D.n2431 D.n2430 0.001
R27520 D.n2417 D.n2416 0.001
R27521 D.n2403 D.n2402 0.001
R27522 D.n2389 D.n2388 0.001
R27523 D.n2375 D.n2374 0.001
R27524 D.n2361 D.n2360 0.001
R27525 D.n2347 D.n2346 0.001
R27526 D.n2333 D.n2332 0.001
R27527 D.n3366 D.n3365 0.001
R27528 D.n3352 D.n3351 0.001
R27529 D.n3338 D.n3337 0.001
R27530 D.n3324 D.n3323 0.001
R27531 D.n3310 D.n3309 0.001
R27532 D.n3296 D.n3295 0.001
R27533 D.n3282 D.n3281 0.001
R27534 D.n3268 D.n3267 0.001
R27535 D.n3254 D.n3253 0.001
R27536 D.n3240 D.n3239 0.001
R27537 D.n3226 D.n3225 0.001
R27538 D.n3212 D.n3211 0.001
R27539 D.n3198 D.n3197 0.001
R27540 D.n3184 D.n3183 0.001
R27541 D.n3170 D.n3169 0.001
R27542 D.n3156 D.n3155 0.001
R27543 D.n3142 D.n3141 0.001
R27544 D.n3128 D.n3127 0.001
R27545 D.n3114 D.n3113 0.001
R27546 D.n3100 D.n3099 0.001
R27547 D.n3086 D.n3085 0.001
R27548 D.n3072 D.n3071 0.001
R27549 D.n3058 D.n3057 0.001
R27550 D.n3044 D.n3043 0.001
R27551 D.n3030 D.n3029 0.001
R27552 D.n3016 D.n3015 0.001
R27553 D.n3002 D.n3001 0.001
R27554 D.n2988 D.n2987 0.001
R27555 D.n2974 D.n2973 0.001
R27556 D.n2960 D.n2959 0.001
R27557 D.n2946 D.n2945 0.001
R27558 D.n2932 D.n2931 0.001
R27559 D.n2918 D.n2917 0.001
R27560 D.n2904 D.n2903 0.001
R27561 D.n2890 D.n2889 0.001
R27562 D.n2876 D.n2875 0.001
R27563 D.n3854 D.n3853 0.001
R27564 D.n3840 D.n3839 0.001
R27565 D.n3826 D.n3825 0.001
R27566 D.n3812 D.n3811 0.001
R27567 D.n3798 D.n3797 0.001
R27568 D.n3784 D.n3783 0.001
R27569 D.n3770 D.n3769 0.001
R27570 D.n3756 D.n3755 0.001
R27571 D.n3742 D.n3741 0.001
R27572 D.n3728 D.n3727 0.001
R27573 D.n3714 D.n3713 0.001
R27574 D.n3700 D.n3699 0.001
R27575 D.n3686 D.n3685 0.001
R27576 D.n3672 D.n3671 0.001
R27577 D.n3658 D.n3657 0.001
R27578 D.n3644 D.n3643 0.001
R27579 D.n3630 D.n3629 0.001
R27580 D.n3616 D.n3615 0.001
R27581 D.n3602 D.n3601 0.001
R27582 D.n3588 D.n3587 0.001
R27583 D.n3574 D.n3573 0.001
R27584 D.n3560 D.n3559 0.001
R27585 D.n3546 D.n3545 0.001
R27586 D.n3532 D.n3531 0.001
R27587 D.n3518 D.n3517 0.001
R27588 D.n3504 D.n3503 0.001
R27589 D.n3490 D.n3489 0.001
R27590 D.n3476 D.n3475 0.001
R27591 D.n3462 D.n3461 0.001
R27592 D.n3448 D.n3447 0.001
R27593 D.n3434 D.n3433 0.001
R27594 D.n3420 D.n3419 0.001
R27595 D.n3406 D.n3405 0.001
R27596 D.n3392 D.n3391 0.001
R27597 D.n4314 D.n4313 0.001
R27598 D.n4300 D.n4299 0.001
R27599 D.n4286 D.n4285 0.001
R27600 D.n4272 D.n4271 0.001
R27601 D.n4258 D.n4257 0.001
R27602 D.n4244 D.n4243 0.001
R27603 D.n4230 D.n4229 0.001
R27604 D.n4216 D.n4215 0.001
R27605 D.n4202 D.n4201 0.001
R27606 D.n4188 D.n4187 0.001
R27607 D.n4174 D.n4173 0.001
R27608 D.n4160 D.n4159 0.001
R27609 D.n4146 D.n4145 0.001
R27610 D.n4132 D.n4131 0.001
R27611 D.n4118 D.n4117 0.001
R27612 D.n4104 D.n4103 0.001
R27613 D.n4090 D.n4089 0.001
R27614 D.n4076 D.n4075 0.001
R27615 D.n4062 D.n4061 0.001
R27616 D.n4048 D.n4047 0.001
R27617 D.n4034 D.n4033 0.001
R27618 D.n4020 D.n4019 0.001
R27619 D.n4006 D.n4005 0.001
R27620 D.n3992 D.n3991 0.001
R27621 D.n3978 D.n3977 0.001
R27622 D.n3964 D.n3963 0.001
R27623 D.n3950 D.n3949 0.001
R27624 D.n3936 D.n3935 0.001
R27625 D.n3922 D.n3921 0.001
R27626 D.n3908 D.n3907 0.001
R27627 D.n3894 D.n3893 0.001
R27628 D.n3880 D.n3879 0.001
R27629 D.n4746 D.n4745 0.001
R27630 D.n4732 D.n4731 0.001
R27631 D.n4718 D.n4717 0.001
R27632 D.n4704 D.n4703 0.001
R27633 D.n4690 D.n4689 0.001
R27634 D.n4676 D.n4675 0.001
R27635 D.n4662 D.n4661 0.001
R27636 D.n4648 D.n4647 0.001
R27637 D.n4634 D.n4633 0.001
R27638 D.n4620 D.n4619 0.001
R27639 D.n4606 D.n4605 0.001
R27640 D.n4592 D.n4591 0.001
R27641 D.n4578 D.n4577 0.001
R27642 D.n4564 D.n4563 0.001
R27643 D.n4550 D.n4549 0.001
R27644 D.n4536 D.n4535 0.001
R27645 D.n4522 D.n4521 0.001
R27646 D.n4508 D.n4507 0.001
R27647 D.n4494 D.n4493 0.001
R27648 D.n4480 D.n4479 0.001
R27649 D.n4466 D.n4465 0.001
R27650 D.n4452 D.n4451 0.001
R27651 D.n4438 D.n4437 0.001
R27652 D.n4424 D.n4423 0.001
R27653 D.n4410 D.n4409 0.001
R27654 D.n4396 D.n4395 0.001
R27655 D.n4382 D.n4381 0.001
R27656 D.n4368 D.n4367 0.001
R27657 D.n4354 D.n4353 0.001
R27658 D.n4340 D.n4339 0.001
R27659 D.n5150 D.n5149 0.001
R27660 D.n5136 D.n5135 0.001
R27661 D.n5122 D.n5121 0.001
R27662 D.n5108 D.n5107 0.001
R27663 D.n5094 D.n5093 0.001
R27664 D.n5080 D.n5079 0.001
R27665 D.n5066 D.n5065 0.001
R27666 D.n5052 D.n5051 0.001
R27667 D.n5038 D.n5037 0.001
R27668 D.n5024 D.n5023 0.001
R27669 D.n5010 D.n5009 0.001
R27670 D.n4996 D.n4995 0.001
R27671 D.n4982 D.n4981 0.001
R27672 D.n4968 D.n4967 0.001
R27673 D.n4954 D.n4953 0.001
R27674 D.n4940 D.n4939 0.001
R27675 D.n4926 D.n4925 0.001
R27676 D.n4912 D.n4911 0.001
R27677 D.n4898 D.n4897 0.001
R27678 D.n4884 D.n4883 0.001
R27679 D.n4870 D.n4869 0.001
R27680 D.n4856 D.n4855 0.001
R27681 D.n4842 D.n4841 0.001
R27682 D.n4828 D.n4827 0.001
R27683 D.n4814 D.n4813 0.001
R27684 D.n4800 D.n4799 0.001
R27685 D.n4786 D.n4785 0.001
R27686 D.n4772 D.n4771 0.001
R27687 D.n5526 D.n5525 0.001
R27688 D.n5512 D.n5511 0.001
R27689 D.n5498 D.n5497 0.001
R27690 D.n5484 D.n5483 0.001
R27691 D.n5470 D.n5469 0.001
R27692 D.n5456 D.n5455 0.001
R27693 D.n5442 D.n5441 0.001
R27694 D.n5428 D.n5427 0.001
R27695 D.n5414 D.n5413 0.001
R27696 D.n5400 D.n5399 0.001
R27697 D.n5386 D.n5385 0.001
R27698 D.n5372 D.n5371 0.001
R27699 D.n5358 D.n5357 0.001
R27700 D.n5344 D.n5343 0.001
R27701 D.n5330 D.n5329 0.001
R27702 D.n5316 D.n5315 0.001
R27703 D.n5302 D.n5301 0.001
R27704 D.n5288 D.n5287 0.001
R27705 D.n5274 D.n5273 0.001
R27706 D.n5260 D.n5259 0.001
R27707 D.n5246 D.n5245 0.001
R27708 D.n5232 D.n5231 0.001
R27709 D.n5218 D.n5217 0.001
R27710 D.n5204 D.n5203 0.001
R27711 D.n5190 D.n5189 0.001
R27712 D.n5176 D.n5175 0.001
R27713 D.n5874 D.n5873 0.001
R27714 D.n5860 D.n5859 0.001
R27715 D.n5846 D.n5845 0.001
R27716 D.n5832 D.n5831 0.001
R27717 D.n5818 D.n5817 0.001
R27718 D.n5804 D.n5803 0.001
R27719 D.n5790 D.n5789 0.001
R27720 D.n5776 D.n5775 0.001
R27721 D.n5762 D.n5761 0.001
R27722 D.n5748 D.n5747 0.001
R27723 D.n5734 D.n5733 0.001
R27724 D.n5720 D.n5719 0.001
R27725 D.n5706 D.n5705 0.001
R27726 D.n5692 D.n5691 0.001
R27727 D.n5678 D.n5677 0.001
R27728 D.n5664 D.n5663 0.001
R27729 D.n5650 D.n5649 0.001
R27730 D.n5636 D.n5635 0.001
R27731 D.n5622 D.n5621 0.001
R27732 D.n5608 D.n5607 0.001
R27733 D.n5594 D.n5593 0.001
R27734 D.n5580 D.n5579 0.001
R27735 D.n5566 D.n5565 0.001
R27736 D.n5552 D.n5551 0.001
R27737 D.n6194 D.n6193 0.001
R27738 D.n6180 D.n6179 0.001
R27739 D.n6166 D.n6165 0.001
R27740 D.n6152 D.n6151 0.001
R27741 D.n6138 D.n6137 0.001
R27742 D.n6124 D.n6123 0.001
R27743 D.n6110 D.n6109 0.001
R27744 D.n6096 D.n6095 0.001
R27745 D.n6082 D.n6081 0.001
R27746 D.n6068 D.n6067 0.001
R27747 D.n6054 D.n6053 0.001
R27748 D.n6040 D.n6039 0.001
R27749 D.n6026 D.n6025 0.001
R27750 D.n6012 D.n6011 0.001
R27751 D.n5998 D.n5997 0.001
R27752 D.n5984 D.n5983 0.001
R27753 D.n5970 D.n5969 0.001
R27754 D.n5956 D.n5955 0.001
R27755 D.n5942 D.n5941 0.001
R27756 D.n5928 D.n5927 0.001
R27757 D.n5914 D.n5913 0.001
R27758 D.n5900 D.n5899 0.001
R27759 D.n6486 D.n6485 0.001
R27760 D.n6472 D.n6471 0.001
R27761 D.n6458 D.n6457 0.001
R27762 D.n6444 D.n6443 0.001
R27763 D.n6430 D.n6429 0.001
R27764 D.n6416 D.n6415 0.001
R27765 D.n6402 D.n6401 0.001
R27766 D.n6388 D.n6387 0.001
R27767 D.n6374 D.n6373 0.001
R27768 D.n6360 D.n6359 0.001
R27769 D.n6346 D.n6345 0.001
R27770 D.n6332 D.n6331 0.001
R27771 D.n6318 D.n6317 0.001
R27772 D.n6304 D.n6303 0.001
R27773 D.n6290 D.n6289 0.001
R27774 D.n6276 D.n6275 0.001
R27775 D.n6262 D.n6261 0.001
R27776 D.n6248 D.n6247 0.001
R27777 D.n6234 D.n6233 0.001
R27778 D.n6220 D.n6219 0.001
R27779 D.n6750 D.n6749 0.001
R27780 D.n6736 D.n6735 0.001
R27781 D.n6722 D.n6721 0.001
R27782 D.n6708 D.n6707 0.001
R27783 D.n6694 D.n6693 0.001
R27784 D.n6680 D.n6679 0.001
R27785 D.n6666 D.n6665 0.001
R27786 D.n6652 D.n6651 0.001
R27787 D.n6638 D.n6637 0.001
R27788 D.n6624 D.n6623 0.001
R27789 D.n6610 D.n6609 0.001
R27790 D.n6596 D.n6595 0.001
R27791 D.n6582 D.n6581 0.001
R27792 D.n6568 D.n6567 0.001
R27793 D.n6554 D.n6553 0.001
R27794 D.n6540 D.n6539 0.001
R27795 D.n6526 D.n6525 0.001
R27796 D.n6512 D.n6511 0.001
R27797 D.n6986 D.n6985 0.001
R27798 D.n6972 D.n6971 0.001
R27799 D.n6958 D.n6957 0.001
R27800 D.n6944 D.n6943 0.001
R27801 D.n6930 D.n6929 0.001
R27802 D.n6916 D.n6915 0.001
R27803 D.n6902 D.n6901 0.001
R27804 D.n6888 D.n6887 0.001
R27805 D.n6874 D.n6873 0.001
R27806 D.n6860 D.n6859 0.001
R27807 D.n6846 D.n6845 0.001
R27808 D.n6832 D.n6831 0.001
R27809 D.n6818 D.n6817 0.001
R27810 D.n6804 D.n6803 0.001
R27811 D.n6790 D.n6789 0.001
R27812 D.n6776 D.n6775 0.001
R27813 D.n7194 D.n7193 0.001
R27814 D.n7180 D.n7179 0.001
R27815 D.n7166 D.n7165 0.001
R27816 D.n7152 D.n7151 0.001
R27817 D.n7138 D.n7137 0.001
R27818 D.n7124 D.n7123 0.001
R27819 D.n7110 D.n7109 0.001
R27820 D.n7096 D.n7095 0.001
R27821 D.n7082 D.n7081 0.001
R27822 D.n7068 D.n7067 0.001
R27823 D.n7054 D.n7053 0.001
R27824 D.n7040 D.n7039 0.001
R27825 D.n7026 D.n7025 0.001
R27826 D.n7012 D.n7011 0.001
R27827 D.n7374 D.n7373 0.001
R27828 D.n7360 D.n7359 0.001
R27829 D.n7346 D.n7345 0.001
R27830 D.n7332 D.n7331 0.001
R27831 D.n7318 D.n7317 0.001
R27832 D.n7304 D.n7303 0.001
R27833 D.n7290 D.n7289 0.001
R27834 D.n7276 D.n7275 0.001
R27835 D.n7262 D.n7261 0.001
R27836 D.n7248 D.n7247 0.001
R27837 D.n7234 D.n7233 0.001
R27838 D.n7220 D.n7219 0.001
R27839 D.n7526 D.n7525 0.001
R27840 D.n7512 D.n7511 0.001
R27841 D.n7498 D.n7497 0.001
R27842 D.n7484 D.n7483 0.001
R27843 D.n7470 D.n7469 0.001
R27844 D.n7456 D.n7455 0.001
R27845 D.n7442 D.n7441 0.001
R27846 D.n7428 D.n7427 0.001
R27847 D.n7414 D.n7413 0.001
R27848 D.n7400 D.n7399 0.001
R27849 D.n7650 D.n7649 0.001
R27850 D.n7636 D.n7635 0.001
R27851 D.n7622 D.n7621 0.001
R27852 D.n7608 D.n7607 0.001
R27853 D.n7594 D.n7593 0.001
R27854 D.n7580 D.n7579 0.001
R27855 D.n7566 D.n7565 0.001
R27856 D.n7552 D.n7551 0.001
R27857 D.n7746 D.n7745 0.001
R27858 D.n7732 D.n7731 0.001
R27859 D.n7718 D.n7717 0.001
R27860 D.n7704 D.n7703 0.001
R27861 D.n7690 D.n7689 0.001
R27862 D.n7676 D.n7675 0.001
R27863 D.n7815 D.n7814 0.001
R27864 D.n7799 D.n7798 0.001
R27865 D.n7785 D.n7784 0.001
R27866 D.n7771 D.n7770 0.001
R27867 D.n508 D.n503 0.001
R27868 D.n7856 D.n7854 0.001
R27869 D.n7849 D.n7818 0.001
R27870 D.n7842 D.n7840 0.001
R27871 D.n7832 D.n7830 0.001
R27872 D.n453 D.n451 0.001
R27873 D.n444 D.n442 0.001
R27874 D.n47 D.n33 0.001
R27875 D.n7933 D.n7931 0.001
R27876 D.n7962 D.n7960 0.001
R27877 D.n7952 D.n7945 0.001
R27878 D.n14067 D.n14065 0.001
R27879 D.n14049 D.n14047 0.001
R27880 D.n14031 D.n14029 0.001
R27881 D.n14013 D.n14011 0.001
R27882 D.n13995 D.n13993 0.001
R27883 D.n13977 D.n13975 0.001
R27884 D.n13959 D.n13957 0.001
R27885 D.n13941 D.n13939 0.001
R27886 D.n13923 D.n13921 0.001
R27887 D.n13905 D.n13903 0.001
R27888 D.n13887 D.n13885 0.001
R27889 D.n13869 D.n13867 0.001
R27890 D.n13851 D.n13849 0.001
R27891 D.n13833 D.n13831 0.001
R27892 D.n13815 D.n13813 0.001
R27893 D.n13797 D.n13795 0.001
R27894 D.n13779 D.n13777 0.001
R27895 D.n13761 D.n13759 0.001
R27896 D.n13743 D.n13741 0.001
R27897 D.n13725 D.n13723 0.001
R27898 D.n13707 D.n13705 0.001
R27899 D.n13689 D.n13686 0.001
R27900 D.n13698 D.n13696 0.001
R27901 D.n13716 D.n13714 0.001
R27902 D.n13734 D.n13732 0.001
R27903 D.n13752 D.n13750 0.001
R27904 D.n13770 D.n13768 0.001
R27905 D.n13788 D.n13786 0.001
R27906 D.n13806 D.n13804 0.001
R27907 D.n13824 D.n13822 0.001
R27908 D.n13842 D.n13840 0.001
R27909 D.n13860 D.n13858 0.001
R27910 D.n13878 D.n13876 0.001
R27911 D.n13896 D.n13894 0.001
R27912 D.n13914 D.n13912 0.001
R27913 D.n13932 D.n13930 0.001
R27914 D.n13950 D.n13948 0.001
R27915 D.n13968 D.n13966 0.001
R27916 D.n13986 D.n13984 0.001
R27917 D.n14004 D.n14002 0.001
R27918 D.n14022 D.n14020 0.001
R27919 D.n14040 D.n14038 0.001
R27920 D.n14058 D.n14056 0.001
R27921 D.n14081 D.n14078 0.001
R27922 D.n14096 D.n14091 0.001
R27923 D.n13212 D.n13211 0.001
R27924 D.n13232 D.n13231 0.001
R27925 D.n13252 D.n13251 0.001
R27926 D.n13272 D.n13271 0.001
R27927 D.n13292 D.n13291 0.001
R27928 D.n13312 D.n13311 0.001
R27929 D.n13332 D.n13331 0.001
R27930 D.n13352 D.n13351 0.001
R27931 D.n13372 D.n13371 0.001
R27932 D.n13392 D.n13391 0.001
R27933 D.n13412 D.n13411 0.001
R27934 D.n13432 D.n13431 0.001
R27935 D.n13452 D.n13451 0.001
R27936 D.n13472 D.n13471 0.001
R27937 D.n13492 D.n13491 0.001
R27938 D.n13512 D.n13511 0.001
R27939 D.n13532 D.n13531 0.001
R27940 D.n13552 D.n13551 0.001
R27941 D.n13572 D.n13571 0.001
R27942 D.n13592 D.n13591 0.001
R27943 D.n13612 D.n13611 0.001
R27944 D.n13602 D.n13600 0.001
R27945 D.n13582 D.n13580 0.001
R27946 D.n13562 D.n13560 0.001
R27947 D.n13542 D.n13540 0.001
R27948 D.n13522 D.n13520 0.001
R27949 D.n13502 D.n13500 0.001
R27950 D.n13482 D.n13480 0.001
R27951 D.n13462 D.n13460 0.001
R27952 D.n13442 D.n13440 0.001
R27953 D.n13422 D.n13420 0.001
R27954 D.n13402 D.n13400 0.001
R27955 D.n13382 D.n13380 0.001
R27956 D.n13362 D.n13360 0.001
R27957 D.n13342 D.n13340 0.001
R27958 D.n13322 D.n13320 0.001
R27959 D.n13302 D.n13300 0.001
R27960 D.n13282 D.n13280 0.001
R27961 D.n13262 D.n13260 0.001
R27962 D.n13242 D.n13240 0.001
R27963 D.n13222 D.n13220 0.001
R27964 D.n13202 D.n13195 0.001
R27965 D.n13183 D.n13178 0.001
R27966 D.n13104 D.n13102 0.001
R27967 D.n13086 D.n13084 0.001
R27968 D.n13068 D.n13066 0.001
R27969 D.n13050 D.n13048 0.001
R27970 D.n13032 D.n13030 0.001
R27971 D.n13014 D.n13012 0.001
R27972 D.n12996 D.n12994 0.001
R27973 D.n12978 D.n12976 0.001
R27974 D.n12960 D.n12958 0.001
R27975 D.n12942 D.n12940 0.001
R27976 D.n12924 D.n12922 0.001
R27977 D.n12906 D.n12904 0.001
R27978 D.n12888 D.n12886 0.001
R27979 D.n12870 D.n12868 0.001
R27980 D.n12852 D.n12850 0.001
R27981 D.n12834 D.n12832 0.001
R27982 D.n12816 D.n12814 0.001
R27983 D.n12798 D.n12796 0.001
R27984 D.n12780 D.n12778 0.001
R27985 D.n12762 D.n12759 0.001
R27986 D.n12771 D.n12769 0.001
R27987 D.n12789 D.n12787 0.001
R27988 D.n12807 D.n12805 0.001
R27989 D.n12825 D.n12823 0.001
R27990 D.n12843 D.n12841 0.001
R27991 D.n12861 D.n12859 0.001
R27992 D.n12879 D.n12877 0.001
R27993 D.n12897 D.n12895 0.001
R27994 D.n12915 D.n12913 0.001
R27995 D.n12933 D.n12931 0.001
R27996 D.n12951 D.n12949 0.001
R27997 D.n12969 D.n12967 0.001
R27998 D.n12987 D.n12985 0.001
R27999 D.n13005 D.n13003 0.001
R28000 D.n13023 D.n13021 0.001
R28001 D.n13041 D.n13039 0.001
R28002 D.n13059 D.n13057 0.001
R28003 D.n13077 D.n13075 0.001
R28004 D.n13095 D.n13093 0.001
R28005 D.n13117 D.n13114 0.001
R28006 D.n13127 D.n13121 0.001
R28007 D.n12329 D.n12328 0.001
R28008 D.n12349 D.n12348 0.001
R28009 D.n12369 D.n12368 0.001
R28010 D.n12389 D.n12388 0.001
R28011 D.n12409 D.n12408 0.001
R28012 D.n12429 D.n12428 0.001
R28013 D.n12449 D.n12448 0.001
R28014 D.n12469 D.n12468 0.001
R28015 D.n12489 D.n12488 0.001
R28016 D.n12509 D.n12508 0.001
R28017 D.n12529 D.n12528 0.001
R28018 D.n12549 D.n12548 0.001
R28019 D.n12569 D.n12568 0.001
R28020 D.n12589 D.n12588 0.001
R28021 D.n12609 D.n12608 0.001
R28022 D.n12629 D.n12628 0.001
R28023 D.n12649 D.n12648 0.001
R28024 D.n12669 D.n12668 0.001
R28025 D.n12689 D.n12688 0.001
R28026 D.n12679 D.n12677 0.001
R28027 D.n12659 D.n12657 0.001
R28028 D.n12639 D.n12637 0.001
R28029 D.n12619 D.n12617 0.001
R28030 D.n12599 D.n12597 0.001
R28031 D.n12579 D.n12577 0.001
R28032 D.n12559 D.n12557 0.001
R28033 D.n12539 D.n12537 0.001
R28034 D.n12519 D.n12517 0.001
R28035 D.n12499 D.n12497 0.001
R28036 D.n12479 D.n12477 0.001
R28037 D.n12459 D.n12457 0.001
R28038 D.n12439 D.n12437 0.001
R28039 D.n12419 D.n12417 0.001
R28040 D.n12399 D.n12397 0.001
R28041 D.n12379 D.n12377 0.001
R28042 D.n12359 D.n12357 0.001
R28043 D.n12339 D.n12337 0.001
R28044 D.n12319 D.n12312 0.001
R28045 D.n12300 D.n12295 0.001
R28046 D.n12219 D.n12217 0.001
R28047 D.n12201 D.n12199 0.001
R28048 D.n12183 D.n12181 0.001
R28049 D.n12165 D.n12163 0.001
R28050 D.n12147 D.n12145 0.001
R28051 D.n12129 D.n12127 0.001
R28052 D.n12111 D.n12109 0.001
R28053 D.n12093 D.n12091 0.001
R28054 D.n12075 D.n12073 0.001
R28055 D.n12057 D.n12055 0.001
R28056 D.n12039 D.n12037 0.001
R28057 D.n12021 D.n12019 0.001
R28058 D.n12003 D.n12001 0.001
R28059 D.n11985 D.n11983 0.001
R28060 D.n11967 D.n11965 0.001
R28061 D.n11949 D.n11947 0.001
R28062 D.n11931 D.n11929 0.001
R28063 D.n11913 D.n11910 0.001
R28064 D.n11922 D.n11920 0.001
R28065 D.n11940 D.n11938 0.001
R28066 D.n11958 D.n11956 0.001
R28067 D.n11976 D.n11974 0.001
R28068 D.n11994 D.n11992 0.001
R28069 D.n12012 D.n12010 0.001
R28070 D.n12030 D.n12028 0.001
R28071 D.n12048 D.n12046 0.001
R28072 D.n12066 D.n12064 0.001
R28073 D.n12084 D.n12082 0.001
R28074 D.n12102 D.n12100 0.001
R28075 D.n12120 D.n12118 0.001
R28076 D.n12138 D.n12136 0.001
R28077 D.n12156 D.n12154 0.001
R28078 D.n12174 D.n12172 0.001
R28079 D.n12192 D.n12190 0.001
R28080 D.n12210 D.n12208 0.001
R28081 D.n12232 D.n12230 0.001
R28082 D.n12248 D.n12243 0.001
R28083 D.n11520 D.n11519 0.001
R28084 D.n11540 D.n11539 0.001
R28085 D.n11560 D.n11559 0.001
R28086 D.n11580 D.n11579 0.001
R28087 D.n11600 D.n11599 0.001
R28088 D.n11620 D.n11619 0.001
R28089 D.n11640 D.n11639 0.001
R28090 D.n11660 D.n11659 0.001
R28091 D.n11680 D.n11679 0.001
R28092 D.n11700 D.n11699 0.001
R28093 D.n11720 D.n11719 0.001
R28094 D.n11740 D.n11739 0.001
R28095 D.n11760 D.n11759 0.001
R28096 D.n11780 D.n11779 0.001
R28097 D.n11800 D.n11799 0.001
R28098 D.n11820 D.n11819 0.001
R28099 D.n11840 D.n11839 0.001
R28100 D.n11830 D.n11828 0.001
R28101 D.n11810 D.n11808 0.001
R28102 D.n11790 D.n11788 0.001
R28103 D.n11770 D.n11768 0.001
R28104 D.n11750 D.n11748 0.001
R28105 D.n11730 D.n11728 0.001
R28106 D.n11710 D.n11708 0.001
R28107 D.n11690 D.n11688 0.001
R28108 D.n11670 D.n11668 0.001
R28109 D.n11650 D.n11648 0.001
R28110 D.n11630 D.n11628 0.001
R28111 D.n11610 D.n11608 0.001
R28112 D.n11590 D.n11588 0.001
R28113 D.n11570 D.n11568 0.001
R28114 D.n11550 D.n11548 0.001
R28115 D.n11530 D.n11528 0.001
R28116 D.n11510 D.n11505 0.001
R28117 D.n11495 D.n11491 0.001
R28118 D.n11420 D.n11418 0.001
R28119 D.n11402 D.n11400 0.001
R28120 D.n11384 D.n11382 0.001
R28121 D.n11366 D.n11364 0.001
R28122 D.n11348 D.n11346 0.001
R28123 D.n11330 D.n11328 0.001
R28124 D.n11312 D.n11310 0.001
R28125 D.n11294 D.n11292 0.001
R28126 D.n11276 D.n11274 0.001
R28127 D.n11258 D.n11256 0.001
R28128 D.n11240 D.n11238 0.001
R28129 D.n11222 D.n11220 0.001
R28130 D.n11204 D.n11202 0.001
R28131 D.n11186 D.n11184 0.001
R28132 D.n11168 D.n11166 0.001
R28133 D.n11150 D.n11147 0.001
R28134 D.n11159 D.n11157 0.001
R28135 D.n11177 D.n11175 0.001
R28136 D.n11195 D.n11193 0.001
R28137 D.n11213 D.n11211 0.001
R28138 D.n11231 D.n11229 0.001
R28139 D.n11249 D.n11247 0.001
R28140 D.n11267 D.n11265 0.001
R28141 D.n11285 D.n11283 0.001
R28142 D.n11303 D.n11301 0.001
R28143 D.n11321 D.n11319 0.001
R28144 D.n11339 D.n11337 0.001
R28145 D.n11357 D.n11355 0.001
R28146 D.n11375 D.n11373 0.001
R28147 D.n11393 D.n11391 0.001
R28148 D.n11411 D.n11409 0.001
R28149 D.n11433 D.n11431 0.001
R28150 D.n11449 D.n11444 0.001
R28151 D.n10797 D.n10796 0.001
R28152 D.n10817 D.n10816 0.001
R28153 D.n10837 D.n10836 0.001
R28154 D.n10857 D.n10856 0.001
R28155 D.n10877 D.n10876 0.001
R28156 D.n10897 D.n10896 0.001
R28157 D.n10917 D.n10916 0.001
R28158 D.n10937 D.n10936 0.001
R28159 D.n10957 D.n10956 0.001
R28160 D.n10977 D.n10976 0.001
R28161 D.n10997 D.n10996 0.001
R28162 D.n11017 D.n11016 0.001
R28163 D.n11037 D.n11036 0.001
R28164 D.n11057 D.n11056 0.001
R28165 D.n11077 D.n11076 0.001
R28166 D.n11067 D.n11065 0.001
R28167 D.n11047 D.n11045 0.001
R28168 D.n11027 D.n11025 0.001
R28169 D.n11007 D.n11005 0.001
R28170 D.n10987 D.n10985 0.001
R28171 D.n10967 D.n10965 0.001
R28172 D.n10947 D.n10945 0.001
R28173 D.n10927 D.n10925 0.001
R28174 D.n10907 D.n10905 0.001
R28175 D.n10887 D.n10885 0.001
R28176 D.n10867 D.n10865 0.001
R28177 D.n10847 D.n10845 0.001
R28178 D.n10827 D.n10825 0.001
R28179 D.n10807 D.n10805 0.001
R28180 D.n10787 D.n10782 0.001
R28181 D.n10772 D.n10768 0.001
R28182 D.n10701 D.n10699 0.001
R28183 D.n10683 D.n10681 0.001
R28184 D.n10665 D.n10663 0.001
R28185 D.n10647 D.n10645 0.001
R28186 D.n10629 D.n10627 0.001
R28187 D.n10611 D.n10609 0.001
R28188 D.n10593 D.n10591 0.001
R28189 D.n10575 D.n10573 0.001
R28190 D.n10557 D.n10555 0.001
R28191 D.n10539 D.n10537 0.001
R28192 D.n10521 D.n10519 0.001
R28193 D.n10503 D.n10501 0.001
R28194 D.n10485 D.n10483 0.001
R28195 D.n10467 D.n10464 0.001
R28196 D.n10476 D.n10474 0.001
R28197 D.n10494 D.n10492 0.001
R28198 D.n10512 D.n10510 0.001
R28199 D.n10530 D.n10528 0.001
R28200 D.n10548 D.n10546 0.001
R28201 D.n10566 D.n10564 0.001
R28202 D.n10584 D.n10582 0.001
R28203 D.n10602 D.n10600 0.001
R28204 D.n10620 D.n10618 0.001
R28205 D.n10638 D.n10636 0.001
R28206 D.n10656 D.n10654 0.001
R28207 D.n10674 D.n10672 0.001
R28208 D.n10692 D.n10690 0.001
R28209 D.n10714 D.n10712 0.001
R28210 D.n10730 D.n10725 0.001
R28211 D.n10154 D.n10153 0.001
R28212 D.n10174 D.n10173 0.001
R28213 D.n10194 D.n10193 0.001
R28214 D.n10214 D.n10213 0.001
R28215 D.n10234 D.n10233 0.001
R28216 D.n10254 D.n10253 0.001
R28217 D.n10274 D.n10273 0.001
R28218 D.n10294 D.n10293 0.001
R28219 D.n10314 D.n10313 0.001
R28220 D.n10334 D.n10333 0.001
R28221 D.n10354 D.n10353 0.001
R28222 D.n10374 D.n10373 0.001
R28223 D.n10394 D.n10393 0.001
R28224 D.n10384 D.n10382 0.001
R28225 D.n10364 D.n10362 0.001
R28226 D.n10344 D.n10342 0.001
R28227 D.n10324 D.n10322 0.001
R28228 D.n10304 D.n10302 0.001
R28229 D.n10284 D.n10282 0.001
R28230 D.n10264 D.n10262 0.001
R28231 D.n10244 D.n10242 0.001
R28232 D.n10224 D.n10222 0.001
R28233 D.n10204 D.n10202 0.001
R28234 D.n10184 D.n10182 0.001
R28235 D.n10164 D.n10162 0.001
R28236 D.n10144 D.n10137 0.001
R28237 D.n10125 D.n10120 0.001
R28238 D.n10062 D.n10060 0.001
R28239 D.n10044 D.n10042 0.001
R28240 D.n10026 D.n10024 0.001
R28241 D.n10008 D.n10006 0.001
R28242 D.n9990 D.n9988 0.001
R28243 D.n9972 D.n9970 0.001
R28244 D.n9954 D.n9952 0.001
R28245 D.n9936 D.n9934 0.001
R28246 D.n9918 D.n9916 0.001
R28247 D.n9900 D.n9898 0.001
R28248 D.n9882 D.n9880 0.001
R28249 D.n9864 D.n9861 0.001
R28250 D.n9873 D.n9871 0.001
R28251 D.n9891 D.n9889 0.001
R28252 D.n9909 D.n9907 0.001
R28253 D.n9927 D.n9925 0.001
R28254 D.n9945 D.n9943 0.001
R28255 D.n9963 D.n9961 0.001
R28256 D.n9981 D.n9979 0.001
R28257 D.n9999 D.n9997 0.001
R28258 D.n10017 D.n10015 0.001
R28259 D.n10035 D.n10033 0.001
R28260 D.n10053 D.n10051 0.001
R28261 D.n10075 D.n10072 0.001
R28262 D.n10085 D.n10079 0.001
R28263 D.n9591 D.n9590 0.001
R28264 D.n9611 D.n9610 0.001
R28265 D.n9631 D.n9630 0.001
R28266 D.n9651 D.n9650 0.001
R28267 D.n9671 D.n9670 0.001
R28268 D.n9691 D.n9690 0.001
R28269 D.n9711 D.n9710 0.001
R28270 D.n9731 D.n9730 0.001
R28271 D.n9751 D.n9750 0.001
R28272 D.n9771 D.n9770 0.001
R28273 D.n9791 D.n9790 0.001
R28274 D.n9781 D.n9779 0.001
R28275 D.n9761 D.n9759 0.001
R28276 D.n9741 D.n9739 0.001
R28277 D.n9721 D.n9719 0.001
R28278 D.n9701 D.n9699 0.001
R28279 D.n9681 D.n9679 0.001
R28280 D.n9661 D.n9659 0.001
R28281 D.n9641 D.n9639 0.001
R28282 D.n9621 D.n9619 0.001
R28283 D.n9601 D.n9599 0.001
R28284 D.n9581 D.n9574 0.001
R28285 D.n9562 D.n9557 0.001
R28286 D.n9497 D.n9495 0.001
R28287 D.n9479 D.n9477 0.001
R28288 D.n9461 D.n9459 0.001
R28289 D.n9443 D.n9441 0.001
R28290 D.n9425 D.n9423 0.001
R28291 D.n9407 D.n9405 0.001
R28292 D.n9389 D.n9387 0.001
R28293 D.n9371 D.n9369 0.001
R28294 D.n9353 D.n9351 0.001
R28295 D.n9335 D.n9332 0.001
R28296 D.n9344 D.n9342 0.001
R28297 D.n9362 D.n9360 0.001
R28298 D.n9380 D.n9378 0.001
R28299 D.n9398 D.n9396 0.001
R28300 D.n9416 D.n9414 0.001
R28301 D.n9434 D.n9432 0.001
R28302 D.n9452 D.n9450 0.001
R28303 D.n9470 D.n9468 0.001
R28304 D.n9488 D.n9486 0.001
R28305 D.n9510 D.n9508 0.001
R28306 D.n9526 D.n9521 0.001
R28307 D.n9102 D.n9101 0.001
R28308 D.n9122 D.n9121 0.001
R28309 D.n9142 D.n9141 0.001
R28310 D.n9162 D.n9161 0.001
R28311 D.n9182 D.n9181 0.001
R28312 D.n9202 D.n9201 0.001
R28313 D.n9222 D.n9221 0.001
R28314 D.n9242 D.n9241 0.001
R28315 D.n9262 D.n9261 0.001
R28316 D.n9252 D.n9250 0.001
R28317 D.n9232 D.n9230 0.001
R28318 D.n9212 D.n9210 0.001
R28319 D.n9192 D.n9190 0.001
R28320 D.n9172 D.n9170 0.001
R28321 D.n9152 D.n9150 0.001
R28322 D.n9132 D.n9130 0.001
R28323 D.n9112 D.n9110 0.001
R28324 D.n9092 D.n9087 0.001
R28325 D.n9077 D.n9073 0.001
R28326 D.n9018 D.n9016 0.001
R28327 D.n9000 D.n8998 0.001
R28328 D.n8982 D.n8980 0.001
R28329 D.n8964 D.n8962 0.001
R28330 D.n8946 D.n8944 0.001
R28331 D.n8928 D.n8926 0.001
R28332 D.n8910 D.n8908 0.001
R28333 D.n8892 D.n8889 0.001
R28334 D.n8901 D.n8899 0.001
R28335 D.n8919 D.n8917 0.001
R28336 D.n8937 D.n8935 0.001
R28337 D.n8955 D.n8953 0.001
R28338 D.n8973 D.n8971 0.001
R28339 D.n8991 D.n8989 0.001
R28340 D.n9009 D.n9007 0.001
R28341 D.n9031 D.n9029 0.001
R28342 D.n9047 D.n9042 0.001
R28343 D.n8699 D.n8698 0.001
R28344 D.n8719 D.n8718 0.001
R28345 D.n8739 D.n8738 0.001
R28346 D.n8759 D.n8758 0.001
R28347 D.n8779 D.n8778 0.001
R28348 D.n8799 D.n8798 0.001
R28349 D.n8819 D.n8818 0.001
R28350 D.n8809 D.n8807 0.001
R28351 D.n8789 D.n8787 0.001
R28352 D.n8769 D.n8767 0.001
R28353 D.n8749 D.n8747 0.001
R28354 D.n8729 D.n8727 0.001
R28355 D.n8709 D.n8707 0.001
R28356 D.n8689 D.n8682 0.001
R28357 D.n8670 D.n8665 0.001
R28358 D.n8619 D.n8617 0.001
R28359 D.n8601 D.n8599 0.001
R28360 D.n8583 D.n8581 0.001
R28361 D.n8565 D.n8563 0.001
R28362 D.n8547 D.n8545 0.001
R28363 D.n8529 D.n8526 0.001
R28364 D.n8538 D.n8536 0.001
R28365 D.n8556 D.n8554 0.001
R28366 D.n8574 D.n8572 0.001
R28367 D.n8592 D.n8590 0.001
R28368 D.n8610 D.n8608 0.001
R28369 D.n8632 D.n8629 0.001
R28370 D.n8642 D.n8636 0.001
R28371 D.n8376 D.n8375 0.001
R28372 D.n8396 D.n8395 0.001
R28373 D.n8416 D.n8415 0.001
R28374 D.n8436 D.n8435 0.001
R28375 D.n8456 D.n8455 0.001
R28376 D.n8446 D.n8444 0.001
R28377 D.n8426 D.n8424 0.001
R28378 D.n8406 D.n8404 0.001
R28379 D.n8386 D.n8384 0.001
R28380 D.n8366 D.n8359 0.001
R28381 D.n8347 D.n8342 0.001
R28382 D.n8294 D.n8292 0.001
R28383 D.n8276 D.n8274 0.001
R28384 D.n8258 D.n8256 0.001
R28385 D.n8240 D.n8237 0.001
R28386 D.n8249 D.n8247 0.001
R28387 D.n8267 D.n8265 0.001
R28388 D.n8285 D.n8283 0.001
R28389 D.n8307 D.n8305 0.001
R28390 D.n8323 D.n8318 0.001
R28391 D.n8127 D.n8126 0.001
R28392 D.n8147 D.n8146 0.001
R28393 D.n8167 D.n8166 0.001
R28394 D.n8157 D.n8155 0.001
R28395 D.n8137 D.n8135 0.001
R28396 D.n8117 D.n8112 0.001
R28397 D.n8102 D.n8098 0.001
R28398 D.n8055 D.n8053 0.001
R28399 D.n8037 D.n8034 0.001
R28400 D.n8046 D.n8044 0.001
R28401 D.n8068 D.n8066 0.001
R28402 D.n8084 D.n8079 0.001
R28403 D.n7917 D.n7910 0.001
R28404 D.n57 D.n55 0.001
R28405 D.n66 D.n64 0.001
R28406 D.n75 D.n73 0.001
R28407 D.n84 D.n82 0.001
R28408 D.n93 D.n91 0.001
R28409 D.n102 D.n100 0.001
R28410 D.n111 D.n109 0.001
R28411 D.n120 D.n118 0.001
R28412 D.n129 D.n127 0.001
R28413 D.n138 D.n136 0.001
R28414 D.n147 D.n145 0.001
R28415 D.n156 D.n154 0.001
R28416 D.n165 D.n163 0.001
R28417 D.n174 D.n172 0.001
R28418 D.n183 D.n181 0.001
R28419 D.n192 D.n190 0.001
R28420 D.n201 D.n199 0.001
R28421 D.n210 D.n208 0.001
R28422 D.n219 D.n217 0.001
R28423 D.n228 D.n226 0.001
R28424 D.n237 D.n235 0.001
R28425 D.n246 D.n244 0.001
R28426 D.n255 D.n253 0.001
R28427 D.n264 D.n262 0.001
R28428 D.n273 D.n271 0.001
R28429 D.n282 D.n280 0.001
R28430 D.n291 D.n289 0.001
R28431 D.n300 D.n298 0.001
R28432 D.n309 D.n307 0.001
R28433 D.n318 D.n316 0.001
R28434 D.n327 D.n325 0.001
R28435 D.n336 D.n334 0.001
R28436 D.n345 D.n343 0.001
R28437 D.n354 D.n352 0.001
R28438 D.n363 D.n361 0.001
R28439 D.n372 D.n370 0.001
R28440 D.n381 D.n379 0.001
R28441 D.n390 D.n388 0.001
R28442 D.n399 D.n397 0.001
R28443 D.n408 D.n406 0.001
R28444 D.n417 D.n415 0.001
R28445 D.n426 D.n424 0.001
R28446 D.n435 D.n433 0.001
R28447 D.n535 D.n527 0.001
R28448 D.n549 D.n543 0.001
R28449 D.n1141 D.n514 0.001
R28450 D.n1137 D.n1131 0.001
R28451 D.n1123 D.n1117 0.001
R28452 D.n1109 D.n1103 0.001
R28453 D.n1095 D.n1089 0.001
R28454 D.n1081 D.n1075 0.001
R28455 D.n1067 D.n1061 0.001
R28456 D.n1053 D.n1047 0.001
R28457 D.n1039 D.n1033 0.001
R28458 D.n1025 D.n1019 0.001
R28459 D.n1011 D.n1005 0.001
R28460 D.n997 D.n991 0.001
R28461 D.n983 D.n977 0.001
R28462 D.n969 D.n963 0.001
R28463 D.n955 D.n949 0.001
R28464 D.n941 D.n935 0.001
R28465 D.n927 D.n921 0.001
R28466 D.n913 D.n907 0.001
R28467 D.n899 D.n893 0.001
R28468 D.n885 D.n879 0.001
R28469 D.n871 D.n865 0.001
R28470 D.n857 D.n851 0.001
R28471 D.n843 D.n837 0.001
R28472 D.n829 D.n823 0.001
R28473 D.n815 D.n809 0.001
R28474 D.n801 D.n795 0.001
R28475 D.n787 D.n781 0.001
R28476 D.n773 D.n767 0.001
R28477 D.n759 D.n753 0.001
R28478 D.n745 D.n739 0.001
R28479 D.n731 D.n725 0.001
R28480 D.n717 D.n711 0.001
R28481 D.n703 D.n697 0.001
R28482 D.n689 D.n683 0.001
R28483 D.n675 D.n669 0.001
R28484 D.n661 D.n655 0.001
R28485 D.n647 D.n641 0.001
R28486 D.n633 D.n627 0.001
R28487 D.n619 D.n613 0.001
R28488 D.n605 D.n599 0.001
R28489 D.n591 D.n585 0.001
R28490 D.n577 D.n571 0.001
R28491 D.n563 D.n557 0.001
R28492 D.n1162 D.n1154 0.001
R28493 D.n1176 D.n1170 0.001
R28494 D.n1740 D.n1144 0.001
R28495 D.n1736 D.n1730 0.001
R28496 D.n1722 D.n1716 0.001
R28497 D.n1708 D.n1702 0.001
R28498 D.n1694 D.n1688 0.001
R28499 D.n1680 D.n1674 0.001
R28500 D.n1666 D.n1660 0.001
R28501 D.n1652 D.n1646 0.001
R28502 D.n1638 D.n1632 0.001
R28503 D.n1624 D.n1618 0.001
R28504 D.n1610 D.n1604 0.001
R28505 D.n1596 D.n1590 0.001
R28506 D.n1582 D.n1576 0.001
R28507 D.n1568 D.n1562 0.001
R28508 D.n1554 D.n1548 0.001
R28509 D.n1540 D.n1534 0.001
R28510 D.n1526 D.n1520 0.001
R28511 D.n1512 D.n1506 0.001
R28512 D.n1498 D.n1492 0.001
R28513 D.n1484 D.n1478 0.001
R28514 D.n1470 D.n1464 0.001
R28515 D.n1456 D.n1450 0.001
R28516 D.n1442 D.n1436 0.001
R28517 D.n1428 D.n1422 0.001
R28518 D.n1414 D.n1408 0.001
R28519 D.n1400 D.n1394 0.001
R28520 D.n1386 D.n1380 0.001
R28521 D.n1372 D.n1366 0.001
R28522 D.n1358 D.n1352 0.001
R28523 D.n1344 D.n1338 0.001
R28524 D.n1330 D.n1324 0.001
R28525 D.n1316 D.n1310 0.001
R28526 D.n1302 D.n1296 0.001
R28527 D.n1288 D.n1282 0.001
R28528 D.n1274 D.n1268 0.001
R28529 D.n1260 D.n1254 0.001
R28530 D.n1246 D.n1240 0.001
R28531 D.n1232 D.n1226 0.001
R28532 D.n1218 D.n1212 0.001
R28533 D.n1204 D.n1198 0.001
R28534 D.n1190 D.n1184 0.001
R28535 D.n1761 D.n1753 0.001
R28536 D.n1775 D.n1769 0.001
R28537 D.n2311 D.n1743 0.001
R28538 D.n2307 D.n2301 0.001
R28539 D.n2293 D.n2287 0.001
R28540 D.n2279 D.n2273 0.001
R28541 D.n2265 D.n2259 0.001
R28542 D.n2251 D.n2245 0.001
R28543 D.n2237 D.n2231 0.001
R28544 D.n2223 D.n2217 0.001
R28545 D.n2209 D.n2203 0.001
R28546 D.n2195 D.n2189 0.001
R28547 D.n2181 D.n2175 0.001
R28548 D.n2167 D.n2161 0.001
R28549 D.n2153 D.n2147 0.001
R28550 D.n2139 D.n2133 0.001
R28551 D.n2125 D.n2119 0.001
R28552 D.n2111 D.n2105 0.001
R28553 D.n2097 D.n2091 0.001
R28554 D.n2083 D.n2077 0.001
R28555 D.n2069 D.n2063 0.001
R28556 D.n2055 D.n2049 0.001
R28557 D.n2041 D.n2035 0.001
R28558 D.n2027 D.n2021 0.001
R28559 D.n2013 D.n2007 0.001
R28560 D.n1999 D.n1993 0.001
R28561 D.n1985 D.n1979 0.001
R28562 D.n1971 D.n1965 0.001
R28563 D.n1957 D.n1951 0.001
R28564 D.n1943 D.n1937 0.001
R28565 D.n1929 D.n1923 0.001
R28566 D.n1915 D.n1909 0.001
R28567 D.n1901 D.n1895 0.001
R28568 D.n1887 D.n1881 0.001
R28569 D.n1873 D.n1867 0.001
R28570 D.n1859 D.n1853 0.001
R28571 D.n1845 D.n1839 0.001
R28572 D.n1831 D.n1825 0.001
R28573 D.n1817 D.n1811 0.001
R28574 D.n1803 D.n1797 0.001
R28575 D.n1789 D.n1783 0.001
R28576 D.n2332 D.n2324 0.001
R28577 D.n2346 D.n2340 0.001
R28578 D.n2854 D.n2314 0.001
R28579 D.n2850 D.n2844 0.001
R28580 D.n2836 D.n2830 0.001
R28581 D.n2822 D.n2816 0.001
R28582 D.n2808 D.n2802 0.001
R28583 D.n2794 D.n2788 0.001
R28584 D.n2780 D.n2774 0.001
R28585 D.n2766 D.n2760 0.001
R28586 D.n2752 D.n2746 0.001
R28587 D.n2738 D.n2732 0.001
R28588 D.n2724 D.n2718 0.001
R28589 D.n2710 D.n2704 0.001
R28590 D.n2696 D.n2690 0.001
R28591 D.n2682 D.n2676 0.001
R28592 D.n2668 D.n2662 0.001
R28593 D.n2654 D.n2648 0.001
R28594 D.n2640 D.n2634 0.001
R28595 D.n2626 D.n2620 0.001
R28596 D.n2612 D.n2606 0.001
R28597 D.n2598 D.n2592 0.001
R28598 D.n2584 D.n2578 0.001
R28599 D.n2570 D.n2564 0.001
R28600 D.n2556 D.n2550 0.001
R28601 D.n2542 D.n2536 0.001
R28602 D.n2528 D.n2522 0.001
R28603 D.n2514 D.n2508 0.001
R28604 D.n2500 D.n2494 0.001
R28605 D.n2486 D.n2480 0.001
R28606 D.n2472 D.n2466 0.001
R28607 D.n2458 D.n2452 0.001
R28608 D.n2444 D.n2438 0.001
R28609 D.n2430 D.n2424 0.001
R28610 D.n2416 D.n2410 0.001
R28611 D.n2402 D.n2396 0.001
R28612 D.n2388 D.n2382 0.001
R28613 D.n2374 D.n2368 0.001
R28614 D.n2360 D.n2354 0.001
R28615 D.n2875 D.n2867 0.001
R28616 D.n2889 D.n2883 0.001
R28617 D.n3369 D.n2857 0.001
R28618 D.n3365 D.n3359 0.001
R28619 D.n3351 D.n3345 0.001
R28620 D.n3337 D.n3331 0.001
R28621 D.n3323 D.n3317 0.001
R28622 D.n3309 D.n3303 0.001
R28623 D.n3295 D.n3289 0.001
R28624 D.n3281 D.n3275 0.001
R28625 D.n3267 D.n3261 0.001
R28626 D.n3253 D.n3247 0.001
R28627 D.n3239 D.n3233 0.001
R28628 D.n3225 D.n3219 0.001
R28629 D.n3211 D.n3205 0.001
R28630 D.n3197 D.n3191 0.001
R28631 D.n3183 D.n3177 0.001
R28632 D.n3169 D.n3163 0.001
R28633 D.n3155 D.n3149 0.001
R28634 D.n3141 D.n3135 0.001
R28635 D.n3127 D.n3121 0.001
R28636 D.n3113 D.n3107 0.001
R28637 D.n3099 D.n3093 0.001
R28638 D.n3085 D.n3079 0.001
R28639 D.n3071 D.n3065 0.001
R28640 D.n3057 D.n3051 0.001
R28641 D.n3043 D.n3037 0.001
R28642 D.n3029 D.n3023 0.001
R28643 D.n3015 D.n3009 0.001
R28644 D.n3001 D.n2995 0.001
R28645 D.n2987 D.n2981 0.001
R28646 D.n2973 D.n2967 0.001
R28647 D.n2959 D.n2953 0.001
R28648 D.n2945 D.n2939 0.001
R28649 D.n2931 D.n2925 0.001
R28650 D.n2917 D.n2911 0.001
R28651 D.n2903 D.n2897 0.001
R28652 D.n3391 D.n3383 0.001
R28653 D.n3405 D.n3399 0.001
R28654 D.n3857 D.n3373 0.001
R28655 D.n3853 D.n3847 0.001
R28656 D.n3839 D.n3833 0.001
R28657 D.n3825 D.n3819 0.001
R28658 D.n3811 D.n3805 0.001
R28659 D.n3797 D.n3791 0.001
R28660 D.n3783 D.n3777 0.001
R28661 D.n3769 D.n3763 0.001
R28662 D.n3755 D.n3749 0.001
R28663 D.n3741 D.n3735 0.001
R28664 D.n3727 D.n3721 0.001
R28665 D.n3713 D.n3707 0.001
R28666 D.n3699 D.n3693 0.001
R28667 D.n3685 D.n3679 0.001
R28668 D.n3671 D.n3665 0.001
R28669 D.n3657 D.n3651 0.001
R28670 D.n3643 D.n3637 0.001
R28671 D.n3629 D.n3623 0.001
R28672 D.n3615 D.n3609 0.001
R28673 D.n3601 D.n3595 0.001
R28674 D.n3587 D.n3581 0.001
R28675 D.n3573 D.n3567 0.001
R28676 D.n3559 D.n3553 0.001
R28677 D.n3545 D.n3539 0.001
R28678 D.n3531 D.n3525 0.001
R28679 D.n3517 D.n3511 0.001
R28680 D.n3503 D.n3497 0.001
R28681 D.n3489 D.n3483 0.001
R28682 D.n3475 D.n3469 0.001
R28683 D.n3461 D.n3455 0.001
R28684 D.n3447 D.n3441 0.001
R28685 D.n3433 D.n3427 0.001
R28686 D.n3419 D.n3413 0.001
R28687 D.n3879 D.n3871 0.001
R28688 D.n3893 D.n3887 0.001
R28689 D.n4317 D.n3861 0.001
R28690 D.n4313 D.n4307 0.001
R28691 D.n4299 D.n4293 0.001
R28692 D.n4285 D.n4279 0.001
R28693 D.n4271 D.n4265 0.001
R28694 D.n4257 D.n4251 0.001
R28695 D.n4243 D.n4237 0.001
R28696 D.n4229 D.n4223 0.001
R28697 D.n4215 D.n4209 0.001
R28698 D.n4201 D.n4195 0.001
R28699 D.n4187 D.n4181 0.001
R28700 D.n4173 D.n4167 0.001
R28701 D.n4159 D.n4153 0.001
R28702 D.n4145 D.n4139 0.001
R28703 D.n4131 D.n4125 0.001
R28704 D.n4117 D.n4111 0.001
R28705 D.n4103 D.n4097 0.001
R28706 D.n4089 D.n4083 0.001
R28707 D.n4075 D.n4069 0.001
R28708 D.n4061 D.n4055 0.001
R28709 D.n4047 D.n4041 0.001
R28710 D.n4033 D.n4027 0.001
R28711 D.n4019 D.n4013 0.001
R28712 D.n4005 D.n3999 0.001
R28713 D.n3991 D.n3985 0.001
R28714 D.n3977 D.n3971 0.001
R28715 D.n3963 D.n3957 0.001
R28716 D.n3949 D.n3943 0.001
R28717 D.n3935 D.n3929 0.001
R28718 D.n3921 D.n3915 0.001
R28719 D.n3907 D.n3901 0.001
R28720 D.n4339 D.n4331 0.001
R28721 D.n4353 D.n4347 0.001
R28722 D.n4749 D.n4321 0.001
R28723 D.n4745 D.n4739 0.001
R28724 D.n4731 D.n4725 0.001
R28725 D.n4717 D.n4711 0.001
R28726 D.n4703 D.n4697 0.001
R28727 D.n4689 D.n4683 0.001
R28728 D.n4675 D.n4669 0.001
R28729 D.n4661 D.n4655 0.001
R28730 D.n4647 D.n4641 0.001
R28731 D.n4633 D.n4627 0.001
R28732 D.n4619 D.n4613 0.001
R28733 D.n4605 D.n4599 0.001
R28734 D.n4591 D.n4585 0.001
R28735 D.n4577 D.n4571 0.001
R28736 D.n4563 D.n4557 0.001
R28737 D.n4549 D.n4543 0.001
R28738 D.n4535 D.n4529 0.001
R28739 D.n4521 D.n4515 0.001
R28740 D.n4507 D.n4501 0.001
R28741 D.n4493 D.n4487 0.001
R28742 D.n4479 D.n4473 0.001
R28743 D.n4465 D.n4459 0.001
R28744 D.n4451 D.n4445 0.001
R28745 D.n4437 D.n4431 0.001
R28746 D.n4423 D.n4417 0.001
R28747 D.n4409 D.n4403 0.001
R28748 D.n4395 D.n4389 0.001
R28749 D.n4381 D.n4375 0.001
R28750 D.n4367 D.n4361 0.001
R28751 D.n4771 D.n4763 0.001
R28752 D.n4785 D.n4779 0.001
R28753 D.n5153 D.n4753 0.001
R28754 D.n5149 D.n5143 0.001
R28755 D.n5135 D.n5129 0.001
R28756 D.n5121 D.n5115 0.001
R28757 D.n5107 D.n5101 0.001
R28758 D.n5093 D.n5087 0.001
R28759 D.n5079 D.n5073 0.001
R28760 D.n5065 D.n5059 0.001
R28761 D.n5051 D.n5045 0.001
R28762 D.n5037 D.n5031 0.001
R28763 D.n5023 D.n5017 0.001
R28764 D.n5009 D.n5003 0.001
R28765 D.n4995 D.n4989 0.001
R28766 D.n4981 D.n4975 0.001
R28767 D.n4967 D.n4961 0.001
R28768 D.n4953 D.n4947 0.001
R28769 D.n4939 D.n4933 0.001
R28770 D.n4925 D.n4919 0.001
R28771 D.n4911 D.n4905 0.001
R28772 D.n4897 D.n4891 0.001
R28773 D.n4883 D.n4877 0.001
R28774 D.n4869 D.n4863 0.001
R28775 D.n4855 D.n4849 0.001
R28776 D.n4841 D.n4835 0.001
R28777 D.n4827 D.n4821 0.001
R28778 D.n4813 D.n4807 0.001
R28779 D.n4799 D.n4793 0.001
R28780 D.n5175 D.n5167 0.001
R28781 D.n5189 D.n5183 0.001
R28782 D.n5529 D.n5157 0.001
R28783 D.n5525 D.n5519 0.001
R28784 D.n5511 D.n5505 0.001
R28785 D.n5497 D.n5491 0.001
R28786 D.n5483 D.n5477 0.001
R28787 D.n5469 D.n5463 0.001
R28788 D.n5455 D.n5449 0.001
R28789 D.n5441 D.n5435 0.001
R28790 D.n5427 D.n5421 0.001
R28791 D.n5413 D.n5407 0.001
R28792 D.n5399 D.n5393 0.001
R28793 D.n5385 D.n5379 0.001
R28794 D.n5371 D.n5365 0.001
R28795 D.n5357 D.n5351 0.001
R28796 D.n5343 D.n5337 0.001
R28797 D.n5329 D.n5323 0.001
R28798 D.n5315 D.n5309 0.001
R28799 D.n5301 D.n5295 0.001
R28800 D.n5287 D.n5281 0.001
R28801 D.n5273 D.n5267 0.001
R28802 D.n5259 D.n5253 0.001
R28803 D.n5245 D.n5239 0.001
R28804 D.n5231 D.n5225 0.001
R28805 D.n5217 D.n5211 0.001
R28806 D.n5203 D.n5197 0.001
R28807 D.n5551 D.n5543 0.001
R28808 D.n5565 D.n5559 0.001
R28809 D.n5877 D.n5533 0.001
R28810 D.n5873 D.n5867 0.001
R28811 D.n5859 D.n5853 0.001
R28812 D.n5845 D.n5839 0.001
R28813 D.n5831 D.n5825 0.001
R28814 D.n5817 D.n5811 0.001
R28815 D.n5803 D.n5797 0.001
R28816 D.n5789 D.n5783 0.001
R28817 D.n5775 D.n5769 0.001
R28818 D.n5761 D.n5755 0.001
R28819 D.n5747 D.n5741 0.001
R28820 D.n5733 D.n5727 0.001
R28821 D.n5719 D.n5713 0.001
R28822 D.n5705 D.n5699 0.001
R28823 D.n5691 D.n5685 0.001
R28824 D.n5677 D.n5671 0.001
R28825 D.n5663 D.n5657 0.001
R28826 D.n5649 D.n5643 0.001
R28827 D.n5635 D.n5629 0.001
R28828 D.n5621 D.n5615 0.001
R28829 D.n5607 D.n5601 0.001
R28830 D.n5593 D.n5587 0.001
R28831 D.n5579 D.n5573 0.001
R28832 D.n5899 D.n5891 0.001
R28833 D.n5913 D.n5907 0.001
R28834 D.n6197 D.n5881 0.001
R28835 D.n6193 D.n6187 0.001
R28836 D.n6179 D.n6173 0.001
R28837 D.n6165 D.n6159 0.001
R28838 D.n6151 D.n6145 0.001
R28839 D.n6137 D.n6131 0.001
R28840 D.n6123 D.n6117 0.001
R28841 D.n6109 D.n6103 0.001
R28842 D.n6095 D.n6089 0.001
R28843 D.n6081 D.n6075 0.001
R28844 D.n6067 D.n6061 0.001
R28845 D.n6053 D.n6047 0.001
R28846 D.n6039 D.n6033 0.001
R28847 D.n6025 D.n6019 0.001
R28848 D.n6011 D.n6005 0.001
R28849 D.n5997 D.n5991 0.001
R28850 D.n5983 D.n5977 0.001
R28851 D.n5969 D.n5963 0.001
R28852 D.n5955 D.n5949 0.001
R28853 D.n5941 D.n5935 0.001
R28854 D.n5927 D.n5921 0.001
R28855 D.n6219 D.n6211 0.001
R28856 D.n6233 D.n6227 0.001
R28857 D.n6489 D.n6201 0.001
R28858 D.n6485 D.n6479 0.001
R28859 D.n6471 D.n6465 0.001
R28860 D.n6457 D.n6451 0.001
R28861 D.n6443 D.n6437 0.001
R28862 D.n6429 D.n6423 0.001
R28863 D.n6415 D.n6409 0.001
R28864 D.n6401 D.n6395 0.001
R28865 D.n6387 D.n6381 0.001
R28866 D.n6373 D.n6367 0.001
R28867 D.n6359 D.n6353 0.001
R28868 D.n6345 D.n6339 0.001
R28869 D.n6331 D.n6325 0.001
R28870 D.n6317 D.n6311 0.001
R28871 D.n6303 D.n6297 0.001
R28872 D.n6289 D.n6283 0.001
R28873 D.n6275 D.n6269 0.001
R28874 D.n6261 D.n6255 0.001
R28875 D.n6247 D.n6241 0.001
R28876 D.n6511 D.n6503 0.001
R28877 D.n6525 D.n6519 0.001
R28878 D.n6753 D.n6493 0.001
R28879 D.n6749 D.n6743 0.001
R28880 D.n6735 D.n6729 0.001
R28881 D.n6721 D.n6715 0.001
R28882 D.n6707 D.n6701 0.001
R28883 D.n6693 D.n6687 0.001
R28884 D.n6679 D.n6673 0.001
R28885 D.n6665 D.n6659 0.001
R28886 D.n6651 D.n6645 0.001
R28887 D.n6637 D.n6631 0.001
R28888 D.n6623 D.n6617 0.001
R28889 D.n6609 D.n6603 0.001
R28890 D.n6595 D.n6589 0.001
R28891 D.n6581 D.n6575 0.001
R28892 D.n6567 D.n6561 0.001
R28893 D.n6553 D.n6547 0.001
R28894 D.n6539 D.n6533 0.001
R28895 D.n6775 D.n6767 0.001
R28896 D.n6789 D.n6783 0.001
R28897 D.n6989 D.n6757 0.001
R28898 D.n6985 D.n6979 0.001
R28899 D.n6971 D.n6965 0.001
R28900 D.n6957 D.n6951 0.001
R28901 D.n6943 D.n6937 0.001
R28902 D.n6929 D.n6923 0.001
R28903 D.n6915 D.n6909 0.001
R28904 D.n6901 D.n6895 0.001
R28905 D.n6887 D.n6881 0.001
R28906 D.n6873 D.n6867 0.001
R28907 D.n6859 D.n6853 0.001
R28908 D.n6845 D.n6839 0.001
R28909 D.n6831 D.n6825 0.001
R28910 D.n6817 D.n6811 0.001
R28911 D.n6803 D.n6797 0.001
R28912 D.n7011 D.n7003 0.001
R28913 D.n7025 D.n7019 0.001
R28914 D.n7197 D.n6993 0.001
R28915 D.n7193 D.n7187 0.001
R28916 D.n7179 D.n7173 0.001
R28917 D.n7165 D.n7159 0.001
R28918 D.n7151 D.n7145 0.001
R28919 D.n7137 D.n7131 0.001
R28920 D.n7123 D.n7117 0.001
R28921 D.n7109 D.n7103 0.001
R28922 D.n7095 D.n7089 0.001
R28923 D.n7081 D.n7075 0.001
R28924 D.n7067 D.n7061 0.001
R28925 D.n7053 D.n7047 0.001
R28926 D.n7039 D.n7033 0.001
R28927 D.n7219 D.n7211 0.001
R28928 D.n7233 D.n7227 0.001
R28929 D.n7377 D.n7201 0.001
R28930 D.n7373 D.n7367 0.001
R28931 D.n7359 D.n7353 0.001
R28932 D.n7345 D.n7339 0.001
R28933 D.n7331 D.n7325 0.001
R28934 D.n7317 D.n7311 0.001
R28935 D.n7303 D.n7297 0.001
R28936 D.n7289 D.n7283 0.001
R28937 D.n7275 D.n7269 0.001
R28938 D.n7261 D.n7255 0.001
R28939 D.n7247 D.n7241 0.001
R28940 D.n7399 D.n7391 0.001
R28941 D.n7413 D.n7407 0.001
R28942 D.n7529 D.n7381 0.001
R28943 D.n7525 D.n7519 0.001
R28944 D.n7511 D.n7505 0.001
R28945 D.n7497 D.n7491 0.001
R28946 D.n7483 D.n7477 0.001
R28947 D.n7469 D.n7463 0.001
R28948 D.n7455 D.n7449 0.001
R28949 D.n7441 D.n7435 0.001
R28950 D.n7427 D.n7421 0.001
R28951 D.n7551 D.n7543 0.001
R28952 D.n7565 D.n7559 0.001
R28953 D.n7653 D.n7533 0.001
R28954 D.n7649 D.n7643 0.001
R28955 D.n7635 D.n7629 0.001
R28956 D.n7621 D.n7615 0.001
R28957 D.n7607 D.n7601 0.001
R28958 D.n7593 D.n7587 0.001
R28959 D.n7579 D.n7573 0.001
R28960 D.n7675 D.n7667 0.001
R28961 D.n7689 D.n7683 0.001
R28962 D.n7749 D.n7657 0.001
R28963 D.n7745 D.n7739 0.001
R28964 D.n7731 D.n7725 0.001
R28965 D.n7717 D.n7711 0.001
R28966 D.n7703 D.n7697 0.001
R28967 D.n7770 D.n7762 0.001
R28968 D.n7784 D.n7778 0.001
R28969 D.n7816 D.n7752 0.001
R28970 D.n7814 D.n7806 0.001
R28971 D.n7798 D.n7792 0.001
R28972 D.n7842 D.n7837 0.001
R28973 D.n7832 D.n7827 0.001
R28974 D.n453 D.n448 0.001
R28975 D.n444 D.n439 0.001
R28976 D.n47 D.n30 0.001
R28977 D.n7962 D.n7957 0.001
R28978 D.n7952 D.n7942 0.001
R28979 D.n14067 D.n14062 0.001
R28980 D.n14049 D.n14044 0.001
R28981 D.n14031 D.n14026 0.001
R28982 D.n14013 D.n14008 0.001
R28983 D.n13995 D.n13990 0.001
R28984 D.n13977 D.n13972 0.001
R28985 D.n13959 D.n13954 0.001
R28986 D.n13941 D.n13936 0.001
R28987 D.n13923 D.n13918 0.001
R28988 D.n13905 D.n13900 0.001
R28989 D.n13887 D.n13882 0.001
R28990 D.n13869 D.n13864 0.001
R28991 D.n13851 D.n13846 0.001
R28992 D.n13833 D.n13828 0.001
R28993 D.n13815 D.n13810 0.001
R28994 D.n13797 D.n13792 0.001
R28995 D.n13779 D.n13774 0.001
R28996 D.n13761 D.n13756 0.001
R28997 D.n13743 D.n13738 0.001
R28998 D.n13725 D.n13720 0.001
R28999 D.n13707 D.n13702 0.001
R29000 D.n13689 D.n13683 0.001
R29001 D.n13698 D.n13693 0.001
R29002 D.n13716 D.n13711 0.001
R29003 D.n13734 D.n13729 0.001
R29004 D.n13752 D.n13747 0.001
R29005 D.n13770 D.n13765 0.001
R29006 D.n13788 D.n13783 0.001
R29007 D.n13806 D.n13801 0.001
R29008 D.n13824 D.n13819 0.001
R29009 D.n13842 D.n13837 0.001
R29010 D.n13860 D.n13855 0.001
R29011 D.n13878 D.n13873 0.001
R29012 D.n13896 D.n13891 0.001
R29013 D.n13914 D.n13909 0.001
R29014 D.n13932 D.n13927 0.001
R29015 D.n13950 D.n13945 0.001
R29016 D.n13968 D.n13963 0.001
R29017 D.n13986 D.n13981 0.001
R29018 D.n14004 D.n13999 0.001
R29019 D.n14022 D.n14017 0.001
R29020 D.n14040 D.n14035 0.001
R29021 D.n14058 D.n14053 0.001
R29022 D.n14081 D.n14075 0.001
R29023 D.n13212 D.n13208 0.001
R29024 D.n13232 D.n13228 0.001
R29025 D.n13252 D.n13248 0.001
R29026 D.n13272 D.n13268 0.001
R29027 D.n13292 D.n13288 0.001
R29028 D.n13312 D.n13308 0.001
R29029 D.n13332 D.n13328 0.001
R29030 D.n13352 D.n13348 0.001
R29031 D.n13372 D.n13368 0.001
R29032 D.n13392 D.n13388 0.001
R29033 D.n13412 D.n13408 0.001
R29034 D.n13432 D.n13428 0.001
R29035 D.n13452 D.n13448 0.001
R29036 D.n13472 D.n13468 0.001
R29037 D.n13492 D.n13488 0.001
R29038 D.n13512 D.n13508 0.001
R29039 D.n13532 D.n13528 0.001
R29040 D.n13552 D.n13548 0.001
R29041 D.n13572 D.n13568 0.001
R29042 D.n13592 D.n13588 0.001
R29043 D.n13612 D.n13608 0.001
R29044 D.n13602 D.n13597 0.001
R29045 D.n13582 D.n13577 0.001
R29046 D.n13562 D.n13557 0.001
R29047 D.n13542 D.n13537 0.001
R29048 D.n13522 D.n13517 0.001
R29049 D.n13502 D.n13497 0.001
R29050 D.n13482 D.n13477 0.001
R29051 D.n13462 D.n13457 0.001
R29052 D.n13442 D.n13437 0.001
R29053 D.n13422 D.n13417 0.001
R29054 D.n13402 D.n13397 0.001
R29055 D.n13382 D.n13377 0.001
R29056 D.n13362 D.n13357 0.001
R29057 D.n13342 D.n13337 0.001
R29058 D.n13322 D.n13317 0.001
R29059 D.n13302 D.n13297 0.001
R29060 D.n13282 D.n13277 0.001
R29061 D.n13262 D.n13257 0.001
R29062 D.n13242 D.n13237 0.001
R29063 D.n13222 D.n13217 0.001
R29064 D.n13202 D.n13192 0.001
R29065 D.n13104 D.n13099 0.001
R29066 D.n13086 D.n13081 0.001
R29067 D.n13068 D.n13063 0.001
R29068 D.n13050 D.n13045 0.001
R29069 D.n13032 D.n13027 0.001
R29070 D.n13014 D.n13009 0.001
R29071 D.n12996 D.n12991 0.001
R29072 D.n12978 D.n12973 0.001
R29073 D.n12960 D.n12955 0.001
R29074 D.n12942 D.n12937 0.001
R29075 D.n12924 D.n12919 0.001
R29076 D.n12906 D.n12901 0.001
R29077 D.n12888 D.n12883 0.001
R29078 D.n12870 D.n12865 0.001
R29079 D.n12852 D.n12847 0.001
R29080 D.n12834 D.n12829 0.001
R29081 D.n12816 D.n12811 0.001
R29082 D.n12798 D.n12793 0.001
R29083 D.n12780 D.n12775 0.001
R29084 D.n12762 D.n12756 0.001
R29085 D.n12771 D.n12766 0.001
R29086 D.n12789 D.n12784 0.001
R29087 D.n12807 D.n12802 0.001
R29088 D.n12825 D.n12820 0.001
R29089 D.n12843 D.n12838 0.001
R29090 D.n12861 D.n12856 0.001
R29091 D.n12879 D.n12874 0.001
R29092 D.n12897 D.n12892 0.001
R29093 D.n12915 D.n12910 0.001
R29094 D.n12933 D.n12928 0.001
R29095 D.n12951 D.n12946 0.001
R29096 D.n12969 D.n12964 0.001
R29097 D.n12987 D.n12982 0.001
R29098 D.n13005 D.n13000 0.001
R29099 D.n13023 D.n13018 0.001
R29100 D.n13041 D.n13036 0.001
R29101 D.n13059 D.n13054 0.001
R29102 D.n13077 D.n13072 0.001
R29103 D.n13095 D.n13090 0.001
R29104 D.n13117 D.n13111 0.001
R29105 D.n12329 D.n12325 0.001
R29106 D.n12349 D.n12345 0.001
R29107 D.n12369 D.n12365 0.001
R29108 D.n12389 D.n12385 0.001
R29109 D.n12409 D.n12405 0.001
R29110 D.n12429 D.n12425 0.001
R29111 D.n12449 D.n12445 0.001
R29112 D.n12469 D.n12465 0.001
R29113 D.n12489 D.n12485 0.001
R29114 D.n12509 D.n12505 0.001
R29115 D.n12529 D.n12525 0.001
R29116 D.n12549 D.n12545 0.001
R29117 D.n12569 D.n12565 0.001
R29118 D.n12589 D.n12585 0.001
R29119 D.n12609 D.n12605 0.001
R29120 D.n12629 D.n12625 0.001
R29121 D.n12649 D.n12645 0.001
R29122 D.n12669 D.n12665 0.001
R29123 D.n12689 D.n12685 0.001
R29124 D.n12679 D.n12674 0.001
R29125 D.n12659 D.n12654 0.001
R29126 D.n12639 D.n12634 0.001
R29127 D.n12619 D.n12614 0.001
R29128 D.n12599 D.n12594 0.001
R29129 D.n12579 D.n12574 0.001
R29130 D.n12559 D.n12554 0.001
R29131 D.n12539 D.n12534 0.001
R29132 D.n12519 D.n12514 0.001
R29133 D.n12499 D.n12494 0.001
R29134 D.n12479 D.n12474 0.001
R29135 D.n12459 D.n12454 0.001
R29136 D.n12439 D.n12434 0.001
R29137 D.n12419 D.n12414 0.001
R29138 D.n12399 D.n12394 0.001
R29139 D.n12379 D.n12374 0.001
R29140 D.n12359 D.n12354 0.001
R29141 D.n12339 D.n12334 0.001
R29142 D.n12319 D.n12309 0.001
R29143 D.n12219 D.n12214 0.001
R29144 D.n12201 D.n12196 0.001
R29145 D.n12183 D.n12178 0.001
R29146 D.n12165 D.n12160 0.001
R29147 D.n12147 D.n12142 0.001
R29148 D.n12129 D.n12124 0.001
R29149 D.n12111 D.n12106 0.001
R29150 D.n12093 D.n12088 0.001
R29151 D.n12075 D.n12070 0.001
R29152 D.n12057 D.n12052 0.001
R29153 D.n12039 D.n12034 0.001
R29154 D.n12021 D.n12016 0.001
R29155 D.n12003 D.n11998 0.001
R29156 D.n11985 D.n11980 0.001
R29157 D.n11967 D.n11962 0.001
R29158 D.n11949 D.n11944 0.001
R29159 D.n11931 D.n11926 0.001
R29160 D.n11913 D.n11907 0.001
R29161 D.n11922 D.n11917 0.001
R29162 D.n11940 D.n11935 0.001
R29163 D.n11958 D.n11953 0.001
R29164 D.n11976 D.n11971 0.001
R29165 D.n11994 D.n11989 0.001
R29166 D.n12012 D.n12007 0.001
R29167 D.n12030 D.n12025 0.001
R29168 D.n12048 D.n12043 0.001
R29169 D.n12066 D.n12061 0.001
R29170 D.n12084 D.n12079 0.001
R29171 D.n12102 D.n12097 0.001
R29172 D.n12120 D.n12115 0.001
R29173 D.n12138 D.n12133 0.001
R29174 D.n12156 D.n12151 0.001
R29175 D.n12174 D.n12169 0.001
R29176 D.n12192 D.n12187 0.001
R29177 D.n12210 D.n12205 0.001
R29178 D.n12232 D.n12227 0.001
R29179 D.n11520 D.n11516 0.001
R29180 D.n11540 D.n11536 0.001
R29181 D.n11560 D.n11556 0.001
R29182 D.n11580 D.n11576 0.001
R29183 D.n11600 D.n11596 0.001
R29184 D.n11620 D.n11616 0.001
R29185 D.n11640 D.n11636 0.001
R29186 D.n11660 D.n11656 0.001
R29187 D.n11680 D.n11676 0.001
R29188 D.n11700 D.n11696 0.001
R29189 D.n11720 D.n11716 0.001
R29190 D.n11740 D.n11736 0.001
R29191 D.n11760 D.n11756 0.001
R29192 D.n11780 D.n11776 0.001
R29193 D.n11800 D.n11796 0.001
R29194 D.n11820 D.n11816 0.001
R29195 D.n11840 D.n11836 0.001
R29196 D.n11830 D.n11825 0.001
R29197 D.n11810 D.n11805 0.001
R29198 D.n11790 D.n11785 0.001
R29199 D.n11770 D.n11765 0.001
R29200 D.n11750 D.n11745 0.001
R29201 D.n11730 D.n11725 0.001
R29202 D.n11710 D.n11705 0.001
R29203 D.n11690 D.n11685 0.001
R29204 D.n11670 D.n11665 0.001
R29205 D.n11650 D.n11645 0.001
R29206 D.n11630 D.n11625 0.001
R29207 D.n11610 D.n11605 0.001
R29208 D.n11590 D.n11585 0.001
R29209 D.n11570 D.n11565 0.001
R29210 D.n11550 D.n11545 0.001
R29211 D.n11530 D.n11525 0.001
R29212 D.n11510 D.n11502 0.001
R29213 D.n11420 D.n11415 0.001
R29214 D.n11402 D.n11397 0.001
R29215 D.n11384 D.n11379 0.001
R29216 D.n11366 D.n11361 0.001
R29217 D.n11348 D.n11343 0.001
R29218 D.n11330 D.n11325 0.001
R29219 D.n11312 D.n11307 0.001
R29220 D.n11294 D.n11289 0.001
R29221 D.n11276 D.n11271 0.001
R29222 D.n11258 D.n11253 0.001
R29223 D.n11240 D.n11235 0.001
R29224 D.n11222 D.n11217 0.001
R29225 D.n11204 D.n11199 0.001
R29226 D.n11186 D.n11181 0.001
R29227 D.n11168 D.n11163 0.001
R29228 D.n11150 D.n11144 0.001
R29229 D.n11159 D.n11154 0.001
R29230 D.n11177 D.n11172 0.001
R29231 D.n11195 D.n11190 0.001
R29232 D.n11213 D.n11208 0.001
R29233 D.n11231 D.n11226 0.001
R29234 D.n11249 D.n11244 0.001
R29235 D.n11267 D.n11262 0.001
R29236 D.n11285 D.n11280 0.001
R29237 D.n11303 D.n11298 0.001
R29238 D.n11321 D.n11316 0.001
R29239 D.n11339 D.n11334 0.001
R29240 D.n11357 D.n11352 0.001
R29241 D.n11375 D.n11370 0.001
R29242 D.n11393 D.n11388 0.001
R29243 D.n11411 D.n11406 0.001
R29244 D.n11433 D.n11428 0.001
R29245 D.n10797 D.n10793 0.001
R29246 D.n10817 D.n10813 0.001
R29247 D.n10837 D.n10833 0.001
R29248 D.n10857 D.n10853 0.001
R29249 D.n10877 D.n10873 0.001
R29250 D.n10897 D.n10893 0.001
R29251 D.n10917 D.n10913 0.001
R29252 D.n10937 D.n10933 0.001
R29253 D.n10957 D.n10953 0.001
R29254 D.n10977 D.n10973 0.001
R29255 D.n10997 D.n10993 0.001
R29256 D.n11017 D.n11013 0.001
R29257 D.n11037 D.n11033 0.001
R29258 D.n11057 D.n11053 0.001
R29259 D.n11077 D.n11073 0.001
R29260 D.n11067 D.n11062 0.001
R29261 D.n11047 D.n11042 0.001
R29262 D.n11027 D.n11022 0.001
R29263 D.n11007 D.n11002 0.001
R29264 D.n10987 D.n10982 0.001
R29265 D.n10967 D.n10962 0.001
R29266 D.n10947 D.n10942 0.001
R29267 D.n10927 D.n10922 0.001
R29268 D.n10907 D.n10902 0.001
R29269 D.n10887 D.n10882 0.001
R29270 D.n10867 D.n10862 0.001
R29271 D.n10847 D.n10842 0.001
R29272 D.n10827 D.n10822 0.001
R29273 D.n10807 D.n10802 0.001
R29274 D.n10787 D.n10779 0.001
R29275 D.n10701 D.n10696 0.001
R29276 D.n10683 D.n10678 0.001
R29277 D.n10665 D.n10660 0.001
R29278 D.n10647 D.n10642 0.001
R29279 D.n10629 D.n10624 0.001
R29280 D.n10611 D.n10606 0.001
R29281 D.n10593 D.n10588 0.001
R29282 D.n10575 D.n10570 0.001
R29283 D.n10557 D.n10552 0.001
R29284 D.n10539 D.n10534 0.001
R29285 D.n10521 D.n10516 0.001
R29286 D.n10503 D.n10498 0.001
R29287 D.n10485 D.n10480 0.001
R29288 D.n10467 D.n10461 0.001
R29289 D.n10476 D.n10471 0.001
R29290 D.n10494 D.n10489 0.001
R29291 D.n10512 D.n10507 0.001
R29292 D.n10530 D.n10525 0.001
R29293 D.n10548 D.n10543 0.001
R29294 D.n10566 D.n10561 0.001
R29295 D.n10584 D.n10579 0.001
R29296 D.n10602 D.n10597 0.001
R29297 D.n10620 D.n10615 0.001
R29298 D.n10638 D.n10633 0.001
R29299 D.n10656 D.n10651 0.001
R29300 D.n10674 D.n10669 0.001
R29301 D.n10692 D.n10687 0.001
R29302 D.n10714 D.n10709 0.001
R29303 D.n10154 D.n10150 0.001
R29304 D.n10174 D.n10170 0.001
R29305 D.n10194 D.n10190 0.001
R29306 D.n10214 D.n10210 0.001
R29307 D.n10234 D.n10230 0.001
R29308 D.n10254 D.n10250 0.001
R29309 D.n10274 D.n10270 0.001
R29310 D.n10294 D.n10290 0.001
R29311 D.n10314 D.n10310 0.001
R29312 D.n10334 D.n10330 0.001
R29313 D.n10354 D.n10350 0.001
R29314 D.n10374 D.n10370 0.001
R29315 D.n10394 D.n10390 0.001
R29316 D.n10384 D.n10379 0.001
R29317 D.n10364 D.n10359 0.001
R29318 D.n10344 D.n10339 0.001
R29319 D.n10324 D.n10319 0.001
R29320 D.n10304 D.n10299 0.001
R29321 D.n10284 D.n10279 0.001
R29322 D.n10264 D.n10259 0.001
R29323 D.n10244 D.n10239 0.001
R29324 D.n10224 D.n10219 0.001
R29325 D.n10204 D.n10199 0.001
R29326 D.n10184 D.n10179 0.001
R29327 D.n10164 D.n10159 0.001
R29328 D.n10144 D.n10134 0.001
R29329 D.n10062 D.n10057 0.001
R29330 D.n10044 D.n10039 0.001
R29331 D.n10026 D.n10021 0.001
R29332 D.n10008 D.n10003 0.001
R29333 D.n9990 D.n9985 0.001
R29334 D.n9972 D.n9967 0.001
R29335 D.n9954 D.n9949 0.001
R29336 D.n9936 D.n9931 0.001
R29337 D.n9918 D.n9913 0.001
R29338 D.n9900 D.n9895 0.001
R29339 D.n9882 D.n9877 0.001
R29340 D.n9864 D.n9858 0.001
R29341 D.n9873 D.n9868 0.001
R29342 D.n9891 D.n9886 0.001
R29343 D.n9909 D.n9904 0.001
R29344 D.n9927 D.n9922 0.001
R29345 D.n9945 D.n9940 0.001
R29346 D.n9963 D.n9958 0.001
R29347 D.n9981 D.n9976 0.001
R29348 D.n9999 D.n9994 0.001
R29349 D.n10017 D.n10012 0.001
R29350 D.n10035 D.n10030 0.001
R29351 D.n10053 D.n10048 0.001
R29352 D.n10075 D.n10069 0.001
R29353 D.n9591 D.n9587 0.001
R29354 D.n9611 D.n9607 0.001
R29355 D.n9631 D.n9627 0.001
R29356 D.n9651 D.n9647 0.001
R29357 D.n9671 D.n9667 0.001
R29358 D.n9691 D.n9687 0.001
R29359 D.n9711 D.n9707 0.001
R29360 D.n9731 D.n9727 0.001
R29361 D.n9751 D.n9747 0.001
R29362 D.n9771 D.n9767 0.001
R29363 D.n9791 D.n9787 0.001
R29364 D.n9781 D.n9776 0.001
R29365 D.n9761 D.n9756 0.001
R29366 D.n9741 D.n9736 0.001
R29367 D.n9721 D.n9716 0.001
R29368 D.n9701 D.n9696 0.001
R29369 D.n9681 D.n9676 0.001
R29370 D.n9661 D.n9656 0.001
R29371 D.n9641 D.n9636 0.001
R29372 D.n9621 D.n9616 0.001
R29373 D.n9601 D.n9596 0.001
R29374 D.n9581 D.n9571 0.001
R29375 D.n9497 D.n9492 0.001
R29376 D.n9479 D.n9474 0.001
R29377 D.n9461 D.n9456 0.001
R29378 D.n9443 D.n9438 0.001
R29379 D.n9425 D.n9420 0.001
R29380 D.n9407 D.n9402 0.001
R29381 D.n9389 D.n9384 0.001
R29382 D.n9371 D.n9366 0.001
R29383 D.n9353 D.n9348 0.001
R29384 D.n9335 D.n9329 0.001
R29385 D.n9344 D.n9339 0.001
R29386 D.n9362 D.n9357 0.001
R29387 D.n9380 D.n9375 0.001
R29388 D.n9398 D.n9393 0.001
R29389 D.n9416 D.n9411 0.001
R29390 D.n9434 D.n9429 0.001
R29391 D.n9452 D.n9447 0.001
R29392 D.n9470 D.n9465 0.001
R29393 D.n9488 D.n9483 0.001
R29394 D.n9510 D.n9505 0.001
R29395 D.n9102 D.n9098 0.001
R29396 D.n9122 D.n9118 0.001
R29397 D.n9142 D.n9138 0.001
R29398 D.n9162 D.n9158 0.001
R29399 D.n9182 D.n9178 0.001
R29400 D.n9202 D.n9198 0.001
R29401 D.n9222 D.n9218 0.001
R29402 D.n9242 D.n9238 0.001
R29403 D.n9262 D.n9258 0.001
R29404 D.n9252 D.n9247 0.001
R29405 D.n9232 D.n9227 0.001
R29406 D.n9212 D.n9207 0.001
R29407 D.n9192 D.n9187 0.001
R29408 D.n9172 D.n9167 0.001
R29409 D.n9152 D.n9147 0.001
R29410 D.n9132 D.n9127 0.001
R29411 D.n9112 D.n9107 0.001
R29412 D.n9092 D.n9084 0.001
R29413 D.n9018 D.n9013 0.001
R29414 D.n9000 D.n8995 0.001
R29415 D.n8982 D.n8977 0.001
R29416 D.n8964 D.n8959 0.001
R29417 D.n8946 D.n8941 0.001
R29418 D.n8928 D.n8923 0.001
R29419 D.n8910 D.n8905 0.001
R29420 D.n8892 D.n8886 0.001
R29421 D.n8901 D.n8896 0.001
R29422 D.n8919 D.n8914 0.001
R29423 D.n8937 D.n8932 0.001
R29424 D.n8955 D.n8950 0.001
R29425 D.n8973 D.n8968 0.001
R29426 D.n8991 D.n8986 0.001
R29427 D.n9009 D.n9004 0.001
R29428 D.n9031 D.n9026 0.001
R29429 D.n8699 D.n8695 0.001
R29430 D.n8719 D.n8715 0.001
R29431 D.n8739 D.n8735 0.001
R29432 D.n8759 D.n8755 0.001
R29433 D.n8779 D.n8775 0.001
R29434 D.n8799 D.n8795 0.001
R29435 D.n8819 D.n8815 0.001
R29436 D.n8809 D.n8804 0.001
R29437 D.n8789 D.n8784 0.001
R29438 D.n8769 D.n8764 0.001
R29439 D.n8749 D.n8744 0.001
R29440 D.n8729 D.n8724 0.001
R29441 D.n8709 D.n8704 0.001
R29442 D.n8689 D.n8679 0.001
R29443 D.n8619 D.n8614 0.001
R29444 D.n8601 D.n8596 0.001
R29445 D.n8583 D.n8578 0.001
R29446 D.n8565 D.n8560 0.001
R29447 D.n8547 D.n8542 0.001
R29448 D.n8529 D.n8523 0.001
R29449 D.n8538 D.n8533 0.001
R29450 D.n8556 D.n8551 0.001
R29451 D.n8574 D.n8569 0.001
R29452 D.n8592 D.n8587 0.001
R29453 D.n8610 D.n8605 0.001
R29454 D.n8632 D.n8626 0.001
R29455 D.n8376 D.n8372 0.001
R29456 D.n8396 D.n8392 0.001
R29457 D.n8416 D.n8412 0.001
R29458 D.n8436 D.n8432 0.001
R29459 D.n8456 D.n8452 0.001
R29460 D.n8446 D.n8441 0.001
R29461 D.n8426 D.n8421 0.001
R29462 D.n8406 D.n8401 0.001
R29463 D.n8386 D.n8381 0.001
R29464 D.n8366 D.n8356 0.001
R29465 D.n8294 D.n8289 0.001
R29466 D.n8276 D.n8271 0.001
R29467 D.n8258 D.n8253 0.001
R29468 D.n8240 D.n8234 0.001
R29469 D.n8249 D.n8244 0.001
R29470 D.n8267 D.n8262 0.001
R29471 D.n8285 D.n8280 0.001
R29472 D.n8307 D.n8302 0.001
R29473 D.n8127 D.n8123 0.001
R29474 D.n8147 D.n8143 0.001
R29475 D.n8167 D.n8163 0.001
R29476 D.n8157 D.n8152 0.001
R29477 D.n8137 D.n8132 0.001
R29478 D.n8117 D.n8109 0.001
R29479 D.n8055 D.n8050 0.001
R29480 D.n8037 D.n8031 0.001
R29481 D.n8046 D.n8041 0.001
R29482 D.n8068 D.n8063 0.001
R29483 D.n57 D.n52 0.001
R29484 D.n66 D.n61 0.001
R29485 D.n75 D.n70 0.001
R29486 D.n84 D.n79 0.001
R29487 D.n93 D.n88 0.001
R29488 D.n102 D.n97 0.001
R29489 D.n111 D.n106 0.001
R29490 D.n120 D.n115 0.001
R29491 D.n129 D.n124 0.001
R29492 D.n138 D.n133 0.001
R29493 D.n147 D.n142 0.001
R29494 D.n156 D.n151 0.001
R29495 D.n165 D.n160 0.001
R29496 D.n174 D.n169 0.001
R29497 D.n183 D.n178 0.001
R29498 D.n192 D.n187 0.001
R29499 D.n201 D.n196 0.001
R29500 D.n210 D.n205 0.001
R29501 D.n219 D.n214 0.001
R29502 D.n228 D.n223 0.001
R29503 D.n237 D.n232 0.001
R29504 D.n246 D.n241 0.001
R29505 D.n255 D.n250 0.001
R29506 D.n264 D.n259 0.001
R29507 D.n273 D.n268 0.001
R29508 D.n282 D.n277 0.001
R29509 D.n291 D.n286 0.001
R29510 D.n300 D.n295 0.001
R29511 D.n309 D.n304 0.001
R29512 D.n318 D.n313 0.001
R29513 D.n327 D.n322 0.001
R29514 D.n336 D.n331 0.001
R29515 D.n345 D.n340 0.001
R29516 D.n354 D.n349 0.001
R29517 D.n363 D.n358 0.001
R29518 D.n372 D.n367 0.001
R29519 D.n381 D.n376 0.001
R29520 D.n390 D.n385 0.001
R29521 D.n399 D.n394 0.001
R29522 D.n408 D.n403 0.001
R29523 D.n417 D.n412 0.001
R29524 D.n426 D.n421 0.001
R29525 D.n435 D.n430 0.001
R29526 D.n535 D.n524 0.001
R29527 D.n549 D.n540 0.001
R29528 D.n1137 D.n1128 0.001
R29529 D.n1123 D.n1114 0.001
R29530 D.n1109 D.n1100 0.001
R29531 D.n1095 D.n1086 0.001
R29532 D.n1081 D.n1072 0.001
R29533 D.n1067 D.n1058 0.001
R29534 D.n1053 D.n1044 0.001
R29535 D.n1039 D.n1030 0.001
R29536 D.n1025 D.n1016 0.001
R29537 D.n1011 D.n1002 0.001
R29538 D.n997 D.n988 0.001
R29539 D.n983 D.n974 0.001
R29540 D.n969 D.n960 0.001
R29541 D.n955 D.n946 0.001
R29542 D.n941 D.n932 0.001
R29543 D.n927 D.n918 0.001
R29544 D.n913 D.n904 0.001
R29545 D.n899 D.n890 0.001
R29546 D.n885 D.n876 0.001
R29547 D.n871 D.n862 0.001
R29548 D.n857 D.n848 0.001
R29549 D.n843 D.n834 0.001
R29550 D.n829 D.n820 0.001
R29551 D.n815 D.n806 0.001
R29552 D.n801 D.n792 0.001
R29553 D.n787 D.n778 0.001
R29554 D.n773 D.n764 0.001
R29555 D.n759 D.n750 0.001
R29556 D.n745 D.n736 0.001
R29557 D.n731 D.n722 0.001
R29558 D.n717 D.n708 0.001
R29559 D.n703 D.n694 0.001
R29560 D.n689 D.n680 0.001
R29561 D.n675 D.n666 0.001
R29562 D.n661 D.n652 0.001
R29563 D.n647 D.n638 0.001
R29564 D.n633 D.n624 0.001
R29565 D.n619 D.n610 0.001
R29566 D.n605 D.n596 0.001
R29567 D.n591 D.n582 0.001
R29568 D.n577 D.n568 0.001
R29569 D.n563 D.n554 0.001
R29570 D.n1162 D.n1151 0.001
R29571 D.n1176 D.n1167 0.001
R29572 D.n1736 D.n1727 0.001
R29573 D.n1722 D.n1713 0.001
R29574 D.n1708 D.n1699 0.001
R29575 D.n1694 D.n1685 0.001
R29576 D.n1680 D.n1671 0.001
R29577 D.n1666 D.n1657 0.001
R29578 D.n1652 D.n1643 0.001
R29579 D.n1638 D.n1629 0.001
R29580 D.n1624 D.n1615 0.001
R29581 D.n1610 D.n1601 0.001
R29582 D.n1596 D.n1587 0.001
R29583 D.n1582 D.n1573 0.001
R29584 D.n1568 D.n1559 0.001
R29585 D.n1554 D.n1545 0.001
R29586 D.n1540 D.n1531 0.001
R29587 D.n1526 D.n1517 0.001
R29588 D.n1512 D.n1503 0.001
R29589 D.n1498 D.n1489 0.001
R29590 D.n1484 D.n1475 0.001
R29591 D.n1470 D.n1461 0.001
R29592 D.n1456 D.n1447 0.001
R29593 D.n1442 D.n1433 0.001
R29594 D.n1428 D.n1419 0.001
R29595 D.n1414 D.n1405 0.001
R29596 D.n1400 D.n1391 0.001
R29597 D.n1386 D.n1377 0.001
R29598 D.n1372 D.n1363 0.001
R29599 D.n1358 D.n1349 0.001
R29600 D.n1344 D.n1335 0.001
R29601 D.n1330 D.n1321 0.001
R29602 D.n1316 D.n1307 0.001
R29603 D.n1302 D.n1293 0.001
R29604 D.n1288 D.n1279 0.001
R29605 D.n1274 D.n1265 0.001
R29606 D.n1260 D.n1251 0.001
R29607 D.n1246 D.n1237 0.001
R29608 D.n1232 D.n1223 0.001
R29609 D.n1218 D.n1209 0.001
R29610 D.n1204 D.n1195 0.001
R29611 D.n1190 D.n1181 0.001
R29612 D.n1761 D.n1750 0.001
R29613 D.n1775 D.n1766 0.001
R29614 D.n2307 D.n2298 0.001
R29615 D.n2293 D.n2284 0.001
R29616 D.n2279 D.n2270 0.001
R29617 D.n2265 D.n2256 0.001
R29618 D.n2251 D.n2242 0.001
R29619 D.n2237 D.n2228 0.001
R29620 D.n2223 D.n2214 0.001
R29621 D.n2209 D.n2200 0.001
R29622 D.n2195 D.n2186 0.001
R29623 D.n2181 D.n2172 0.001
R29624 D.n2167 D.n2158 0.001
R29625 D.n2153 D.n2144 0.001
R29626 D.n2139 D.n2130 0.001
R29627 D.n2125 D.n2116 0.001
R29628 D.n2111 D.n2102 0.001
R29629 D.n2097 D.n2088 0.001
R29630 D.n2083 D.n2074 0.001
R29631 D.n2069 D.n2060 0.001
R29632 D.n2055 D.n2046 0.001
R29633 D.n2041 D.n2032 0.001
R29634 D.n2027 D.n2018 0.001
R29635 D.n2013 D.n2004 0.001
R29636 D.n1999 D.n1990 0.001
R29637 D.n1985 D.n1976 0.001
R29638 D.n1971 D.n1962 0.001
R29639 D.n1957 D.n1948 0.001
R29640 D.n1943 D.n1934 0.001
R29641 D.n1929 D.n1920 0.001
R29642 D.n1915 D.n1906 0.001
R29643 D.n1901 D.n1892 0.001
R29644 D.n1887 D.n1878 0.001
R29645 D.n1873 D.n1864 0.001
R29646 D.n1859 D.n1850 0.001
R29647 D.n1845 D.n1836 0.001
R29648 D.n1831 D.n1822 0.001
R29649 D.n1817 D.n1808 0.001
R29650 D.n1803 D.n1794 0.001
R29651 D.n1789 D.n1780 0.001
R29652 D.n2332 D.n2321 0.001
R29653 D.n2346 D.n2337 0.001
R29654 D.n2850 D.n2841 0.001
R29655 D.n2836 D.n2827 0.001
R29656 D.n2822 D.n2813 0.001
R29657 D.n2808 D.n2799 0.001
R29658 D.n2794 D.n2785 0.001
R29659 D.n2780 D.n2771 0.001
R29660 D.n2766 D.n2757 0.001
R29661 D.n2752 D.n2743 0.001
R29662 D.n2738 D.n2729 0.001
R29663 D.n2724 D.n2715 0.001
R29664 D.n2710 D.n2701 0.001
R29665 D.n2696 D.n2687 0.001
R29666 D.n2682 D.n2673 0.001
R29667 D.n2668 D.n2659 0.001
R29668 D.n2654 D.n2645 0.001
R29669 D.n2640 D.n2631 0.001
R29670 D.n2626 D.n2617 0.001
R29671 D.n2612 D.n2603 0.001
R29672 D.n2598 D.n2589 0.001
R29673 D.n2584 D.n2575 0.001
R29674 D.n2570 D.n2561 0.001
R29675 D.n2556 D.n2547 0.001
R29676 D.n2542 D.n2533 0.001
R29677 D.n2528 D.n2519 0.001
R29678 D.n2514 D.n2505 0.001
R29679 D.n2500 D.n2491 0.001
R29680 D.n2486 D.n2477 0.001
R29681 D.n2472 D.n2463 0.001
R29682 D.n2458 D.n2449 0.001
R29683 D.n2444 D.n2435 0.001
R29684 D.n2430 D.n2421 0.001
R29685 D.n2416 D.n2407 0.001
R29686 D.n2402 D.n2393 0.001
R29687 D.n2388 D.n2379 0.001
R29688 D.n2374 D.n2365 0.001
R29689 D.n2360 D.n2351 0.001
R29690 D.n2875 D.n2864 0.001
R29691 D.n2889 D.n2880 0.001
R29692 D.n3365 D.n3356 0.001
R29693 D.n3351 D.n3342 0.001
R29694 D.n3337 D.n3328 0.001
R29695 D.n3323 D.n3314 0.001
R29696 D.n3309 D.n3300 0.001
R29697 D.n3295 D.n3286 0.001
R29698 D.n3281 D.n3272 0.001
R29699 D.n3267 D.n3258 0.001
R29700 D.n3253 D.n3244 0.001
R29701 D.n3239 D.n3230 0.001
R29702 D.n3225 D.n3216 0.001
R29703 D.n3211 D.n3202 0.001
R29704 D.n3197 D.n3188 0.001
R29705 D.n3183 D.n3174 0.001
R29706 D.n3169 D.n3160 0.001
R29707 D.n3155 D.n3146 0.001
R29708 D.n3141 D.n3132 0.001
R29709 D.n3127 D.n3118 0.001
R29710 D.n3113 D.n3104 0.001
R29711 D.n3099 D.n3090 0.001
R29712 D.n3085 D.n3076 0.001
R29713 D.n3071 D.n3062 0.001
R29714 D.n3057 D.n3048 0.001
R29715 D.n3043 D.n3034 0.001
R29716 D.n3029 D.n3020 0.001
R29717 D.n3015 D.n3006 0.001
R29718 D.n3001 D.n2992 0.001
R29719 D.n2987 D.n2978 0.001
R29720 D.n2973 D.n2964 0.001
R29721 D.n2959 D.n2950 0.001
R29722 D.n2945 D.n2936 0.001
R29723 D.n2931 D.n2922 0.001
R29724 D.n2917 D.n2908 0.001
R29725 D.n2903 D.n2894 0.001
R29726 D.n3391 D.n3380 0.001
R29727 D.n3405 D.n3396 0.001
R29728 D.n3853 D.n3844 0.001
R29729 D.n3839 D.n3830 0.001
R29730 D.n3825 D.n3816 0.001
R29731 D.n3811 D.n3802 0.001
R29732 D.n3797 D.n3788 0.001
R29733 D.n3783 D.n3774 0.001
R29734 D.n3769 D.n3760 0.001
R29735 D.n3755 D.n3746 0.001
R29736 D.n3741 D.n3732 0.001
R29737 D.n3727 D.n3718 0.001
R29738 D.n3713 D.n3704 0.001
R29739 D.n3699 D.n3690 0.001
R29740 D.n3685 D.n3676 0.001
R29741 D.n3671 D.n3662 0.001
R29742 D.n3657 D.n3648 0.001
R29743 D.n3643 D.n3634 0.001
R29744 D.n3629 D.n3620 0.001
R29745 D.n3615 D.n3606 0.001
R29746 D.n3601 D.n3592 0.001
R29747 D.n3587 D.n3578 0.001
R29748 D.n3573 D.n3564 0.001
R29749 D.n3559 D.n3550 0.001
R29750 D.n3545 D.n3536 0.001
R29751 D.n3531 D.n3522 0.001
R29752 D.n3517 D.n3508 0.001
R29753 D.n3503 D.n3494 0.001
R29754 D.n3489 D.n3480 0.001
R29755 D.n3475 D.n3466 0.001
R29756 D.n3461 D.n3452 0.001
R29757 D.n3447 D.n3438 0.001
R29758 D.n3433 D.n3424 0.001
R29759 D.n3419 D.n3410 0.001
R29760 D.n3879 D.n3868 0.001
R29761 D.n3893 D.n3884 0.001
R29762 D.n4313 D.n4304 0.001
R29763 D.n4299 D.n4290 0.001
R29764 D.n4285 D.n4276 0.001
R29765 D.n4271 D.n4262 0.001
R29766 D.n4257 D.n4248 0.001
R29767 D.n4243 D.n4234 0.001
R29768 D.n4229 D.n4220 0.001
R29769 D.n4215 D.n4206 0.001
R29770 D.n4201 D.n4192 0.001
R29771 D.n4187 D.n4178 0.001
R29772 D.n4173 D.n4164 0.001
R29773 D.n4159 D.n4150 0.001
R29774 D.n4145 D.n4136 0.001
R29775 D.n4131 D.n4122 0.001
R29776 D.n4117 D.n4108 0.001
R29777 D.n4103 D.n4094 0.001
R29778 D.n4089 D.n4080 0.001
R29779 D.n4075 D.n4066 0.001
R29780 D.n4061 D.n4052 0.001
R29781 D.n4047 D.n4038 0.001
R29782 D.n4033 D.n4024 0.001
R29783 D.n4019 D.n4010 0.001
R29784 D.n4005 D.n3996 0.001
R29785 D.n3991 D.n3982 0.001
R29786 D.n3977 D.n3968 0.001
R29787 D.n3963 D.n3954 0.001
R29788 D.n3949 D.n3940 0.001
R29789 D.n3935 D.n3926 0.001
R29790 D.n3921 D.n3912 0.001
R29791 D.n3907 D.n3898 0.001
R29792 D.n4339 D.n4328 0.001
R29793 D.n4353 D.n4344 0.001
R29794 D.n4745 D.n4736 0.001
R29795 D.n4731 D.n4722 0.001
R29796 D.n4717 D.n4708 0.001
R29797 D.n4703 D.n4694 0.001
R29798 D.n4689 D.n4680 0.001
R29799 D.n4675 D.n4666 0.001
R29800 D.n4661 D.n4652 0.001
R29801 D.n4647 D.n4638 0.001
R29802 D.n4633 D.n4624 0.001
R29803 D.n4619 D.n4610 0.001
R29804 D.n4605 D.n4596 0.001
R29805 D.n4591 D.n4582 0.001
R29806 D.n4577 D.n4568 0.001
R29807 D.n4563 D.n4554 0.001
R29808 D.n4549 D.n4540 0.001
R29809 D.n4535 D.n4526 0.001
R29810 D.n4521 D.n4512 0.001
R29811 D.n4507 D.n4498 0.001
R29812 D.n4493 D.n4484 0.001
R29813 D.n4479 D.n4470 0.001
R29814 D.n4465 D.n4456 0.001
R29815 D.n4451 D.n4442 0.001
R29816 D.n4437 D.n4428 0.001
R29817 D.n4423 D.n4414 0.001
R29818 D.n4409 D.n4400 0.001
R29819 D.n4395 D.n4386 0.001
R29820 D.n4381 D.n4372 0.001
R29821 D.n4367 D.n4358 0.001
R29822 D.n4771 D.n4760 0.001
R29823 D.n4785 D.n4776 0.001
R29824 D.n5149 D.n5140 0.001
R29825 D.n5135 D.n5126 0.001
R29826 D.n5121 D.n5112 0.001
R29827 D.n5107 D.n5098 0.001
R29828 D.n5093 D.n5084 0.001
R29829 D.n5079 D.n5070 0.001
R29830 D.n5065 D.n5056 0.001
R29831 D.n5051 D.n5042 0.001
R29832 D.n5037 D.n5028 0.001
R29833 D.n5023 D.n5014 0.001
R29834 D.n5009 D.n5000 0.001
R29835 D.n4995 D.n4986 0.001
R29836 D.n4981 D.n4972 0.001
R29837 D.n4967 D.n4958 0.001
R29838 D.n4953 D.n4944 0.001
R29839 D.n4939 D.n4930 0.001
R29840 D.n4925 D.n4916 0.001
R29841 D.n4911 D.n4902 0.001
R29842 D.n4897 D.n4888 0.001
R29843 D.n4883 D.n4874 0.001
R29844 D.n4869 D.n4860 0.001
R29845 D.n4855 D.n4846 0.001
R29846 D.n4841 D.n4832 0.001
R29847 D.n4827 D.n4818 0.001
R29848 D.n4813 D.n4804 0.001
R29849 D.n4799 D.n4790 0.001
R29850 D.n5175 D.n5164 0.001
R29851 D.n5189 D.n5180 0.001
R29852 D.n5525 D.n5516 0.001
R29853 D.n5511 D.n5502 0.001
R29854 D.n5497 D.n5488 0.001
R29855 D.n5483 D.n5474 0.001
R29856 D.n5469 D.n5460 0.001
R29857 D.n5455 D.n5446 0.001
R29858 D.n5441 D.n5432 0.001
R29859 D.n5427 D.n5418 0.001
R29860 D.n5413 D.n5404 0.001
R29861 D.n5399 D.n5390 0.001
R29862 D.n5385 D.n5376 0.001
R29863 D.n5371 D.n5362 0.001
R29864 D.n5357 D.n5348 0.001
R29865 D.n5343 D.n5334 0.001
R29866 D.n5329 D.n5320 0.001
R29867 D.n5315 D.n5306 0.001
R29868 D.n5301 D.n5292 0.001
R29869 D.n5287 D.n5278 0.001
R29870 D.n5273 D.n5264 0.001
R29871 D.n5259 D.n5250 0.001
R29872 D.n5245 D.n5236 0.001
R29873 D.n5231 D.n5222 0.001
R29874 D.n5217 D.n5208 0.001
R29875 D.n5203 D.n5194 0.001
R29876 D.n5551 D.n5540 0.001
R29877 D.n5565 D.n5556 0.001
R29878 D.n5873 D.n5864 0.001
R29879 D.n5859 D.n5850 0.001
R29880 D.n5845 D.n5836 0.001
R29881 D.n5831 D.n5822 0.001
R29882 D.n5817 D.n5808 0.001
R29883 D.n5803 D.n5794 0.001
R29884 D.n5789 D.n5780 0.001
R29885 D.n5775 D.n5766 0.001
R29886 D.n5761 D.n5752 0.001
R29887 D.n5747 D.n5738 0.001
R29888 D.n5733 D.n5724 0.001
R29889 D.n5719 D.n5710 0.001
R29890 D.n5705 D.n5696 0.001
R29891 D.n5691 D.n5682 0.001
R29892 D.n5677 D.n5668 0.001
R29893 D.n5663 D.n5654 0.001
R29894 D.n5649 D.n5640 0.001
R29895 D.n5635 D.n5626 0.001
R29896 D.n5621 D.n5612 0.001
R29897 D.n5607 D.n5598 0.001
R29898 D.n5593 D.n5584 0.001
R29899 D.n5579 D.n5570 0.001
R29900 D.n5899 D.n5888 0.001
R29901 D.n5913 D.n5904 0.001
R29902 D.n6193 D.n6184 0.001
R29903 D.n6179 D.n6170 0.001
R29904 D.n6165 D.n6156 0.001
R29905 D.n6151 D.n6142 0.001
R29906 D.n6137 D.n6128 0.001
R29907 D.n6123 D.n6114 0.001
R29908 D.n6109 D.n6100 0.001
R29909 D.n6095 D.n6086 0.001
R29910 D.n6081 D.n6072 0.001
R29911 D.n6067 D.n6058 0.001
R29912 D.n6053 D.n6044 0.001
R29913 D.n6039 D.n6030 0.001
R29914 D.n6025 D.n6016 0.001
R29915 D.n6011 D.n6002 0.001
R29916 D.n5997 D.n5988 0.001
R29917 D.n5983 D.n5974 0.001
R29918 D.n5969 D.n5960 0.001
R29919 D.n5955 D.n5946 0.001
R29920 D.n5941 D.n5932 0.001
R29921 D.n5927 D.n5918 0.001
R29922 D.n6219 D.n6208 0.001
R29923 D.n6233 D.n6224 0.001
R29924 D.n6485 D.n6476 0.001
R29925 D.n6471 D.n6462 0.001
R29926 D.n6457 D.n6448 0.001
R29927 D.n6443 D.n6434 0.001
R29928 D.n6429 D.n6420 0.001
R29929 D.n6415 D.n6406 0.001
R29930 D.n6401 D.n6392 0.001
R29931 D.n6387 D.n6378 0.001
R29932 D.n6373 D.n6364 0.001
R29933 D.n6359 D.n6350 0.001
R29934 D.n6345 D.n6336 0.001
R29935 D.n6331 D.n6322 0.001
R29936 D.n6317 D.n6308 0.001
R29937 D.n6303 D.n6294 0.001
R29938 D.n6289 D.n6280 0.001
R29939 D.n6275 D.n6266 0.001
R29940 D.n6261 D.n6252 0.001
R29941 D.n6247 D.n6238 0.001
R29942 D.n6511 D.n6500 0.001
R29943 D.n6525 D.n6516 0.001
R29944 D.n6749 D.n6740 0.001
R29945 D.n6735 D.n6726 0.001
R29946 D.n6721 D.n6712 0.001
R29947 D.n6707 D.n6698 0.001
R29948 D.n6693 D.n6684 0.001
R29949 D.n6679 D.n6670 0.001
R29950 D.n6665 D.n6656 0.001
R29951 D.n6651 D.n6642 0.001
R29952 D.n6637 D.n6628 0.001
R29953 D.n6623 D.n6614 0.001
R29954 D.n6609 D.n6600 0.001
R29955 D.n6595 D.n6586 0.001
R29956 D.n6581 D.n6572 0.001
R29957 D.n6567 D.n6558 0.001
R29958 D.n6553 D.n6544 0.001
R29959 D.n6539 D.n6530 0.001
R29960 D.n6775 D.n6764 0.001
R29961 D.n6789 D.n6780 0.001
R29962 D.n6985 D.n6976 0.001
R29963 D.n6971 D.n6962 0.001
R29964 D.n6957 D.n6948 0.001
R29965 D.n6943 D.n6934 0.001
R29966 D.n6929 D.n6920 0.001
R29967 D.n6915 D.n6906 0.001
R29968 D.n6901 D.n6892 0.001
R29969 D.n6887 D.n6878 0.001
R29970 D.n6873 D.n6864 0.001
R29971 D.n6859 D.n6850 0.001
R29972 D.n6845 D.n6836 0.001
R29973 D.n6831 D.n6822 0.001
R29974 D.n6817 D.n6808 0.001
R29975 D.n6803 D.n6794 0.001
R29976 D.n7011 D.n7000 0.001
R29977 D.n7025 D.n7016 0.001
R29978 D.n7193 D.n7184 0.001
R29979 D.n7179 D.n7170 0.001
R29980 D.n7165 D.n7156 0.001
R29981 D.n7151 D.n7142 0.001
R29982 D.n7137 D.n7128 0.001
R29983 D.n7123 D.n7114 0.001
R29984 D.n7109 D.n7100 0.001
R29985 D.n7095 D.n7086 0.001
R29986 D.n7081 D.n7072 0.001
R29987 D.n7067 D.n7058 0.001
R29988 D.n7053 D.n7044 0.001
R29989 D.n7039 D.n7030 0.001
R29990 D.n7219 D.n7208 0.001
R29991 D.n7233 D.n7224 0.001
R29992 D.n7373 D.n7364 0.001
R29993 D.n7359 D.n7350 0.001
R29994 D.n7345 D.n7336 0.001
R29995 D.n7331 D.n7322 0.001
R29996 D.n7317 D.n7308 0.001
R29997 D.n7303 D.n7294 0.001
R29998 D.n7289 D.n7280 0.001
R29999 D.n7275 D.n7266 0.001
R30000 D.n7261 D.n7252 0.001
R30001 D.n7247 D.n7238 0.001
R30002 D.n7399 D.n7388 0.001
R30003 D.n7413 D.n7404 0.001
R30004 D.n7525 D.n7516 0.001
R30005 D.n7511 D.n7502 0.001
R30006 D.n7497 D.n7488 0.001
R30007 D.n7483 D.n7474 0.001
R30008 D.n7469 D.n7460 0.001
R30009 D.n7455 D.n7446 0.001
R30010 D.n7441 D.n7432 0.001
R30011 D.n7427 D.n7418 0.001
R30012 D.n7551 D.n7540 0.001
R30013 D.n7565 D.n7556 0.001
R30014 D.n7649 D.n7640 0.001
R30015 D.n7635 D.n7626 0.001
R30016 D.n7621 D.n7612 0.001
R30017 D.n7607 D.n7598 0.001
R30018 D.n7593 D.n7584 0.001
R30019 D.n7579 D.n7570 0.001
R30020 D.n7675 D.n7664 0.001
R30021 D.n7689 D.n7680 0.001
R30022 D.n7745 D.n7736 0.001
R30023 D.n7731 D.n7722 0.001
R30024 D.n7717 D.n7708 0.001
R30025 D.n7703 D.n7694 0.001
R30026 D.n7770 D.n7759 0.001
R30027 D.n7784 D.n7775 0.001
R30028 D.n7814 D.n7803 0.001
R30029 D.n7798 D.n7789 0.001
R30030 D.n7902 D.n7893 0.001
R30031 D.n7988 D.n7977 0.001
R30032 D.n13679 D.n13660 0.001
R30033 D.n13636 D.n13625 0.001
R30034 D.n12752 D.n12737 0.001
R30035 D.n12713 D.n12702 0.001
R30036 D.n11903 D.n11888 0.001
R30037 D.n11864 D.n11853 0.001
R30038 D.n11140 D.n11125 0.001
R30039 D.n11101 D.n11090 0.001
R30040 D.n10457 D.n10442 0.001
R30041 D.n10418 D.n10407 0.001
R30042 D.n9854 D.n9839 0.001
R30043 D.n9815 D.n9804 0.001
R30044 D.n9325 D.n9310 0.001
R30045 D.n9286 D.n9275 0.001
R30046 D.n8882 D.n8867 0.001
R30047 D.n8843 D.n8832 0.001
R30048 D.n8519 D.n8504 0.001
R30049 D.n8480 D.n8469 0.001
R30050 D.n8230 D.n8215 0.001
R30051 D.n8191 D.n8180 0.001
R30052 D.n8027 D.n8012 0.001
R30053 D.n455 D.n454 0.001
R30054 D.n7823 D.n7821 0.001
R30055 D.n533 D.n531 0.001
R30056 D.n1160 D.n1158 0.001
R30057 D.n1759 D.n1757 0.001
R30058 D.n2330 D.n2328 0.001
R30059 D.n2873 D.n2871 0.001
R30060 D.n3389 D.n3387 0.001
R30061 D.n3877 D.n3875 0.001
R30062 D.n4337 D.n4335 0.001
R30063 D.n4769 D.n4767 0.001
R30064 D.n5173 D.n5171 0.001
R30065 D.n5549 D.n5547 0.001
R30066 D.n5897 D.n5895 0.001
R30067 D.n6217 D.n6215 0.001
R30068 D.n6509 D.n6507 0.001
R30069 D.n6773 D.n6771 0.001
R30070 D.n7009 D.n7007 0.001
R30071 D.n7217 D.n7215 0.001
R30072 D.n7397 D.n7395 0.001
R30073 D.n7549 D.n7547 0.001
R30074 D.n7673 D.n7671 0.001
R30075 D.n7768 D.n7766 0.001
R30076 D.n7860 D.n7858 0.001
R30077 D.n7861 D.n7856 0.001
R30078 S.n22291 S.n22290 153.554
R30079 S.n18062 S.n18061 153.554
R30080 S.n18946 S.n18945 153.554
R30081 S.n19817 S.n19816 153.554
R30082 S.n20454 S.n20453 153.554
R30083 S.n21299 S.n21298 153.554
R30084 S.n16235 S.n16234 153.554
R30085 S.n17154 S.n17153 153.554
R30086 S.n14338 S.n14337 153.554
R30087 S.n15292 S.n15291 153.554
R30088 S.n12371 S.n12370 153.554
R30089 S.n13360 S.n13359 153.554
R30090 S.n10334 S.n10333 153.554
R30091 S.n11358 S.n11357 153.554
R30092 S.n8227 S.n8226 153.554
R30093 S.n9286 S.n9285 153.554
R30094 S.n6050 S.n6049 153.554
R30095 S.n7144 S.n7143 153.554
R30096 S.n3802 S.n3801 153.554
R30097 S.n4931 S.n4930 153.554
R30098 S.n1463 S.n1462 153.554
R30099 S.n2656 S.n2655 153.554
R30100 S.n435 S.n434 153.554
R30101 S.n20338 S.n20337 153.118
R30102 S.n21141 S.n21140 153.118
R30103 S.n19498 S.n19497 153.118
R30104 S.n18641 S.n18640 153.118
R30105 S.n17773 S.n17772 153.118
R30106 S.n16879 S.n16878 153.118
R30107 S.n15976 S.n15975 153.118
R30108 S.n15047 S.n15046 153.118
R30109 S.n14109 S.n14108 153.118
R30110 S.n13145 S.n13144 153.118
R30111 S.n12172 S.n12171 153.118
R30112 S.n11173 S.n11172 153.118
R30113 S.n10165 S.n10164 153.118
R30114 S.n9131 S.n9130 153.118
R30115 S.n8088 S.n8087 153.118
R30116 S.n7019 S.n7018 153.118
R30117 S.n5941 S.n5940 153.118
R30118 S.n4835 S.n4834 153.118
R30119 S.n3722 S.n3721 153.118
R30120 S.n2591 S.n2590 153.118
R30121 S.n22773 S.n22772 153.118
R30122 S.n976 S.n975 153.118
R30123 S.n21970 S.n21969 153.118
R30124 S.n1421 S.n1420 146.135
R30125 S.n1300 S.n1299 146.135
R30126 S.n1418 S.n1417 146.135
R30127 S.n1315 S.n1314 146.135
R30128 S.n1362 S.n1361 146.135
R30129 S.n1379 S.n1378 146.135
R30130 S.n1288 S.n1287 146.135
R30131 S.n1414 S.n1413 146.135
R30132 S.n1276 S.n1275 146.135
R30133 S.n1410 S.n1409 146.135
R30134 S.n1263 S.n1262 146.135
R30135 S.n1406 S.n1405 146.135
R30136 S.n1250 S.n1249 146.135
R30137 S.n1402 S.n1401 146.135
R30138 S.n1237 S.n1236 146.135
R30139 S.n1398 S.n1397 146.135
R30140 S.n1224 S.n1223 146.135
R30141 S.n1394 S.n1393 146.135
R30142 S.n1211 S.n1210 146.135
R30143 S.n1390 S.n1389 146.135
R30144 S.n1198 S.n1197 146.135
R30145 S.n1386 S.n1385 146.135
R30146 S.n1382 S.n1381 146.135
R30147 S.n22957 S.n22956 145.699
R30148 S.n22964 S.n22963 145.699
R30149 S.n22950 S.n22949 145.699
R30150 S.n22943 S.n22942 145.699
R30151 S.n22936 S.n22935 145.699
R30152 S.n22929 S.n22928 145.699
R30153 S.n22922 S.n22921 145.699
R30154 S.n22915 S.n22914 145.699
R30155 S.n22908 S.n22907 145.699
R30156 S.n22901 S.n22900 145.699
R30157 S.n22894 S.n22893 145.699
R30158 S.n22887 S.n22886 145.699
R30159 S.n22880 S.n22879 145.699
R30160 S.n22873 S.n22872 145.699
R30161 S.n22866 S.n22865 145.699
R30162 S.n22859 S.n22858 145.699
R30163 S.n22852 S.n22851 145.699
R30164 S.n22845 S.n22844 145.699
R30165 S.n22838 S.n22837 145.699
R30166 S.n22829 S.n22828 145.699
R30167 S.n22815 S.n22814 145.699
R30168 S.n22820 S.n22819 145.699
R30169 S.n22995 S.n22994 145.699
R30170 S.n422 S.n421 101.08
R30171 S.n1452 S.n1451 101.08
R30172 S.n2646 S.n2645 101.08
R30173 S.n3791 S.n3790 101.08
R30174 S.n4921 S.n4920 101.08
R30175 S.n6039 S.n6038 101.08
R30176 S.n7134 S.n7133 101.08
R30177 S.n8216 S.n8215 101.08
R30178 S.n9276 S.n9275 101.08
R30179 S.n10323 S.n10322 101.08
R30180 S.n11348 S.n11347 101.08
R30181 S.n12360 S.n12359 101.08
R30182 S.n13350 S.n13349 101.08
R30183 S.n14327 S.n14326 101.08
R30184 S.n15282 S.n15281 101.08
R30185 S.n16224 S.n16223 101.08
R30186 S.n17144 S.n17143 101.08
R30187 S.n18051 S.n18050 101.08
R30188 S.n18936 S.n18935 101.08
R30189 S.n19806 S.n19805 101.08
R30190 S.n20444 S.n20443 101.08
R30191 S.n21288 S.n21287 101.08
R30192 S.n22276 S.n22275 101.08
R30193 S.n961 S.n960 98.123
R30194 S.n22793 S.n22792 88.439
R30195 S.n424 S.n423 68.042
R30196 S.n2602 S.n2601 68.042
R30197 S.n3733 S.n3732 68.042
R30198 S.n4846 S.n4845 68.042
R30199 S.n5951 S.n5950 68.042
R30200 S.n7029 S.n7028 68.042
R30201 S.n8098 S.n8097 68.042
R30202 S.n9141 S.n9140 68.042
R30203 S.n10175 S.n10174 68.042
R30204 S.n11183 S.n11182 68.042
R30205 S.n12182 S.n12181 68.042
R30206 S.n13155 S.n13154 68.042
R30207 S.n14119 S.n14118 68.042
R30208 S.n15057 S.n15056 68.042
R30209 S.n15986 S.n15985 68.042
R30210 S.n16889 S.n16888 68.042
R30211 S.n17783 S.n17782 68.042
R30212 S.n18651 S.n18650 68.042
R30213 S.n19508 S.n19507 68.042
R30214 S.n21158 S.n21157 68.042
R30215 S.n21176 S.n21175 68.042
R30216 S.n22786 S.n22785 68.042
R30217 S.n22278 S.n22277 65.312
R30218 S.n22777 S.n22776 62.872
R30219 S.n21179 S.n21178 62.872
R30220 S.n21161 S.n21160 62.872
R30221 S.n19511 S.n19510 62.872
R30222 S.n18654 S.n18653 62.872
R30223 S.n17786 S.n17785 62.872
R30224 S.n16892 S.n16891 62.872
R30225 S.n15989 S.n15988 62.872
R30226 S.n15060 S.n15059 62.872
R30227 S.n14122 S.n14121 62.872
R30228 S.n13158 S.n13157 62.872
R30229 S.n12185 S.n12184 62.872
R30230 S.n11186 S.n11185 62.872
R30231 S.n10178 S.n10177 62.872
R30232 S.n9144 S.n9143 62.872
R30233 S.n8101 S.n8100 62.872
R30234 S.n7032 S.n7031 62.872
R30235 S.n5954 S.n5953 62.872
R30236 S.n4849 S.n4848 62.872
R30237 S.n3736 S.n3735 62.872
R30238 S.n2605 S.n2604 62.872
R30239 S.n1905 S.n1904 62.872
R30240 S.n964 S.n963 62.872
R30241 S.n22794 S.n22793 10.138
R30242 S.t158 S.t51 9.465
R30243 S.n969 S.t95 8.26
R30244 S.n425 S.t122 8.26
R30245 S.n1909 S.t128 8.26
R30246 S.n1453 S.t143 8.26
R30247 S.n2610 S.t193 8.26
R30248 S.n2647 S.t33 8.26
R30249 S.n3741 S.t116 8.26
R30250 S.n3792 S.t81 8.26
R30251 S.n4854 S.t118 8.26
R30252 S.n4922 S.t11 8.26
R30253 S.n5959 S.t35 8.26
R30254 S.n6040 S.t332 8.26
R30255 S.n7037 S.t152 8.26
R30256 S.n7135 S.t23 8.26
R30257 S.n8106 S.t4 8.26
R30258 S.n8217 S.t216 8.26
R30259 S.n9149 S.t58 8.26
R30260 S.n9277 S.t198 8.26
R30261 S.n10183 S.t45 8.26
R30262 S.n10324 S.t56 8.26
R30263 S.n11191 S.t16 8.26
R30264 S.n11349 S.t25 8.26
R30265 S.n12190 S.t37 8.26
R30266 S.n12361 S.t221 8.26
R30267 S.n13163 S.t43 8.26
R30268 S.n13351 S.t97 8.26
R30269 S.n14127 S.t2 8.26
R30270 S.n14328 S.t139 8.26
R30271 S.n15065 S.t330 8.26
R30272 S.n15283 S.t165 8.26
R30273 S.n15994 S.t231 8.26
R30274 S.n16225 S.t49 8.26
R30275 S.n16897 S.t148 8.26
R30276 S.n17145 S.t126 8.26
R30277 S.n17791 S.t321 8.26
R30278 S.n18052 S.t183 8.26
R30279 S.n18659 S.t174 8.26
R30280 S.n18937 S.t39 8.26
R30281 S.n19516 S.t388 8.26
R30282 S.n19807 S.t114 8.26
R30283 S.n21166 S.t91 8.26
R30284 S.n20445 S.t181 8.26
R30285 S.n21184 S.t200 8.26
R30286 S.n21289 S.t27 8.26
R30287 S.n22782 S.t62 8.26
R30288 S.n22280 S.t70 8.26
R30289 S.t109 S.n921 7.985
R30290 S.t137 S.n793 7.985
R30291 S.t270 S.n1961 7.985
R30292 S.t75 S.n1872 7.985
R30293 S.t163 S.n3121 7.985
R30294 S.t14 S.n3032 7.985
R30295 S.t134 S.n4257 7.985
R30296 S.t176 S.n4158 7.985
R30297 S.t288 S.n5391 7.985
R30298 S.t214 S.n5271 7.985
R30299 S.t130 S.n6502 7.985
R30300 S.t83 S.n6371 7.985
R30301 S.t406 S.n7600 7.985
R30302 S.t47 S.n7448 7.985
R30303 S.t141 S.n8675 7.985
R30304 S.t19 S.n8512 7.985
R30305 S.t160 S.n9738 7.985
R30306 S.t366 S.n9554 7.985
R30307 S.t172 S.n10778 7.985
R30308 S.t31 S.n10583 7.985
R30309 S.t67 S.n11806 7.985
R30310 S.t54 S.n11590 7.985
R30311 S.t443 S.n12811 7.985
R30312 S.t357 S.n12584 7.985
R30313 S.t538 S.n13804 7.985
R30314 S.t73 S.n13556 7.985
R30315 S.t102 S.n14774 7.985
R30316 S.t0 S.n14515 7.985
R30317 S.t29 S.n15732 7.985
R30318 S.t60 S.n15452 7.985
R30319 S.t187 S.n16667 7.985
R30320 S.t167 S.n16376 7.985
R30321 S.t169 S.n17590 7.985
R30322 S.t218 S.n17278 7.985
R30323 S.t77 S.n18490 7.985
R30324 S.t79 S.n18167 7.985
R30325 S.t21 S.n19377 7.985
R30326 S.t150 S.n19033 7.985
R30327 S.t262 S.n20245 7.985
R30328 S.t209 S.n19887 7.985
R30329 S.t7 S.n20405 7.985
R30330 S.t64 S.n20498 7.985
R30331 S.t105 S.n21224 7.985
R30332 S.t100 S.n21335 7.985
R30333 S.t88 S.n22748 7.985
R30334 S.t9 S.n22340 7.985
R30335 S.t41 S.n22817 7.985
R30336 S.n22997 S.t2791 6.541
R30337 S.n22805 S.t1797 6.541
R30338 S.n20338 S.t263 6.541
R30339 S.n20177 S.n20176 6.541
R30340 S.n20185 S.t3797 6.541
R30341 S.n20188 S.t1924 6.541
R30342 S.n20180 S.n20179 6.541
R30343 S.n21131 S.n21130 6.541
R30344 S.n21135 S.t2724 6.541
R30345 S.n21138 S.t384 6.541
R30346 S.n21128 S.n21127 6.541
R30347 S.n22957 S.t269 6.541
R30348 S.n22955 S.t4049 6.541
R30349 S.n22637 S.n22636 6.541
R30350 S.n22642 S.t4285 6.541
R30351 S.n22645 S.t3260 6.541
R30352 S.n22634 S.n22633 6.541
R30353 S.n22008 S.n22007 6.541
R30354 S.n22015 S.t1155 6.541
R30355 S.n22012 S.t1991 6.541
R30356 S.n22005 S.n22004 6.541
R30357 S.n21614 S.n21613 6.541
R30358 S.n21619 S.t4391 6.541
R30359 S.n21622 S.t339 6.541
R30360 S.n21611 S.n21610 6.541
R30361 S.n21940 S.n21939 6.541
R30362 S.n21944 S.t2773 6.541
R30363 S.n21947 S.t1944 6.541
R30364 S.n21937 S.n21936 6.541
R30365 S.n20791 S.n20790 6.541
R30366 S.n20796 S.t4336 6.541
R30367 S.n20799 S.t295 6.541
R30368 S.n20788 S.n20787 6.541
R30369 S.n21141 S.t2349 6.541
R30370 S.n21143 S.t3564 6.541
R30371 S.n22964 S.t3247 6.541
R30372 S.n22962 S.t2508 6.541
R30373 S.n22650 S.n22649 6.541
R30374 S.n22658 S.t2728 6.541
R30375 S.n22661 S.t1705 6.541
R30376 S.n22653 S.n22652 6.541
R30377 S.n21989 S.n21988 6.541
R30378 S.n22000 S.t4108 6.541
R30379 S.n21997 S.t435 6.541
R30380 S.n21992 S.n21991 6.541
R30381 S.n21632 S.n21631 6.541
R30382 S.n21640 S.t2836 6.541
R30383 S.n21643 S.t3306 6.541
R30384 S.n21635 S.n21634 6.541
R30385 S.n21955 S.n21954 6.541
R30386 S.n21964 S.t1213 6.541
R30387 S.n21967 S.t2446 6.541
R30388 S.n21958 S.n21957 6.541
R30389 S.n20809 S.n20808 6.541
R30390 S.n20820 S.t1324 6.541
R30391 S.n20823 S.t3916 6.541
R30392 S.n20812 S.n20811 6.541
R30393 S.n20342 S.t556 6.541
R30394 S.n19498 S.t3847 6.541
R30395 S.n19307 S.n19306 6.541
R30396 S.n19315 S.t1734 6.541
R30397 S.n19318 S.t4413 6.541
R30398 S.n19310 S.n19309 6.541
R30399 S.n19531 S.n19530 6.541
R30400 S.n19538 S.t4224 6.541
R30401 S.n19535 S.t2823 6.541
R30402 S.n19528 S.n19527 6.541
R30403 S.n22950 S.t1833 6.541
R30404 S.n22948 S.t1083 6.541
R30405 S.n22621 S.n22620 6.541
R30406 S.n22626 S.t1337 6.541
R30407 S.n22629 S.t285 6.541
R30408 S.n22618 S.n22617 6.541
R30409 S.n22023 S.n22022 6.541
R30410 S.n22030 S.t2716 6.541
R30411 S.n22027 S.t3540 6.541
R30412 S.n22020 S.n22019 6.541
R30413 S.n21598 S.n21597 6.541
R30414 S.n21603 S.t1442 6.541
R30415 S.n21606 S.t1896 6.541
R30416 S.n21595 S.n21594 6.541
R30417 S.n21925 S.n21924 6.541
R30418 S.n21929 S.t4328 6.541
R30419 S.n21932 S.t3490 6.541
R30420 S.n21922 S.n21921 6.541
R30421 S.n20775 S.n20774 6.541
R30422 S.n20780 S.t1385 6.541
R30423 S.n20783 S.t1855 6.541
R30424 S.n20772 S.n20771 6.541
R30425 S.n21115 S.n21114 6.541
R30426 S.n21119 S.t4278 6.541
R30427 S.n21122 S.t3448 6.541
R30428 S.n21112 S.n21111 6.541
R30429 S.n20164 S.n20163 6.541
R30430 S.n20169 S.t1334 6.541
R30431 S.n20172 S.t1811 6.541
R30432 S.n20161 S.n20160 6.541
R30433 S.n19502 S.t2071 6.541
R30434 S.n18641 S.t1786 6.541
R30435 S.n18425 S.n18424 6.541
R30436 S.n18433 S.t4131 6.541
R30437 S.n18436 S.t1212 6.541
R30438 S.n18428 S.n18427 6.541
R30439 S.n18674 S.n18673 6.541
R30440 S.n18681 S.t4204 6.541
R30441 S.n18678 S.t789 6.541
R30442 S.n18671 S.n18670 6.541
R30443 S.n22943 S.t3168 6.541
R30444 S.n22941 S.t2642 6.541
R30445 S.n22605 S.n22604 6.541
R30446 S.n22610 S.t2647 6.541
R30447 S.n22613 S.t1846 6.541
R30448 S.n22602 S.n22601 6.541
R30449 S.n22038 S.n22037 6.541
R30450 S.n22045 S.t4268 6.541
R30451 S.n22042 S.t589 6.541
R30452 S.n22035 S.n22034 6.541
R30453 S.n21582 S.n21581 6.541
R30454 S.n21587 S.t3001 6.541
R30455 S.n21590 S.t3441 6.541
R30456 S.n21579 S.n21578 6.541
R30457 S.n21910 S.n21909 6.541
R30458 S.n21914 S.t1381 6.541
R30459 S.n21917 S.t534 6.541
R30460 S.n21907 S.n21906 6.541
R30461 S.n20759 S.n20758 6.541
R30462 S.n20764 S.t2950 6.541
R30463 S.n20767 S.t3398 6.541
R30464 S.n20756 S.n20755 6.541
R30465 S.n21100 S.n21099 6.541
R30466 S.n21104 S.t1327 6.541
R30467 S.n21107 S.t487 6.541
R30468 S.n21097 S.n21096 6.541
R30469 S.n20148 S.n20147 6.541
R30470 S.n20153 S.t2899 6.541
R30471 S.n20156 S.t3356 6.541
R30472 S.n20145 S.n20144 6.541
R30473 S.n19546 S.n19545 6.541
R30474 S.n19553 S.t1273 6.541
R30475 S.n19550 S.t447 6.541
R30476 S.n19543 S.n19542 6.541
R30477 S.n19294 S.n19293 6.541
R30478 S.n19299 S.t2847 6.541
R30479 S.n19302 S.t3315 6.541
R30480 S.n19291 S.n19290 6.541
R30481 S.n18645 S.t3572 6.541
R30482 S.n17773 S.t4189 6.541
R30483 S.n17520 S.n17519 6.541
R30484 S.n17528 S.t2116 6.541
R30485 S.n17531 S.t3764 6.541
R30486 S.n17523 S.n17522 6.541
R30487 S.n17806 S.n17805 6.541
R30488 S.n17813 S.t1197 6.541
R30489 S.n17810 S.t3234 6.541
R30490 S.n17803 S.n17802 6.541
R30491 S.n22936 S.t185 6.541
R30492 S.n22934 S.t4191 6.541
R30493 S.n22589 S.n22588 6.541
R30494 S.n22594 S.t4196 6.541
R30495 S.n22597 S.t3389 6.541
R30496 S.n22586 S.n22585 6.541
R30497 S.n22053 S.n22052 6.541
R30498 S.n22060 S.t1317 6.541
R30499 S.n22057 S.t1917 6.541
R30500 S.n22050 S.n22049 6.541
R30501 S.n21566 S.n21565 6.541
R30502 S.n21571 S.t4298 6.541
R30503 S.n21574 S.t480 6.541
R30504 S.n21563 S.n21562 6.541
R30505 S.n21895 S.n21894 6.541
R30506 S.n21899 S.t2945 6.541
R30507 S.n21902 S.t2103 6.541
R30508 S.n21892 S.n21891 6.541
R30509 S.n20743 S.n20742 6.541
R30510 S.n20748 S.t4506 6.541
R30511 S.n20751 S.t440 6.541
R30512 S.n20740 S.n20739 6.541
R30513 S.n21085 S.n21084 6.541
R30514 S.n21089 S.t2893 6.541
R30515 S.n21092 S.t2051 6.541
R30516 S.n21082 S.n21081 6.541
R30517 S.n20132 S.n20131 6.541
R30518 S.n20137 S.t4455 6.541
R30519 S.n20140 S.t389 6.541
R30520 S.n20129 S.n20128 6.541
R30521 S.n19561 S.n19560 6.541
R30522 S.n19568 S.t2841 6.541
R30523 S.n19565 S.t2001 6.541
R30524 S.n19558 S.n19557 6.541
R30525 S.n19278 S.n19277 6.541
R30526 S.n19283 S.t4399 6.541
R30527 S.n19286 S.t347 6.541
R30528 S.n19275 S.n19274 6.541
R30529 S.n18689 S.n18688 6.541
R30530 S.n18696 S.t1249 6.541
R30531 S.n18693 S.t1956 6.541
R30532 S.n18686 S.n18685 6.541
R30533 S.n18412 S.n18411 6.541
R30534 S.n18417 S.t4345 6.541
R30535 S.n18420 S.t3292 6.541
R30536 S.n18409 S.n18408 6.541
R30537 S.n17777 S.t567 6.541
R30538 S.n16879 S.t2180 6.541
R30539 S.n16602 S.n16601 6.541
R30540 S.n16610 S.t4563 6.541
R30541 S.n16613 S.t1753 6.541
R30542 S.n16605 S.n16604 6.541
R30543 S.n16912 S.n16911 6.541
R30544 S.n16919 S.t2707 6.541
R30545 S.n16916 S.t1116 6.541
R30546 S.n16909 S.n16908 6.541
R30547 S.n22929 S.t1754 6.541
R30548 S.n22927 S.t1236 6.541
R30549 S.n22573 S.n22572 6.541
R30550 S.n22578 S.t1243 6.541
R30551 S.n22581 S.t428 6.541
R30552 S.n22570 S.n22569 6.541
R30553 S.n22068 S.n22067 6.541
R30554 S.n22075 S.t2885 6.541
R30555 S.n22072 S.t3463 6.541
R30556 S.n22065 S.n22064 6.541
R30557 S.n21550 S.n21549 6.541
R30558 S.n21555 S.t1349 6.541
R30559 S.n21558 S.t2043 6.541
R30560 S.n21547 S.n21546 6.541
R30561 S.n21880 S.n21879 6.541
R30562 S.n21884 S.t4501 6.541
R30563 S.n21887 S.t3418 6.541
R30564 S.n21877 S.n21876 6.541
R30565 S.n20727 S.n20726 6.541
R30566 S.n20732 S.t1292 6.541
R30567 S.n20735 S.t1997 6.541
R30568 S.n20724 S.n20723 6.541
R30569 S.n21070 S.n21069 6.541
R30570 S.n21074 S.t4448 6.541
R30571 S.n21077 S.t3607 6.541
R30572 S.n21067 S.n21066 6.541
R30573 S.n20116 S.n20115 6.541
R30574 S.n20121 S.t1508 6.541
R30575 S.n20124 S.t1948 6.541
R30576 S.n20113 S.n20112 6.541
R30577 S.n19576 S.n19575 6.541
R30578 S.n19583 S.t4396 6.541
R30579 S.n19580 S.t3551 6.541
R30580 S.n19573 S.n19572 6.541
R30581 S.n19262 S.n19261 6.541
R30582 S.n19267 S.t1451 6.541
R30583 S.n19270 S.t1906 6.541
R30584 S.n19259 S.n19258 6.541
R30585 S.n18704 S.n18703 6.541
R30586 S.n18711 S.t2812 6.541
R30587 S.n18708 S.t3500 6.541
R30588 S.n18701 S.n18700 6.541
R30589 S.n18396 S.n18395 6.541
R30590 S.n18401 S.t1395 6.541
R30591 S.n18404 S.t322 6.541
R30592 S.n18393 S.n18392 6.541
R30593 S.n17821 S.n17820 6.541
R30594 S.n17828 S.t2756 6.541
R30595 S.n17825 S.t3455 6.541
R30596 S.n17818 S.n17817 6.541
R30597 S.n17507 S.n17506 6.541
R30598 S.n17512 S.t1345 6.541
R30599 S.n17515 S.t282 6.541
R30600 S.n17504 S.n17503 6.541
R30601 S.n16883 S.t2084 6.541
R30602 S.n15976 S.t30 6.541
R30603 S.n15662 S.n15661 6.541
R30604 S.n15670 S.t2472 6.541
R30605 S.n15673 S.t4210 6.541
R30606 S.n15665 S.n15664 6.541
R30607 S.n16009 S.n16008 6.541
R30608 S.n16016 S.t4211 6.541
R30609 S.n16013 S.t3609 6.541
R30610 S.n16006 S.n16005 6.541
R30611 S.n22922 S.t3302 6.541
R30612 S.n22920 S.t2799 6.541
R30613 S.n22557 S.n22556 6.541
R30614 S.n22562 S.t2808 6.541
R30615 S.n22565 S.t1987 6.541
R30616 S.n22554 S.n22553 6.541
R30617 S.n22083 S.n22082 6.541
R30618 S.n22090 S.t4444 6.541
R30619 S.n22087 S.t503 6.541
R30620 S.n22080 S.n22079 6.541
R30621 S.n21534 S.n21533 6.541
R30622 S.n21539 S.t2914 6.541
R30623 S.n21542 S.t3598 6.541
R30624 S.n21531 S.n21530 6.541
R30625 S.n21865 S.n21864 6.541
R30626 S.n21869 S.t1556 6.541
R30627 S.n21872 S.t459 6.541
R30628 S.n21862 S.n21861 6.541
R30629 S.n20711 S.n20710 6.541
R30630 S.n20716 S.t2860 6.541
R30631 S.n20719 S.t3546 6.541
R30632 S.n20708 S.n20707 6.541
R30633 S.n21055 S.n21054 6.541
R30634 S.n21059 S.t1501 6.541
R30635 S.n21062 S.t412 6.541
R30636 S.n21052 S.n21051 6.541
R30637 S.n20100 S.n20099 6.541
R30638 S.n20105 S.t2802 6.541
R30639 S.n20108 S.t3495 6.541
R30640 S.n20097 S.n20096 6.541
R30641 S.n19591 S.n19590 6.541
R30642 S.n19598 S.t1445 6.541
R30643 S.n19595 S.t597 6.541
R30644 S.n19588 S.n19587 6.541
R30645 S.n19246 S.n19245 6.541
R30646 S.n19251 S.t3012 6.541
R30647 S.n19254 S.t3450 6.541
R30648 S.n19243 S.n19242 6.541
R30649 S.n18719 S.n18718 6.541
R30650 S.n18726 S.t4365 6.541
R30651 S.n18723 S.t544 6.541
R30652 S.n18716 S.n18715 6.541
R30653 S.n18380 S.n18379 6.541
R30654 S.n18385 S.t2963 6.541
R30655 S.n18388 S.t1882 6.541
R30656 S.n18377 S.n18376 6.541
R30657 S.n17836 S.n17835 6.541
R30658 S.n17843 S.t4312 6.541
R30659 S.n17840 S.t495 6.541
R30660 S.n17833 S.n17832 6.541
R30661 S.n17491 S.n17490 6.541
R30662 S.n17496 S.t2909 6.541
R30663 S.n17499 S.t1845 6.541
R30664 S.n17488 S.n17487 6.541
R30665 S.n16927 S.n16926 6.541
R30666 S.n16934 S.t4261 6.541
R30667 S.n16931 S.t455 6.541
R30668 S.n16924 S.n16923 6.541
R30669 S.n16589 S.n16588 6.541
R30670 S.n16594 S.t2854 6.541
R30671 S.n16597 S.t1793 6.541
R30672 S.n16586 S.n16585 6.541
R30673 S.n15980 S.t3583 6.541
R30674 S.n15047 S.t2627 6.541
R30675 S.n14709 S.n14708 6.541
R30676 S.n14717 S.t418 6.541
R30677 S.n14720 S.t1862 6.541
R30678 S.n14712 S.n14711 6.541
R30679 S.n15080 S.n15079 6.541
R30680 S.n15087 S.t1208 6.541
R30681 S.n15084 S.t1552 6.541
R30682 S.n15077 S.n15076 6.541
R30683 S.n22915 S.t771 6.541
R30684 S.n22913 S.t1742 6.541
R30685 S.n22541 S.n22540 6.541
R30686 S.n22546 S.t4306 6.541
R30687 S.n22549 S.t3533 6.541
R30688 S.n22538 S.n22537 6.541
R30689 S.n22098 S.n22097 6.541
R30690 S.n22105 S.t1496 6.541
R30691 S.n22102 S.t2068 6.541
R30692 S.n22095 S.n22094 6.541
R30693 S.n21518 S.n21517 6.541
R30694 S.n21523 S.t4469 6.541
R30695 S.n21526 S.t645 6.541
R30696 S.n21515 S.n21514 6.541
R30697 S.n21850 S.n21849 6.541
R30698 S.n21854 S.t3108 6.541
R30699 S.n21857 S.t2019 6.541
R30700 S.n21847 S.n21846 6.541
R30701 S.n20695 S.n20694 6.541
R30702 S.n20700 S.t4412 6.541
R30703 S.n20703 S.t592 6.541
R30704 S.n20692 S.n20691 6.541
R30705 S.n21040 S.n21039 6.541
R30706 S.n21044 S.t3056 6.541
R30707 S.n21047 S.t1965 6.541
R30708 S.n21037 S.n21036 6.541
R30709 S.n20084 S.n20083 6.541
R30710 S.n20089 S.t4359 6.541
R30711 S.n20092 S.t540 6.541
R30712 S.n20081 S.n20080 6.541
R30713 S.n19606 S.n19605 6.541
R30714 S.n19613 S.t3008 6.541
R30715 S.n19610 S.t1923 6.541
R30716 S.n19603 S.n19602 6.541
R30717 S.n19230 S.n19229 6.541
R30718 S.n19235 S.t4302 6.541
R30719 S.n19238 S.t492 6.541
R30720 S.n19227 S.n19226 6.541
R30721 S.n18734 S.n18733 6.541
R30722 S.n18741 S.t1419 6.541
R30723 S.n18738 S.t2111 6.541
R30724 S.n18731 S.n18730 6.541
R30725 S.n18364 S.n18363 6.541
R30726 S.n18369 S.t4520 6.541
R30727 S.n18372 S.t3428 6.541
R30728 S.n18361 S.n18360 6.541
R30729 S.n17851 S.n17850 6.541
R30730 S.n17858 S.t1363 6.541
R30731 S.n17855 S.t2061 6.541
R30732 S.n17848 S.n17847 6.541
R30733 S.n17475 S.n17474 6.541
R30734 S.n17480 S.t4465 6.541
R30735 S.n17483 S.t3387 6.541
R30736 S.n17472 S.n17471 6.541
R30737 S.n16942 S.n16941 6.541
R30738 S.n16949 S.t1311 6.541
R30739 S.n16946 S.t2012 6.541
R30740 S.n16939 S.n16938 6.541
R30741 S.n16573 S.n16572 6.541
R30742 S.n16578 S.t4407 6.541
R30743 S.n16581 S.t3342 6.541
R30744 S.n16570 S.n16569 6.541
R30745 S.n16024 S.n16023 6.541
R30746 S.n16031 S.t1256 6.541
R30747 S.n16028 S.t1962 6.541
R30748 S.n16021 S.n16020 6.541
R30749 S.n15649 S.n15648 6.541
R30750 S.n15654 S.t4353 6.541
R30751 S.n15657 S.t3297 6.541
R30752 S.n15646 S.n15645 6.541
R30753 S.n15051 S.t4400 6.541
R30754 S.n14109 S.t604 6.541
R30755 S.n13734 S.n13733 6.541
R30756 S.n13742 S.t4081 6.541
R30757 S.n13745 S.t4341 6.541
R30758 S.n13737 S.n13736 6.541
R30759 S.n14142 S.n14141 6.541
R30760 S.n14149 S.t3613 6.541
R30761 S.n14146 S.t734 6.541
R30762 S.n14139 S.n14138 6.541
R30763 S.n22908 S.t2326 6.541
R30764 S.n22906 S.t3070 6.541
R30765 S.n22525 S.n22524 6.541
R30766 S.n22530 S.t1355 6.541
R30767 S.n22533 S.t619 6.541
R30768 S.n22522 S.n22521 6.541
R30769 S.n22113 S.n22112 6.541
R30770 S.n22120 S.t3317 6.541
R30771 S.n22117 S.t1759 6.541
R30772 S.n22110 S.n22109 6.541
R30773 S.n21502 S.n21501 6.541
R30774 S.n21507 S.t2342 6.541
R30775 S.n21510 S.t2206 6.541
R30776 S.n21499 S.n21498 6.541
R30777 S.n21835 S.n21834 6.541
R30778 S.n21839 S.t106 6.541
R30779 S.n21842 S.t3569 6.541
R30780 S.n21832 S.n21831 6.541
R30781 S.n20679 S.n20678 6.541
R30782 S.n20684 S.t1464 6.541
R30783 S.n20687 S.t2154 6.541
R30784 S.n20676 S.n20675 6.541
R30785 S.n21025 S.n21024 6.541
R30786 S.n21029 S.t13 6.541
R30787 S.n21032 S.t3516 6.541
R30788 S.n21022 S.n21021 6.541
R30789 S.n20068 S.n20067 6.541
R30790 S.n20073 S.t1412 6.541
R30791 S.n20076 S.t2107 6.541
R30792 S.n20065 S.n20064 6.541
R30793 S.n19621 S.n19620 6.541
R30794 S.n19628 S.t4566 6.541
R30795 S.n19625 S.t3470 6.541
R30796 S.n19618 S.n19617 6.541
R30797 S.n19214 S.n19213 6.541
R30798 S.n19219 S.t1357 6.541
R30799 S.n19222 S.t2057 6.541
R30800 S.n19211 S.n19210 6.541
R30801 S.n18749 S.n18748 6.541
R30802 S.n18756 S.t2982 6.541
R30803 S.n18753 S.t3424 6.541
R30804 S.n18746 S.n18745 6.541
R30805 S.n18348 S.n18347 6.541
R30806 S.n18353 S.t1298 6.541
R30807 S.n18356 S.t468 6.541
R30808 S.n18345 S.n18344 6.541
R30809 S.n17866 S.n17865 6.541
R30810 S.n17873 S.t2928 6.541
R30811 S.n17870 S.t3620 6.541
R30812 S.n17863 S.n17862 6.541
R30813 S.n17459 S.n17458 6.541
R30814 S.n17464 S.t1520 6.541
R30815 S.n17467 S.t423 6.541
R30816 S.n17456 S.n17455 6.541
R30817 S.n16957 S.n16956 6.541
R30818 S.n16964 S.t2878 6.541
R30819 S.n16961 S.t3562 6.541
R30820 S.n16954 S.n16953 6.541
R30821 S.n16557 S.n16556 6.541
R30822 S.n16562 S.t1459 6.541
R30823 S.n16565 S.t376 6.541
R30824 S.n16554 S.n16553 6.541
R30825 S.n16039 S.n16038 6.541
R30826 S.n16046 S.t2821 6.541
R30827 S.n16043 S.t3511 6.541
R30828 S.n16036 S.n16035 6.541
R30829 S.n15633 S.n15632 6.541
R30830 S.n15638 S.t1405 6.541
R30831 S.n15641 S.t331 6.541
R30832 S.n15630 S.n15629 6.541
R30833 S.n15095 S.n15094 6.541
R30834 S.n15102 S.t2768 6.541
R30835 S.n15099 S.t3466 6.541
R30836 S.n15092 S.n15091 6.541
R30837 S.n14696 S.n14695 6.541
R30838 S.n14701 S.t1352 6.541
R30839 S.n14704 S.t1102 6.541
R30840 S.n14693 S.n14692 6.541
R30841 S.n14113 S.t1396 6.541
R30842 S.n13145 S.t3054 6.541
R30843 S.n12746 S.n12745 6.541
R30844 S.n12754 S.t2064 6.541
R30845 S.n12757 S.t2365 6.541
R30846 S.n12749 S.n12748 6.541
R30847 S.n13178 S.n13177 6.541
R30848 S.n13185 S.t601 6.541
R30849 S.n13182 S.t3185 6.541
R30850 S.n13175 S.n13174 6.541
R30851 S.n22901 S.t3864 6.541
R30852 S.n22899 S.t42 6.541
R30853 S.n22509 S.n22508 6.541
R30854 S.n22514 S.t2920 6.541
R30855 S.n22517 S.t2181 6.541
R30856 S.n22506 S.n22505 6.541
R30857 S.n22128 S.n22127 6.541
R30858 S.n22135 S.t89 6.541
R30859 S.n22132 S.t3310 6.541
R30860 S.n22125 S.n22124 6.541
R30861 S.n21486 S.n21485 6.541
R30862 S.n21491 S.t3878 6.541
R30863 S.n21494 S.t1466 6.541
R30864 S.n21483 S.n21482 6.541
R30865 S.n21820 S.n21819 6.541
R30866 S.n21824 S.t4124 6.541
R30867 S.n21827 S.t2281 6.541
R30868 S.n21817 S.n21816 6.541
R30869 S.n20663 S.n20662 6.541
R30870 S.n20668 S.t2820 6.541
R30871 S.n20671 S.t3700 6.541
R30872 S.n20660 S.n20659 6.541
R30873 S.n21010 S.n21009 6.541
R30874 S.n21014 S.t1659 6.541
R30875 S.n21017 S.t563 6.541
R30876 S.n21007 S.n21006 6.541
R30877 S.n20052 S.n20051 6.541
R30878 S.n20057 S.t2980 6.541
R30879 S.n20060 S.t3655 6.541
R30880 S.n20049 S.n20048 6.541
R30881 S.n19636 S.n19635 6.541
R30882 S.n19643 S.t1607 6.541
R30883 S.n19640 S.t512 6.541
R30884 S.n19633 S.n19632 6.541
R30885 S.n19198 S.n19197 6.541
R30886 S.n19203 S.t2922 6.541
R30887 S.n19206 S.t3612 6.541
R30888 S.n19195 S.n19194 6.541
R30889 S.n18764 S.n18763 6.541
R30890 S.n18771 S.t4541 6.541
R30891 S.n18768 S.t462 6.541
R30892 S.n18761 S.n18760 6.541
R30893 S.n18332 S.n18331 6.541
R30894 S.n18337 S.t2867 6.541
R30895 S.n18340 S.t2029 6.541
R30896 S.n18329 S.n18328 6.541
R30897 S.n17881 S.n17880 6.541
R30898 S.n17888 S.t4482 6.541
R30899 S.n17885 S.t421 6.541
R30900 S.n17878 S.n17877 6.541
R30901 S.n17443 S.n17442 6.541
R30902 S.n17448 S.t2816 6.541
R30903 S.n17451 S.t1980 6.541
R30904 S.n17440 S.n17439 6.541
R30905 S.n16972 S.n16971 6.541
R30906 S.n16979 S.t4434 6.541
R30907 S.n16976 S.t611 6.541
R30908 S.n16969 S.n16968 6.541
R30909 S.n16541 S.n16540 6.541
R30910 S.n16546 S.t3019 6.541
R30911 S.n16549 S.t1936 6.541
R30912 S.n16538 S.n16537 6.541
R30913 S.n16054 S.n16053 6.541
R30914 S.n16061 S.t4375 6.541
R30915 S.n16058 S.t555 6.541
R30916 S.n16051 S.n16050 6.541
R30917 S.n15617 S.n15616 6.541
R30918 S.n15622 S.t2973 6.541
R30919 S.n15625 S.t1891 6.541
R30920 S.n15614 S.n15613 6.541
R30921 S.n15110 S.n15109 6.541
R30922 S.n15117 S.t4324 6.541
R30923 S.n15114 S.t506 6.541
R30924 S.n15107 S.n15106 6.541
R30925 S.n14680 S.n14679 6.541
R30926 S.n14685 S.t2917 6.541
R30927 S.n14688 S.t2662 6.541
R30928 S.n14677 S.n14676 6.541
R30929 S.n14157 S.n14156 6.541
R30930 S.n14164 S.t653 6.541
R30931 S.n14161 S.t4269 6.541
R30932 S.n14154 S.n14153 6.541
R30933 S.n13721 S.n13720 6.541
R30934 S.n13726 S.t2219 6.541
R30935 S.n13729 S.t2610 6.541
R30936 S.n13718 S.n13717 6.541
R30937 S.n13149 S.t2910 6.541
R30938 S.n12172 S.t960 6.541
R30939 S.n11736 S.n11735 6.541
R30940 S.n11744 S.t4508 6.541
R30941 S.n11747 S.t342 6.541
R30942 S.n11739 S.n11738 6.541
R30943 S.n12205 S.n12204 6.541
R30944 S.n12212 S.t2113 6.541
R30945 S.n12209 S.t1066 6.541
R30946 S.n12202 S.n12201 6.541
R30947 S.n22894 S.t901 6.541
R30948 S.n22892 S.t1671 6.541
R30949 S.n22493 S.n22492 6.541
R30950 S.n22498 S.t4474 6.541
R30951 S.n22501 S.t3724 6.541
R30952 S.n22490 S.n22489 6.541
R30953 S.n22143 S.n22142 6.541
R30954 S.n22150 S.t1694 6.541
R30955 S.n22147 S.t340 6.541
R30956 S.n22140 S.n22139 6.541
R30957 S.n21470 S.n21469 6.541
R30958 S.n21475 S.t914 6.541
R30959 S.n21478 S.t3022 6.541
R30960 S.n21467 S.n21466 6.541
R30961 S.n21805 S.n21804 6.541
R30962 S.n21809 S.t961 6.541
R30963 S.n21812 S.t3820 6.541
R30964 S.n21802 S.n21801 6.541
R30965 S.n20647 S.n20646 6.541
R30966 S.n20652 S.t4372 6.541
R30967 S.n20655 S.t1977 6.541
R30968 S.n20644 S.n20643 6.541
R30969 S.n20995 S.n20994 6.541
R30970 S.n20999 S.t146 6.541
R30971 S.n21002 S.t2741 6.541
R30972 S.n20992 S.n20991 6.541
R30973 S.n20036 S.n20035 6.541
R30974 S.n20041 S.t3349 6.541
R30975 S.n20044 S.t698 6.541
R30976 S.n20033 S.n20032 6.541
R30977 S.n19651 S.n19650 6.541
R30978 S.n19658 S.t3162 6.541
R30979 S.n19655 S.t2077 6.541
R30980 S.n19648 S.n19647 6.541
R30981 S.n19182 S.n19181 6.541
R30982 S.n19187 S.t4478 6.541
R30983 S.n19190 S.t655 6.541
R30984 S.n19179 S.n19178 6.541
R30985 S.n18779 S.n18778 6.541
R30986 S.n18786 S.t1588 6.541
R30987 S.n18783 S.t2025 6.541
R30988 S.n18776 S.n18775 6.541
R30989 S.n18316 S.n18315 6.541
R30990 S.n18321 S.t4422 6.541
R30991 S.n18324 S.t3579 6.541
R30992 S.n18313 S.n18312 6.541
R30993 S.n17896 S.n17895 6.541
R30994 S.n17903 S.t1536 6.541
R30995 S.n17900 S.t1975 6.541
R30996 S.n17893 S.n17892 6.541
R30997 S.n17427 S.n17426 6.541
R30998 S.n17432 S.t4368 6.541
R30999 S.n17435 S.t3527 6.541
R31000 S.n17424 S.n17423 6.541
R31001 S.n16987 S.n16986 6.541
R31002 S.n16994 S.t1486 6.541
R31003 S.n16991 S.t1933 6.541
R31004 S.n16984 S.n16983 6.541
R31005 S.n16525 S.n16524 6.541
R31006 S.n16530 S.t4316 6.541
R31007 S.n16533 S.t3484 6.541
R31008 S.n16522 S.n16521 6.541
R31009 S.n16069 S.n16068 6.541
R31010 S.n16076 S.t1429 6.541
R31011 S.n16073 S.t2118 6.541
R31012 S.n16066 S.n16065 6.541
R31013 S.n15601 S.n15600 6.541
R31014 S.n15606 S.t4533 6.541
R31015 S.n15609 S.t3437 6.541
R31016 S.n15598 S.n15597 6.541
R31017 S.n15125 S.n15124 6.541
R31018 S.n15132 S.t1376 6.541
R31019 S.n15129 S.t2070 6.541
R31020 S.n15122 S.n15121 6.541
R31021 S.n14664 S.n14663 6.541
R31022 S.n14669 S.t4472 6.541
R31023 S.n14672 S.t4209 6.541
R31024 S.n14661 S.n14660 6.541
R31025 S.n14172 S.n14171 6.541
R31026 S.n14179 S.t2214 6.541
R31027 S.n14176 S.t1321 6.541
R31028 S.n14169 S.n14168 6.541
R31029 S.n13705 S.n13704 6.541
R31030 S.n13710 S.t3762 6.541
R31031 S.n13713 S.t4160 6.541
R31032 S.n13702 S.n13701 6.541
R31033 S.n13193 S.n13192 6.541
R31034 S.n13200 S.t2160 6.541
R31035 S.n13197 S.t1265 6.541
R31036 S.n13190 S.n13189 6.541
R31037 S.n12733 S.n12732 6.541
R31038 S.n12738 S.t3713 6.541
R31039 S.n12741 S.t4111 6.541
R31040 S.n12730 S.n12729 6.541
R31041 S.n12176 S.t4408 6.541
R31042 S.n11173 S.t3422 6.541
R31043 S.n10713 S.n10712 6.541
R31044 S.n10721 S.t2430 6.541
R31045 S.n10724 S.t2835 6.541
R31046 S.n10716 S.n10715 6.541
R31047 S.n11206 S.n11205 6.541
R31048 S.n11213 S.t3622 6.541
R31049 S.n11210 S.t3550 6.541
R31050 S.n11203 S.n11202 6.541
R31051 S.n22887 S.t2448 6.541
R31052 S.n22885 S.t3221 6.541
R31053 S.n22477 S.n22476 6.541
R31054 S.n22482 S.t1530 6.541
R31055 S.n22485 S.t770 6.541
R31056 S.n22474 S.n22473 6.541
R31057 S.n22158 S.n22157 6.541
R31058 S.n22165 S.t3249 6.541
R31059 S.n22162 S.t1902 6.541
R31060 S.n22155 S.n22154 6.541
R31061 S.n21454 S.n21453 6.541
R31062 S.n21459 S.t2459 6.541
R31063 S.n21462 S.t4582 6.541
R31064 S.n21451 S.n21450 6.541
R31065 S.n21790 S.n21789 6.541
R31066 S.n21794 S.t2509 6.541
R31067 S.n21797 S.t861 6.541
R31068 S.n21787 S.n21786 6.541
R31069 S.n20631 S.n20630 6.541
R31070 S.n20636 S.t1426 6.541
R31071 S.n20639 S.t3525 6.541
R31072 S.n20628 S.n20627 6.541
R31073 S.n20980 S.n20979 6.541
R31074 S.n20984 S.t1502 6.541
R31075 S.n20987 S.t4299 6.541
R31076 S.n20977 S.n20976 6.541
R31077 S.n20020 S.n20019 6.541
R31078 S.n20025 S.t382 6.541
R31079 S.n20028 S.t2474 6.541
R31080 S.n20017 S.n20016 6.541
R31081 S.n19666 S.n19665 6.541
R31082 S.n19673 S.t686 6.541
R31083 S.n19670 S.t3290 6.541
R31084 S.n19663 S.n19662 6.541
R31085 S.n19166 S.n19165 6.541
R31086 S.n19171 S.t3860 6.541
R31087 S.n19174 S.t2216 6.541
R31088 S.n19163 S.n19162 6.541
R31089 S.n18794 S.n18793 6.541
R31090 S.n18801 S.t3143 6.541
R31091 S.n18798 S.t3576 6.541
R31092 S.n18791 S.n18790 6.541
R31093 S.n18300 S.n18299 6.541
R31094 S.n18305 S.t1475 6.541
R31095 S.n18308 S.t629 6.541
R31096 S.n18297 S.n18296 6.541
R31097 S.n17911 S.n17910 6.541
R31098 S.n17918 S.t3090 6.541
R31099 S.n17915 S.t3523 6.541
R31100 S.n17908 S.n17907 6.541
R31101 S.n17411 S.n17410 6.541
R31102 S.n17416 S.t1422 6.541
R31103 S.n17419 S.t575 6.541
R31104 S.n17408 S.n17407 6.541
R31105 S.n17002 S.n17001 6.541
R31106 S.n17009 S.t3043 6.541
R31107 S.n17006 S.t3479 6.541
R31108 S.n16999 S.n16998 6.541
R31109 S.n16509 S.n16508 6.541
R31110 S.n16514 S.t1368 6.541
R31111 S.n16517 S.t525 6.541
R31112 S.n16506 S.n16505 6.541
R31113 S.n16084 S.n16083 6.541
R31114 S.n16091 S.t2989 6.541
R31115 S.n16088 S.t3433 6.541
R31116 S.n16081 S.n16080 6.541
R31117 S.n15585 S.n15584 6.541
R31118 S.n15590 S.t1314 6.541
R31119 S.n15593 S.t475 6.541
R31120 S.n15582 S.n15581 6.541
R31121 S.n15140 S.n15139 6.541
R31122 S.n15147 S.t2941 6.541
R31123 S.n15144 S.t3625 6.541
R31124 S.n15137 S.n15136 6.541
R31125 S.n14648 S.n14647 6.541
R31126 S.n14653 S.t1527 6.541
R31127 S.n14656 S.t1259 6.541
R31128 S.n14645 S.n14644 6.541
R31129 S.n14187 S.n14186 6.541
R31130 S.n14194 S.t3757 6.541
R31131 S.n14191 S.t2886 6.541
R31132 S.n14184 S.n14183 6.541
R31133 S.n13689 S.n13688 6.541
R31134 S.n13694 S.t806 6.541
R31135 S.n13697 S.t1207 6.541
R31136 S.n13686 S.n13685 6.541
R31137 S.n13208 S.n13207 6.541
R31138 S.n13215 S.t3706 6.541
R31139 S.n13212 S.t2834 6.541
R31140 S.n13205 S.n13204 6.541
R31141 S.n12717 S.n12716 6.541
R31142 S.n12722 S.t758 6.541
R31143 S.n12725 S.t1158 6.541
R31144 S.n12714 S.n12713 6.541
R31145 S.n12220 S.n12219 6.541
R31146 S.n12227 S.t3662 6.541
R31147 S.n12224 S.t2777 6.541
R31148 S.n12217 S.n12216 6.541
R31149 S.n11723 S.n11722 6.541
R31150 S.n11728 S.t706 6.541
R31151 S.n11731 S.t1110 6.541
R31152 S.n11720 S.n11719 6.541
R31153 S.n11177 S.t1402 6.541
R31154 S.n10165 S.t2477 6.541
R31155 S.n9668 S.n9667 6.541
R31156 S.n9676 S.t367 6.541
R31157 S.n9679 S.t843 6.541
R31158 S.n9671 S.n9670 6.541
R31159 S.n10198 S.n10197 6.541
R31160 S.n10205 S.t614 6.541
R31161 S.n10202 S.t1493 6.541
R31162 S.n10195 S.n10194 6.541
R31163 S.n22880 S.t3987 6.541
R31164 S.n22878 S.t242 6.541
R31165 S.n22461 S.n22460 6.541
R31166 S.n22466 S.t3084 6.541
R31167 S.n22469 S.t2324 6.541
R31168 S.n22458 S.n22457 6.541
R31169 S.n22173 S.n22172 6.541
R31170 S.n22180 S.t272 6.541
R31171 S.n22177 S.t3446 6.541
R31172 S.n22170 S.n22169 6.541
R31173 S.n21438 S.n21437 6.541
R31174 S.n21443 S.t4001 6.541
R31175 S.n21446 S.t1628 6.541
R31176 S.n21435 S.n21434 6.541
R31177 S.n21775 S.n21774 6.541
R31178 S.n21779 S.t4052 6.541
R31179 S.n21782 S.t2407 6.541
R31180 S.n21772 S.n21771 6.541
R31181 S.n20615 S.n20614 6.541
R31182 S.n20620 S.t2988 6.541
R31183 S.n20623 S.t570 6.541
R31184 S.n20612 S.n20611 6.541
R31185 S.n20965 S.n20964 6.541
R31186 S.n20969 S.t3055 6.541
R31187 S.n20972 S.t1351 6.541
R31188 S.n20962 S.n20961 6.541
R31189 S.n20004 S.n20003 6.541
R31190 S.n20009 S.t1941 6.541
R31191 S.n20012 S.t4011 6.541
R31192 S.n20001 S.n20000 6.541
R31193 S.n19681 S.n19680 6.541
R31194 S.n19688 S.t2008 6.541
R31195 S.n19685 S.t319 6.541
R31196 S.n19678 S.n19677 6.541
R31197 S.n19150 S.n19149 6.541
R31198 S.n19155 S.t895 6.541
R31199 S.n19158 S.t3006 6.541
R31200 S.n19147 S.n19146 6.541
R31201 S.n18809 S.n18808 6.541
R31202 S.n18816 S.t1711 6.541
R31203 S.n18813 S.t3803 6.541
R31204 S.n18806 S.n18805 6.541
R31205 S.n18284 S.n18283 6.541
R31206 S.n18289 S.t4354 6.541
R31207 S.n18292 S.t2188 6.541
R31208 S.n18281 S.n18280 6.541
R31209 S.n17926 S.n17925 6.541
R31210 S.n17933 S.t78 6.541
R31211 S.n17930 S.t569 6.541
R31212 S.n17923 S.n17922 6.541
R31213 S.n17395 S.n17394 6.541
R31214 S.n17400 S.t2986 6.541
R31215 S.n17403 S.t2139 6.541
R31216 S.n17392 S.n17391 6.541
R31217 S.n17017 S.n17016 6.541
R31218 S.n17024 S.t4601 6.541
R31219 S.n17021 S.t522 6.541
R31220 S.n17014 S.n17013 6.541
R31221 S.n16493 S.n16492 6.541
R31222 S.n16498 S.t2932 6.541
R31223 S.n16501 S.t2091 6.541
R31224 S.n16490 S.n16489 6.541
R31225 S.n16099 S.n16098 6.541
R31226 S.n16106 S.t4550 6.541
R31227 S.n16103 S.t472 6.541
R31228 S.n16096 S.n16095 6.541
R31229 S.n15569 S.n15568 6.541
R31230 S.n15574 S.t2882 6.541
R31231 S.n15577 S.t2037 6.541
R31232 S.n15566 S.n15565 6.541
R31233 S.n15155 S.n15154 6.541
R31234 S.n15162 S.t4497 6.541
R31235 S.n15159 S.t426 6.541
R31236 S.n15152 S.n15151 6.541
R31237 S.n14632 S.n14631 6.541
R31238 S.n14637 S.t2826 6.541
R31239 S.n14640 S.t2827 6.541
R31240 S.n14629 S.n14628 6.541
R31241 S.n14202 S.n14201 6.541
R31242 S.n14209 S.t803 6.541
R31243 S.n14206 S.t4443 6.541
R31244 S.n14199 S.n14198 6.541
R31245 S.n13673 S.n13672 6.541
R31246 S.n13678 S.t2360 6.541
R31247 S.n13681 S.t2771 6.541
R31248 S.n13670 S.n13669 6.541
R31249 S.n13223 S.n13222 6.541
R31250 S.n13230 S.t750 6.541
R31251 S.n13227 S.t4387 6.541
R31252 S.n13220 S.n13219 6.541
R31253 S.n12701 S.n12700 6.541
R31254 S.n12706 S.t2318 6.541
R31255 S.n12709 S.t2717 6.541
R31256 S.n12698 S.n12697 6.541
R31257 S.n12235 S.n12234 6.541
R31258 S.n12242 S.t701 6.541
R31259 S.n12239 S.t4329 6.541
R31260 S.n12232 S.n12231 6.541
R31261 S.n11707 S.n11706 6.541
R31262 S.n11712 S.t2270 6.541
R31263 S.n11715 S.t2669 6.541
R31264 S.n11704 S.n11703 6.541
R31265 S.n11221 S.n11220 6.541
R31266 S.n11228 S.t664 6.541
R31267 S.n11225 S.t4281 6.541
R31268 S.n11218 S.n11217 6.541
R31269 S.n10700 S.n10699 6.541
R31270 S.n10705 S.t2227 6.541
R31271 S.n10708 S.t2619 6.541
R31272 S.n10697 S.n10696 6.541
R31273 S.n10169 S.t2915 6.541
R31274 S.n9131 S.t424 6.541
R31275 S.n8610 S.n8609 6.541
R31276 S.n8618 S.t2794 6.541
R31277 S.n8621 S.t2197 6.541
R31278 S.n8613 S.n8612 6.541
R31279 S.n9164 S.n9163 6.541
R31280 S.n9171 S.t585 6.541
R31281 S.n9168 S.t3922 6.541
R31282 S.n9161 S.n9160 6.541
R31283 S.n22873 S.t828 6.541
R31284 S.n22871 S.t1810 6.541
R31285 S.n22445 S.n22444 6.541
R31286 S.n22450 S.t4384 6.541
R31287 S.n22453 S.t3861 6.541
R31288 S.n22442 S.n22441 6.541
R31289 S.n22188 S.n22187 6.541
R31290 S.n22195 S.t1836 6.541
R31291 S.n22192 S.t486 6.541
R31292 S.n22185 S.n22184 6.541
R31293 S.n21422 S.n21421 6.541
R31294 S.n21427 S.t1035 6.541
R31295 S.n21430 S.t3181 6.541
R31296 S.n21419 S.n21418 6.541
R31297 S.n21760 S.n21759 6.541
R31298 S.n21764 S.t1088 6.541
R31299 S.n21767 S.t3946 6.541
R31300 S.n21757 S.n21756 6.541
R31301 S.n20599 S.n20598 6.541
R31302 S.n20604 S.t4548 6.541
R31303 S.n20607 S.t2136 6.541
R31304 S.n20596 S.n20595 6.541
R31305 S.n20950 S.n20949 6.541
R31306 S.n20954 S.t8 6.541
R31307 S.n20957 S.t2916 6.541
R31308 S.n20947 S.n20946 6.541
R31309 S.n19988 S.n19987 6.541
R31310 S.n19993 S.t3488 6.541
R31311 S.n19996 S.t1044 6.541
R31312 S.n19985 S.n19984 6.541
R31313 S.n19696 S.n19695 6.541
R31314 S.n19703 S.t3558 6.541
R31315 S.n19700 S.t1881 6.541
R31316 S.n19693 S.n19692 6.541
R31317 S.n19134 S.n19133 6.541
R31318 S.n19139 S.t2442 6.541
R31319 S.n19142 S.t4564 6.541
R31320 S.n19131 S.n19130 6.541
R31321 S.n18824 S.n18823 6.541
R31322 S.n18831 S.t3030 6.541
R31323 S.n18828 S.t838 6.541
R31324 S.n18821 S.n18820 6.541
R31325 S.n18268 S.n18267 6.541
R31326 S.n18273 S.t1403 6.541
R31327 S.n18276 S.t3994 6.541
R31328 S.n18265 S.n18264 6.541
R31329 S.n17941 S.n17940 6.541
R31330 S.n17948 S.t2229 6.541
R31331 S.n17945 S.t4279 6.541
R31332 S.n17938 S.n17937 6.541
R31333 S.n17379 S.n17378 6.541
R31334 S.n17384 S.t368 6.541
R31335 S.n17387 S.t3686 6.541
R31336 S.n17376 S.n17375 6.541
R31337 S.n17032 S.n17031 6.541
R31338 S.n17039 S.t1647 6.541
R31339 S.n17036 S.t2086 6.541
R31340 S.n17029 S.n17028 6.541
R31341 S.n16477 S.n16476 6.541
R31342 S.n16482 S.t4490 6.541
R31343 S.n16485 S.t3640 6.541
R31344 S.n16474 S.n16473 6.541
R31345 S.n16114 S.n16113 6.541
R31346 S.n16121 S.t1595 6.541
R31347 S.n16118 S.t2035 6.541
R31348 S.n16111 S.n16110 6.541
R31349 S.n15553 S.n15552 6.541
R31350 S.n15558 S.t4439 6.541
R31351 S.n15561 S.t3593 6.541
R31352 S.n15550 S.n15549 6.541
R31353 S.n15170 S.n15169 6.541
R31354 S.n15177 S.t1548 6.541
R31355 S.n15174 S.t1982 6.541
R31356 S.n15167 S.n15166 6.541
R31357 S.n14616 S.n14615 6.541
R31358 S.n14621 S.t4378 6.541
R31359 S.n14624 S.t4374 6.541
R31360 S.n14613 S.n14612 6.541
R31361 S.n14217 S.n14216 6.541
R31362 S.n14224 S.t2358 6.541
R31363 S.n14221 S.t1230 6.541
R31364 S.n14214 S.n14213 6.541
R31365 S.n13657 S.n13656 6.541
R31366 S.n13662 S.t3680 6.541
R31367 S.n13665 S.t4323 6.541
R31368 S.n13654 S.n13653 6.541
R31369 S.n13238 S.n13237 6.541
R31370 S.n13245 S.t2313 6.541
R31371 S.n13242 S.t1439 6.541
R31372 S.n13235 S.n13234 6.541
R31373 S.n12685 S.n12684 6.541
R31374 S.n12690 S.t3852 6.541
R31375 S.n12693 S.t4271 6.541
R31376 S.n12682 S.n12681 6.541
R31377 S.n12250 S.n12249 6.541
R31378 S.n12257 S.t2263 6.541
R31379 S.n12254 S.t1382 6.541
R31380 S.n12247 S.n12246 6.541
R31381 S.n11691 S.n11690 6.541
R31382 S.n11696 S.t3808 6.541
R31383 S.n11699 S.t4220 6.541
R31384 S.n11688 S.n11687 6.541
R31385 S.n11236 S.n11235 6.541
R31386 S.n11243 S.t2224 6.541
R31387 S.n11240 S.t1328 6.541
R31388 S.n11233 S.n11232 6.541
R31389 S.n10684 S.n10683 6.541
R31390 S.n10689 S.t3771 6.541
R31391 S.n10692 S.t4170 6.541
R31392 S.n10681 S.n10680 6.541
R31393 S.n10213 S.n10212 6.541
R31394 S.n10220 S.t2175 6.541
R31395 S.n10217 S.t1279 6.541
R31396 S.n10210 S.n10209 6.541
R31397 S.n9655 S.n9654 6.541
R31398 S.n9660 S.t3722 6.541
R31399 S.n9663 S.t4122 6.541
R31400 S.n9652 S.n9651 6.541
R31401 S.n9135 S.t4415 6.541
R31402 S.n8088 S.t2862 6.541
R31403 S.n7530 S.n7529 6.541
R31404 S.n7538 S.t766 6.541
R31405 S.n7541 S.t153 6.541
R31406 S.n7533 S.n7532 6.541
R31407 S.n8121 S.n8120 6.541
R31408 S.n8128 S.t2096 6.541
R31409 S.n8125 S.t1873 6.541
R31410 S.n8118 S.n8117 6.541
R31411 S.n22866 S.t2383 6.541
R31412 S.n22864 S.t3355 6.541
R31413 S.n22429 S.n22428 6.541
R31414 S.n22434 S.t1437 6.541
R31415 S.n22437 S.t896 6.541
R31416 S.n22426 S.n22425 6.541
R31417 S.n22203 S.n22202 6.541
R31418 S.n22210 S.t3381 6.541
R31419 S.n22207 S.t1826 6.541
R31420 S.n22200 S.n22199 6.541
R31421 S.n21406 S.n21405 6.541
R31422 S.n21411 S.t2396 6.541
R31423 S.n21414 S.t201 6.541
R31424 S.n21403 S.n21402 6.541
R31425 S.n21745 S.n21744 6.541
R31426 S.n21749 S.t2649 6.541
R31427 S.n21752 S.t982 6.541
R31428 S.n21742 S.n21741 6.541
R31429 S.n20583 S.n20582 6.541
R31430 S.n20588 S.t1591 6.541
R31431 S.n20591 S.t3683 6.541
R31432 S.n20580 S.n20579 6.541
R31433 S.n20935 S.n20934 6.541
R31434 S.n20939 S.t1656 6.541
R31435 S.n20942 S.t4470 6.541
R31436 S.n20932 S.n20931 6.541
R31437 S.n19972 S.n19971 6.541
R31438 S.n19977 S.t531 6.541
R31439 S.n19980 S.t2597 6.541
R31440 S.n19969 S.n19968 6.541
R31441 S.n19711 S.n19710 6.541
R31442 S.n19718 S.t602 6.541
R31443 S.n19715 S.t3427 6.541
R31444 S.n19708 S.n19707 6.541
R31445 S.n19118 S.n19117 6.541
R31446 S.n19123 S.t3984 6.541
R31447 S.n19126 S.t1604 6.541
R31448 S.n19115 S.n19114 6.541
R31449 S.n18839 S.n18838 6.541
R31450 S.n18846 S.t4592 6.541
R31451 S.n18843 S.t2391 6.541
R31452 S.n18836 S.n18835 6.541
R31453 S.n18252 S.n18251 6.541
R31454 S.n18257 S.t2971 6.541
R31455 S.n18260 S.t1031 6.541
R31456 S.n18249 S.n18248 6.541
R31457 S.n17956 S.n17955 6.541
R31458 S.n17963 S.t3531 6.541
R31459 S.n17960 S.t1330 6.541
R31460 S.n17953 S.n17952 6.541
R31461 S.n17363 S.n17362 6.541
R31462 S.n17368 S.t1926 6.541
R31463 S.n17371 S.t4543 6.541
R31464 S.n17360 S.n17359 6.541
R31465 S.n17047 S.n17046 6.541
R31466 S.n17054 S.t2688 6.541
R31467 S.n17051 S.t305 6.541
R31468 S.n17044 S.n17043 6.541
R31469 S.n16461 S.n16460 6.541
R31470 S.n16466 S.t881 6.541
R31471 S.n16469 S.t683 6.541
R31472 S.n16458 S.n16457 6.541
R31473 S.n16129 S.n16128 6.541
R31474 S.n16136 S.t3150 6.541
R31475 S.n16133 S.t3587 6.541
R31476 S.n16126 S.n16125 6.541
R31477 S.n15537 S.n15536 6.541
R31478 S.n15542 S.t1492 6.541
R31479 S.n15545 S.t639 6.541
R31480 S.n15534 S.n15533 6.541
R31481 S.n15185 S.n15184 6.541
R31482 S.n15192 S.t3101 6.541
R31483 S.n15189 S.t3529 6.541
R31484 S.n15182 S.n15181 6.541
R31485 S.n14600 S.n14599 6.541
R31486 S.n14605 S.t1432 6.541
R31487 S.n14608 S.t1428 6.541
R31488 S.n14597 S.n14596 6.541
R31489 S.n14232 S.n14231 6.541
R31490 S.n14239 S.t3894 6.541
R31491 S.n14236 S.t2790 6.541
R31492 S.n14229 S.n14228 6.541
R31493 S.n13641 S.n13640 6.541
R31494 S.n13646 S.t722 6.541
R31495 S.n13649 S.t1375 6.541
R31496 S.n13638 S.n13637 6.541
R31497 S.n13253 S.n13252 6.541
R31498 S.n13260 S.t3850 6.541
R31499 S.n13257 S.t2738 6.541
R31500 S.n13250 S.n13249 6.541
R31501 S.n12669 S.n12668 6.541
R31502 S.n12674 S.t674 6.541
R31503 S.n12677 S.t1320 6.541
R31504 S.n12666 S.n12665 6.541
R31505 S.n12265 S.n12264 6.541
R31506 S.n12272 S.t3805 6.541
R31507 S.n12269 S.t2947 6.541
R31508 S.n12262 S.n12261 6.541
R31509 S.n11675 S.n11674 6.541
R31510 S.n11680 S.t847 6.541
R31511 S.n11683 S.t1269 6.541
R31512 S.n11672 S.n11671 6.541
R31513 S.n11251 S.n11250 6.541
R31514 S.n11258 S.t3767 6.541
R31515 S.n11255 S.t2894 6.541
R31516 S.n11248 S.n11247 6.541
R31517 S.n10668 S.n10667 6.541
R31518 S.n10673 S.t810 6.541
R31519 S.n10676 S.t1218 6.541
R31520 S.n10665 S.n10664 6.541
R31521 S.n10228 S.n10227 6.541
R31522 S.n10235 S.t3719 6.541
R31523 S.n10232 S.t2842 6.541
R31524 S.n10225 S.n10224 6.541
R31525 S.n9639 S.n9638 6.541
R31526 S.n9644 S.t768 6.541
R31527 S.n9647 S.t1167 6.541
R31528 S.n9636 S.n9635 6.541
R31529 S.n9179 S.n9178 6.541
R31530 S.n9186 S.t2148 6.541
R31531 S.n9183 S.t2784 6.541
R31532 S.n9176 S.n9175 6.541
R31533 S.n8597 S.n8596 6.541
R31534 S.n8602 S.t717 6.541
R31535 S.n8605 S.t4099 6.541
R31536 S.n8594 S.n8593 6.541
R31537 S.n8092 S.t1414 6.541
R31538 S.n7019 S.t817 6.541
R31539 S.n6437 S.n6436 6.541
R31540 S.n6445 S.t3214 6.541
R31541 S.n6448 S.t2637 6.541
R31542 S.n6440 S.n6439 6.541
R31543 S.n7052 S.n7051 6.541
R31544 S.n7059 S.t3603 6.541
R31545 S.n7056 S.t4286 6.541
R31546 S.n7049 S.n7048 6.541
R31547 S.n22859 S.t3921 6.541
R31548 S.n22857 S.t392 6.541
R31549 S.n22413 S.n22412 6.541
R31550 S.n22418 S.t2998 6.541
R31551 S.n22421 S.t2443 6.541
R31552 S.n22410 S.n22409 6.541
R31553 S.n22218 S.n22217 6.541
R31554 S.n22225 S.t417 6.541
R31555 S.n22222 S.t3371 6.541
R31556 S.n22215 S.n22214 6.541
R31557 S.n21390 S.n21389 6.541
R31558 S.n21395 S.t3935 6.541
R31559 S.n21398 S.t1766 6.541
R31560 S.n21387 S.n21386 6.541
R31561 S.n21730 S.n21729 6.541
R31562 S.n21734 S.t4198 6.541
R31563 S.n21737 S.t2343 6.541
R31564 S.n21727 S.n21726 6.541
R31565 S.n20567 S.n20566 6.541
R31566 S.n20572 S.t2901 6.541
R31567 S.n20575 S.t724 6.541
R31568 S.n20564 S.n20563 6.541
R31569 S.n20920 S.n20919 6.541
R31570 S.n20924 S.t3206 6.541
R31571 S.n20927 S.t1525 6.541
R31572 S.n20917 S.n20916 6.541
R31573 S.n19956 S.n19955 6.541
R31574 S.n19961 S.t2098 6.541
R31575 S.n19964 S.t4146 6.541
R31576 S.n19953 S.n19952 6.541
R31577 S.n19726 S.n19725 6.541
R31578 S.n19733 S.t2166 6.541
R31579 S.n19730 S.t467 6.541
R31580 S.n19723 S.n19722 6.541
R31581 S.n19102 S.n19101 6.541
R31582 S.n19107 S.t1020 6.541
R31583 S.n19110 S.t3160 6.541
R31584 S.n19099 S.n19098 6.541
R31585 S.n18854 S.n18853 6.541
R31586 S.n18861 S.t1638 6.541
R31587 S.n18858 S.t3931 6.541
R31588 S.n18851 S.n18850 6.541
R31589 S.n18236 S.n18235 6.541
R31590 S.n18241 S.t4532 6.541
R31591 S.n18244 S.t2582 6.541
R31592 S.n18233 S.n18232 6.541
R31593 S.n17971 S.n17970 6.541
R31594 S.n17978 S.t580 6.541
R31595 S.n17975 S.t2891 6.541
R31596 S.n17968 S.n17967 6.541
R31597 S.n17347 S.n17346 6.541
R31598 S.n17352 S.t3473 6.541
R31599 S.n17355 S.t1585 6.541
R31600 S.n17344 S.n17343 6.541
R31601 S.n17062 S.n17061 6.541
R31602 S.n17069 S.t4017 6.541
R31603 S.n17066 S.t1866 6.541
R31604 S.n17059 S.n17058 6.541
R31605 S.n16445 S.n16444 6.541
R31606 S.n16450 S.t2428 6.541
R31607 S.n16453 S.t527 6.541
R31608 S.n16442 S.n16441 6.541
R31609 S.n16144 S.n16143 6.541
R31610 S.n16151 S.t3248 6.541
R31611 S.n16148 S.t820 6.541
R31612 S.n16141 S.n16140 6.541
R31613 S.n15521 S.n15520 6.541
R31614 S.n15526 S.t1383 6.541
R31615 S.n15529 S.t2203 6.541
R31616 S.n15518 S.n15517 6.541
R31617 S.n15200 S.n15199 6.541
R31618 S.n15207 S.t93 6.541
R31619 S.n15204 S.t578 6.541
R31620 S.n15197 S.n15196 6.541
R31621 S.n14584 S.n14583 6.541
R31622 S.n14589 S.t2996 6.541
R31623 S.n14592 S.t2991 6.541
R31624 S.n14581 S.n14580 6.541
R31625 S.n14247 S.n14246 6.541
R31626 S.n14254 S.t927 6.541
R31627 S.n14251 S.t4348 6.541
R31628 S.n14244 S.n14243 6.541
R31629 S.n13625 S.n13624 6.541
R31630 S.n13630 S.t2285 6.541
R31631 S.n13633 S.t2940 6.541
R31632 S.n13622 S.n13621 6.541
R31633 S.n13268 S.n13267 6.541
R31634 S.n13275 S.t886 6.541
R31635 S.n13272 S.t4294 6.541
R31636 S.n13265 S.n13264 6.541
R31637 S.n12653 S.n12652 6.541
R31638 S.n12658 S.t2236 6.541
R31639 S.n12661 S.t2889 6.541
R31640 S.n12650 S.n12649 6.541
R31641 S.n12280 S.n12279 6.541
R31642 S.n12287 S.t844 6.541
R31643 S.n12284 S.t4241 6.541
R31644 S.n12277 S.n12276 6.541
R31645 S.n11659 S.n11658 6.541
R31646 S.n11664 S.t2192 6.541
R31647 S.n11667 S.t2833 6.541
R31648 S.n11656 S.n11655 6.541
R31649 S.n11266 S.n11265 6.541
R31650 S.n11273 S.t808 6.541
R31651 S.n11270 S.t4451 6.541
R31652 S.n11263 S.n11262 6.541
R31653 S.n10652 S.n10651 6.541
R31654 S.n10657 S.t2364 6.541
R31655 S.n10660 S.t2776 6.541
R31656 S.n10649 S.n10648 6.541
R31657 S.n10243 S.n10242 6.541
R31658 S.n10250 S.t762 6.541
R31659 S.n10247 S.t4397 6.541
R31660 S.n10240 S.n10239 6.541
R31661 S.n9623 S.n9622 6.541
R31662 S.n9628 S.t2323 6.541
R31663 S.n9631 S.t2726 6.541
R31664 S.n9620 S.n9619 6.541
R31665 S.n9194 S.n9193 6.541
R31666 S.n9201 S.t3695 6.541
R31667 S.n9198 S.t4342 6.541
R31668 S.n9191 S.n9190 6.541
R31669 S.n8581 S.n8580 6.541
R31670 S.n8586 S.t2280 6.541
R31671 S.n8589 S.t1141 6.541
R31672 S.n8578 S.n8577 6.541
R31673 S.n8136 S.n8135 6.541
R31674 S.n8143 S.t3645 6.541
R31675 S.n8140 S.t4288 6.541
R31676 S.n8133 S.n8132 6.541
R31677 S.n7517 S.n7516 6.541
R31678 S.n7522 S.t2232 6.541
R31679 S.n7525 S.t1097 6.541
R31680 S.n7514 S.n7513 6.541
R31681 S.n7023 S.t2925 6.541
R31682 S.n5941 S.t1733 6.541
R31683 S.n5321 S.n5320 6.541
R31684 S.n5329 S.t1096 6.541
R31685 S.n5332 S.t1804 6.541
R31686 S.n5324 S.n5323 6.541
R31687 S.n5974 S.n5973 6.541
R31688 S.n5981 S.t594 6.541
R31689 S.n5978 S.t2261 6.541
R31690 S.n5971 S.n5970 6.541
R31691 S.n22852 S.t3087 6.541
R31692 S.n22850 S.t4018 6.541
R31693 S.n22397 S.n22396 6.541
R31694 S.n22402 S.t2146 6.541
R31695 S.n22405 S.t3985 6.541
R31696 S.n22394 S.n22393 6.541
R31697 S.n22233 S.n22232 6.541
R31698 S.n22240 S.t1972 6.541
R31699 S.n22237 S.t409 6.541
R31700 S.n22230 S.n22229 6.541
R31701 S.n21374 S.n21373 6.541
R31702 S.n21379 S.t967 6.541
R31703 S.n21382 S.t3316 6.541
R31704 S.n21371 S.n21370 6.541
R31705 S.n21715 S.n21714 6.541
R31706 S.n21719 S.t1241 6.541
R31707 S.n21722 S.t3879 6.541
R31708 S.n21712 S.n21711 6.541
R31709 S.n20551 S.n20550 6.541
R31710 S.n20556 S.t4457 6.541
R31711 S.n20559 S.t2288 6.541
R31712 S.n20548 S.n20547 6.541
R31713 S.n20905 S.n20904 6.541
R31714 S.n20909 S.t228 6.541
R31715 S.n20912 S.t2825 6.541
R31716 S.n20902 S.n20901 6.541
R31717 S.n19940 S.n19939 6.541
R31718 S.n19945 S.t3414 6.541
R31719 S.n19948 S.t1190 6.541
R31720 S.n19937 S.n19936 6.541
R31721 S.n19741 S.n19740 6.541
R31722 S.n19748 S.t3711 6.541
R31723 S.n19745 S.t2028 6.541
R31724 S.n19738 S.n19737 6.541
R31725 S.n19086 S.n19085 6.541
R31726 S.n19091 S.t2569 6.541
R31727 S.n19094 S.t175 6.541
R31728 S.n19083 S.n19082 6.541
R31729 S.n18869 S.n18868 6.541
R31730 S.n18876 S.t3189 6.541
R31731 S.n18873 S.t964 6.541
R31732 S.n18866 S.n18865 6.541
R31733 S.n18220 S.n18219 6.541
R31734 S.n18225 S.t1578 6.541
R31735 S.n18228 S.t4125 6.541
R31736 S.n18217 S.n18216 6.541
R31737 S.n17986 S.n17985 6.541
R31738 S.n17993 S.t2144 6.541
R31739 S.n17990 S.t4450 6.541
R31740 S.n17983 S.n17982 6.541
R31741 S.n17331 S.n17330 6.541
R31742 S.n17336 S.t515 6.541
R31743 S.n17339 S.t3144 6.541
R31744 S.n17328 S.n17327 6.541
R31745 S.n17077 S.n17076 6.541
R31746 S.n17084 S.t1050 6.541
R31747 S.n17081 S.t3409 6.541
R31748 S.n17074 S.n17073 6.541
R31749 S.n16429 S.n16428 6.541
R31750 S.n16434 S.t3969 6.541
R31751 S.n16437 S.t2093 6.541
R31752 S.n16426 S.n16425 6.541
R31753 S.n16159 S.n16158 6.541
R31754 S.n16166 S.t4574 6.541
R31755 S.n16163 S.t2376 6.541
R31756 S.n16156 S.n16155 6.541
R31757 S.n15505 S.n15504 6.541
R31758 S.n15510 S.t2948 6.541
R31759 S.n15513 S.t1015 6.541
R31760 S.n15502 S.n15501 6.541
R31761 S.n15215 S.n15214 6.541
R31762 S.n15222 S.t3752 6.541
R31763 S.n15219 S.t1304 6.541
R31764 S.n15212 S.n15211 6.541
R31765 S.n14568 S.n14567 6.541
R31766 S.n14573 S.t1908 6.541
R31767 S.n14576 S.t4553 6.541
R31768 S.n14565 S.n14564 6.541
R31769 S.n14262 S.n14261 6.541
R31770 S.n14269 S.t2473 6.541
R31771 S.n14266 S.t1398 6.541
R31772 S.n14259 S.n14258 6.541
R31773 S.n13609 S.n13608 6.541
R31774 S.n13614 S.t3821 6.541
R31775 S.n13617 S.t4498 6.541
R31776 S.n13606 S.n13605 6.541
R31777 S.n13283 S.n13282 6.541
R31778 S.n13290 S.t2434 6.541
R31779 S.n13287 S.t1347 6.541
R31780 S.n13280 S.n13279 6.541
R31781 S.n12637 S.n12636 6.541
R31782 S.n12642 S.t3780 6.541
R31783 S.n12645 S.t4446 6.541
R31784 S.n12634 S.n12633 6.541
R31785 S.n12295 S.n12294 6.541
R31786 S.n12302 S.t2398 6.541
R31787 S.n12299 S.t1289 6.541
R31788 S.n12292 S.n12291 6.541
R31789 S.n11643 S.n11642 6.541
R31790 S.n11648 S.t3738 6.541
R31791 S.n11651 S.t4390 6.541
R31792 S.n11640 S.n11639 6.541
R31793 S.n11281 S.n11280 6.541
R31794 S.n11288 S.t2362 6.541
R31795 S.n11285 S.t1237 6.541
R31796 S.n11278 S.n11277 6.541
R31797 S.n10636 S.n10635 6.541
R31798 S.n10641 S.t3688 6.541
R31799 S.n10644 S.t4333 6.541
R31800 S.n10633 S.n10632 6.541
R31801 S.n10258 S.n10257 6.541
R31802 S.n10265 S.t2320 6.541
R31803 S.n10262 S.t1450 6.541
R31804 S.n10255 S.n10254 6.541
R31805 S.n9607 S.n9606 6.541
R31806 S.n9612 S.t3859 6.541
R31807 S.n9615 S.t4280 6.541
R31808 S.n9604 S.n9603 6.541
R31809 S.n9209 S.n9208 6.541
R31810 S.n9216 S.t739 6.541
R31811 S.n9213 S.t1394 6.541
R31812 S.n9206 S.n9205 6.541
R31813 S.n8565 S.n8564 6.541
R31814 S.n8570 S.t3819 6.541
R31815 S.n8573 S.t2702 6.541
R31816 S.n8562 S.n8561 6.541
R31817 S.n8151 S.n8150 6.541
R31818 S.n8158 S.t690 6.541
R31819 S.n8155 S.t1339 6.541
R31820 S.n8148 S.n8147 6.541
R31821 S.n7501 S.n7500 6.541
R31822 S.n7506 S.t3777 6.541
R31823 S.n7509 S.t2658 6.541
R31824 S.n7498 S.n7497 6.541
R31825 S.n7067 S.n7066 6.541
R31826 S.n7074 S.t648 6.541
R31827 S.n7071 S.t1283 6.541
R31828 S.n7064 S.n7063 6.541
R31829 S.n6424 S.n6423 6.541
R31830 S.n6429 S.t3731 6.541
R31831 S.n6432 S.t2605 6.541
R31832 S.n6421 S.n6420 6.541
R31833 S.n5945 S.t427 6.541
R31834 S.n4835 S.t4128 6.541
R31835 S.n4192 S.n4191 6.541
R31836 S.n4200 S.t2058 6.541
R31837 S.n4203 S.t4272 6.541
R31838 S.n4195 S.n4194 6.541
R31839 S.n4869 S.n4868 6.541
R31840 S.n4876 S.t2576 6.541
R31841 S.n4873 S.t3180 6.541
R31842 S.n4866 S.n4865 6.541
R31843 S.n22845 S.t71 6.541
R31844 S.n22843 S.t1051 6.541
R31845 S.n22381 S.n22380 6.541
R31846 S.n22386 S.t3694 6.541
R31847 S.n22389 S.t3165 6.541
R31848 S.n22378 S.n22377 6.541
R31849 S.n22248 S.n22247 6.541
R31850 S.n22255 S.t1076 6.541
R31851 S.n22252 S.t4033 6.541
R31852 S.n22245 S.n22244 6.541
R31853 S.n21358 S.n21357 6.541
R31854 S.n21363 S.t101 6.541
R31855 S.n21366 S.t348 6.541
R31856 S.n21355 S.n21354 6.541
R31857 S.n21700 S.n21699 6.541
R31858 S.n21704 S.t2805 6.541
R31859 S.n21707 S.t916 6.541
R31860 S.n21697 S.n21696 6.541
R31861 S.n20535 S.n20534 6.541
R31862 S.n20540 S.t1512 6.541
R31863 S.n20543 S.t3826 6.541
R31864 S.n20532 S.n20531 6.541
R31865 S.n20890 S.n20889 6.541
R31866 S.n20894 S.t1794 6.541
R31867 S.n20897 S.t4373 6.541
R31868 S.n20887 S.n20886 6.541
R31869 S.n19924 S.n19923 6.541
R31870 S.n19929 S.t458 6.541
R31871 S.n19932 S.t2749 6.541
R31872 S.n19921 S.n19920 6.541
R31873 S.n19756 S.n19755 6.541
R31874 S.n19763 S.t755 6.541
R31875 S.n19760 S.t3351 6.541
R31876 S.n19753 S.n19752 6.541
R31877 S.n19070 S.n19069 6.541
R31878 S.n19075 S.t3917 6.541
R31879 S.n19078 S.t1745 6.541
R31880 S.n19067 S.n19066 6.541
R31881 S.n18884 S.n18883 6.541
R31882 S.n18891 S.t207 6.541
R31883 S.n18888 S.t2513 6.541
R31884 S.n18881 S.n18880 6.541
R31885 S.n18204 S.n18203 6.541
R31886 S.n18209 S.t3133 6.541
R31887 S.n18212 S.t1169 6.541
R31888 S.n18201 S.n18200 6.541
R31889 S.n18001 S.n18000 6.541
R31890 S.n18008 S.t3691 6.541
R31891 S.n18005 S.t1505 6.541
R31892 S.n17998 S.n17997 6.541
R31893 S.n17315 S.n17314 6.541
R31894 S.n17320 S.t2081 6.541
R31895 S.n17323 S.t149 6.541
R31896 S.n17312 S.n17311 6.541
R31897 S.n17092 S.n17091 6.541
R31898 S.n17099 S.t2604 6.541
R31899 S.n17096 S.t450 6.541
R31900 S.n17089 S.n17088 6.541
R31901 S.n16413 S.n16412 6.541
R31902 S.n16418 S.t1007 6.541
R31903 S.n16421 S.t3644 6.541
R31904 S.n16410 S.n16409 6.541
R31905 S.n16174 S.n16173 6.541
R31906 S.n16181 S.t1618 6.541
R31907 S.n16178 S.t3910 6.541
R31908 S.n16171 S.n16170 6.541
R31909 S.n15489 S.n15488 6.541
R31910 S.n15494 S.t4504 6.541
R31911 S.n15497 S.t2562 6.541
R31912 S.n15486 S.n15485 6.541
R31913 S.n15230 S.n15229 6.541
R31914 S.n15237 S.t561 6.541
R31915 S.n15234 S.t2871 6.541
R31916 S.n15227 S.n15226 6.541
R31917 S.n14552 S.n14551 6.541
R31918 S.n14557 S.t3452 6.541
R31919 S.n14560 S.t679 6.541
R31920 S.n14549 S.n14548 6.541
R31921 S.n14277 S.n14276 6.541
R31922 S.n14284 S.t3372 6.541
R31923 S.n14281 S.t1465 6.541
R31924 S.n14274 S.n14273 6.541
R31925 S.n13593 S.n13592 6.541
R31926 S.n13598 S.t2049 6.541
R31927 S.n13601 S.t1553 6.541
R31928 S.n13590 S.n13589 6.541
R31929 S.n13298 S.n13297 6.541
R31930 S.n13305 S.t3974 6.541
R31931 S.n13302 S.t2912 6.541
R31932 S.n13295 S.n13294 6.541
R31933 S.n12621 S.n12620 6.541
R31934 S.n12626 S.t818 6.541
R31935 S.n12629 S.t1499 6.541
R31936 S.n12618 S.n12617 6.541
R31937 S.n12310 S.n12309 6.541
R31938 S.n12317 S.t3936 6.541
R31939 S.n12314 S.t2856 6.541
R31940 S.n12307 S.n12306 6.541
R31941 S.n11627 S.n11626 6.541
R31942 S.n11632 S.t781 6.541
R31943 S.n11635 S.t1441 6.541
R31944 S.n11624 S.n11623 6.541
R31945 S.n11296 S.n11295 6.541
R31946 S.n11303 S.t3896 6.541
R31947 S.n11300 S.t2798 6.541
R31948 S.n11293 S.n11292 6.541
R31949 S.n10620 S.n10619 6.541
R31950 S.n10625 S.t731 6.541
R31951 S.n10628 S.t1384 6.541
R31952 S.n10617 S.n10616 6.541
R31953 S.n10273 S.n10272 6.541
R31954 S.n10280 S.t3857 6.541
R31955 S.n10277 S.t2743 6.541
R31956 S.n10270 S.n10269 6.541
R31957 S.n9591 S.n9590 6.541
R31958 S.n9596 S.t685 6.541
R31959 S.n9599 S.t1332 6.541
R31960 S.n9588 S.n9587 6.541
R31961 S.n9227 S.n9226 6.541
R31962 S.n9231 S.t2299 6.541
R31963 S.n9219 S.t2962 6.541
R31964 S.n9224 S.n9223 6.541
R31965 S.n8549 S.n8548 6.541
R31966 S.n8554 S.t859 6.541
R31967 S.n8557 S.t4252 6.541
R31968 S.n8546 S.n8545 6.541
R31969 S.n8166 S.n8165 6.541
R31970 S.n8173 S.t2246 6.541
R31971 S.n8170 S.t2906 6.541
R31972 S.n8163 S.n8162 6.541
R31973 S.n7485 S.n7484 6.541
R31974 S.n7490 S.t816 6.541
R31975 S.n7493 S.t4206 6.541
R31976 S.n7482 S.n7481 6.541
R31977 S.n7082 S.n7081 6.541
R31978 S.n7089 S.t2210 6.541
R31979 S.n7086 S.t2852 6.541
R31980 S.n7079 S.n7078 6.541
R31981 S.n6408 S.n6407 6.541
R31982 S.n6413 S.t774 6.541
R31983 S.n6416 S.t4153 6.541
R31984 S.n6405 S.n6404 6.541
R31985 S.n5989 S.n5988 6.541
R31986 S.n5996 S.t2156 6.541
R31987 S.n5993 S.t2793 6.541
R31988 S.n5986 S.n5985 6.541
R31989 S.n5308 S.n5307 6.541
R31990 S.n5313 S.t723 6.541
R31991 S.n5316 S.t119 6.541
R31992 S.n5305 S.n5304 6.541
R31993 S.n4839 S.t408 6.541
R31994 S.n3722 S.t2115 6.541
R31995 S.n3051 S.n3050 6.541
R31996 S.n3059 S.t1081 6.541
R31997 S.n3062 S.t2309 6.541
R31998 S.n3054 S.n3053 6.541
R31999 S.n3756 S.n3755 6.541
R32000 S.n3764 S.t4075 6.541
R32001 S.n3761 S.t2245 6.541
R32002 S.n3753 S.n3752 6.541
R32003 S.n22838 S.t1684 6.541
R32004 S.n22836 S.t2413 6.541
R32005 S.n22670 S.n22669 6.541
R32006 S.n22667 S.t737 6.541
R32007 S.n22664 S.t4475 6.541
R32008 S.n22268 S.n22267 6.541
R32009 S.n22263 S.n22262 6.541
R32010 S.n22680 S.t2632 6.541
R32011 S.n22677 S.t1065 6.541
R32012 S.n22260 S.n22259 6.541
R32013 S.n21683 S.n21682 6.541
R32014 S.n21680 S.t1698 6.541
R32015 S.n21677 S.t3982 6.541
R32016 S.n21674 S.n21673 6.541
R32017 S.n21669 S.n21668 6.541
R32018 S.n21689 S.t1969 6.541
R32019 S.n21692 S.t4588 6.541
R32020 S.n21666 S.n21665 6.541
R32021 S.n20520 S.n20519 6.541
R32022 S.n20524 S.t658 6.541
R32023 S.n20527 S.t864 6.541
R32024 S.n20517 S.n20516 6.541
R32025 S.n20874 S.n20873 6.541
R32026 S.n20879 S.t3339 6.541
R32027 S.n20882 S.t1427 6.541
R32028 S.n20871 S.n20870 6.541
R32029 S.n19909 S.n19908 6.541
R32030 S.n19913 S.t2016 6.541
R32031 S.n19916 S.t4309 6.541
R32032 S.n19906 S.n19905 6.541
R32033 S.n19771 S.n19770 6.541
R32034 S.n19779 S.t2316 6.541
R32035 S.n19776 S.t386 6.541
R32036 S.n19768 S.n19767 6.541
R32037 S.n19055 S.n19054 6.541
R32038 S.n19059 S.t953 6.541
R32039 S.n19062 S.t3295 6.541
R32040 S.n19052 S.n19051 6.541
R32041 S.n18899 S.n18898 6.541
R32042 S.n18907 S.t1774 6.541
R32043 S.n18904 S.t3862 6.541
R32044 S.n18896 S.n18895 6.541
R32045 S.n18189 S.n18188 6.541
R32046 S.n18193 S.t4437 6.541
R32047 S.n18196 S.t2730 6.541
R32048 S.n18186 S.n18185 6.541
R32049 S.n18016 S.n18015 6.541
R32050 S.n18024 S.t735 6.541
R32051 S.n18021 S.t3059 6.541
R32052 S.n18013 S.n18012 6.541
R32053 S.n17300 S.n17299 6.541
R32054 S.n17304 S.t3634 6.541
R32055 S.n17307 S.t1726 6.541
R32056 S.n17297 S.n17296 6.541
R32057 S.n17107 S.n17106 6.541
R32058 S.n17115 S.t4155 6.541
R32059 S.n17112 S.t2009 6.541
R32060 S.n17104 S.n17103 6.541
R32061 S.n16398 S.n16397 6.541
R32062 S.n16402 S.t2551 6.541
R32063 S.n16405 S.t687 6.541
R32064 S.n16395 S.n16394 6.541
R32065 S.n16189 S.n16188 6.541
R32066 S.n16197 S.t3171 6.541
R32067 S.n16194 S.t948 6.541
R32068 S.n16186 S.n16185 6.541
R32069 S.n15474 S.n15473 6.541
R32070 S.n15478 S.t1559 6.541
R32071 S.n15481 S.t4105 6.541
R32072 S.n15471 S.n15470 6.541
R32073 S.n15245 S.n15244 6.541
R32074 S.n15253 S.t2128 6.541
R32075 S.n15250 S.t4427 6.541
R32076 S.n15242 S.n15241 6.541
R32077 S.n14537 S.n14536 6.541
R32078 S.n14541 S.t494 6.541
R32079 S.n14544 S.t2240 6.541
R32080 S.n14534 S.n14533 6.541
R32081 S.n14292 S.n14291 6.541
R32082 S.n14300 S.t178 6.541
R32083 S.n14297 S.t3025 6.541
R32084 S.n14289 S.n14288 6.541
R32085 S.n13578 S.n13577 6.541
R32086 S.n13582 S.t3604 6.541
R32087 S.n13585 S.t1143 6.541
R32088 S.n13575 S.n13574 6.541
R32089 S.n13313 S.n13312 6.541
R32090 S.n13321 S.t3883 6.541
R32091 S.n13318 S.t1979 6.541
R32092 S.n13310 S.n13309 6.541
R32093 S.n12606 S.n12605 6.541
R32094 S.n12610 S.t2529 6.541
R32095 S.n12613 S.t3052 6.541
R32096 S.n12603 S.n12602 6.541
R32097 S.n12325 S.n12324 6.541
R32098 S.n12333 S.t969 6.541
R32099 S.n12330 S.t4409 6.541
R32100 S.n12322 S.n12321 6.541
R32101 S.n11612 S.n11611 6.541
R32102 S.n11616 S.t2337 6.541
R32103 S.n11619 S.t3003 6.541
R32104 S.n11609 S.n11608 6.541
R32105 S.n11311 S.n11310 6.541
R32106 S.n11319 S.t929 6.541
R32107 S.n11316 S.t4357 6.541
R32108 S.n11308 S.n11307 6.541
R32109 S.n10605 S.n10604 6.541
R32110 S.n10609 S.t2290 6.541
R32111 S.n10612 S.t2949 6.541
R32112 S.n10602 S.n10601 6.541
R32113 S.n10288 S.n10287 6.541
R32114 S.n10296 S.t893 6.541
R32115 S.n10293 S.t4300 6.541
R32116 S.n10285 S.n10284 6.541
R32117 S.n9576 S.n9575 6.541
R32118 S.n9580 S.t2241 6.541
R32119 S.n9583 S.t2898 6.541
R32120 S.n9573 S.n9572 6.541
R32121 S.n9239 S.n9238 6.541
R32122 S.n9247 S.t3836 6.541
R32123 S.n9244 S.t4246 6.541
R32124 S.n9236 S.n9235 6.541
R32125 S.n8534 S.n8533 6.541
R32126 S.n8538 S.t2204 6.541
R32127 S.n8541 S.t1303 6.541
R32128 S.n8531 S.n8530 6.541
R32129 S.n8181 S.n8180 6.541
R32130 S.n8189 S.t3789 6.541
R32131 S.n8186 S.t4462 6.541
R32132 S.n8178 S.n8177 6.541
R32133 S.n7470 S.n7469 6.541
R32134 S.n7474 S.t2372 6.541
R32135 S.n7477 S.t1253 6.541
R32136 S.n7467 S.n7466 6.541
R32137 S.n7097 S.n7096 6.541
R32138 S.n7105 S.t3747 6.541
R32139 S.n7102 S.t4405 6.541
R32140 S.n7094 S.n7093 6.541
R32141 S.n6393 S.n6392 6.541
R32142 S.n6397 S.t2330 6.541
R32143 S.n6400 S.t1199 6.541
R32144 S.n6390 S.n6389 6.541
R32145 S.n6004 S.n6003 6.541
R32146 S.n6012 S.t3703 6.541
R32147 S.n6009 S.t4351 6.541
R32148 S.n6001 S.n6000 6.541
R32149 S.n5293 S.n5292 6.541
R32150 S.n5297 S.t2286 6.541
R32151 S.n5300 S.t1710 6.541
R32152 S.n5290 S.n5289 6.541
R32153 S.n4884 S.n4883 6.541
R32154 S.n4892 S.t4118 6.541
R32155 S.n4889 S.t316 6.541
R32156 S.n4881 S.n4880 6.541
R32157 S.n4180 S.n4179 6.541
R32158 S.n4184 S.t2699 6.541
R32159 S.n4187 S.t1670 6.541
R32160 S.n4177 S.n4176 6.541
R32161 S.n3726 S.t1919 6.541
R32162 S.n2591 S.t4562 6.541
R32163 S.n1444 S.n1443 6.541
R32164 S.n1890 S.t3567 6.541
R32165 S.n1893 S.t286 6.541
R32166 S.n1896 S.n1895 6.541
R32167 S.n2625 S.n2624 6.541
R32168 S.n2633 S.t1070 6.541
R32169 S.n2630 S.t144 6.541
R32170 S.n2622 S.n2621 6.541
R32171 S.n22829 S.t3235 6.541
R32172 S.n22827 S.t3951 6.541
R32173 S.n22364 S.n22363 6.541
R32174 S.n22370 S.t2302 6.541
R32175 S.n22373 S.t1531 6.541
R32176 S.n22361 S.n22360 6.541
R32177 S.n22688 S.n22687 6.541
R32178 S.n22699 S.t3976 6.541
R32179 S.n22696 S.t2620 6.541
R32180 S.n22685 S.n22684 6.541
R32181 S.n21652 S.n21651 6.541
R32182 S.n21649 S.t3253 6.541
R32183 S.n21646 S.t822 6.541
R32184 S.n21279 S.n21278 6.541
R32185 S.n21274 S.n21273 6.541
R32186 S.n21658 S.t3518 6.541
R32187 S.n21661 S.t1633 6.541
R32188 S.n21271 S.n21270 6.541
R32189 S.n20505 S.n20504 6.541
R32190 S.n20509 S.t2217 6.541
R32191 S.n20512 S.t4529 6.541
R32192 S.n20502 S.n20501 6.541
R32193 S.n20858 S.n20857 6.541
R32194 S.n20863 S.t2464 6.541
R32195 S.n20866 S.t577 6.541
R32196 S.n20855 S.n20854 6.541
R32197 S.n19894 S.n19893 6.541
R32198 S.n19898 S.t1114 6.541
R32199 S.n19901 S.t1360 6.541
R32200 S.n19891 S.n19890 6.541
R32201 S.n19787 S.n19786 6.541
R32202 S.n19795 S.t3853 6.541
R32203 S.n19792 S.t1947 6.541
R32204 S.n19784 S.n19783 6.541
R32205 S.n19040 S.n19039 6.541
R32206 S.n19044 S.t2503 6.541
R32207 S.n19047 S.t328 6.541
R32208 S.n19037 S.n19036 6.541
R32209 S.n18915 S.n18914 6.541
R32210 S.n18923 S.t3325 6.541
R32211 S.n18920 S.t897 6.541
R32212 S.n18912 S.n18911 6.541
R32213 S.n18174 S.n18173 6.541
R32214 S.n18178 S.t1488 6.541
R32215 S.n18181 S.t4283 6.541
R32216 S.n18171 S.n18170 6.541
R32217 S.n18032 S.n18031 6.541
R32218 S.n18040 S.t2296 6.541
R32219 S.n18037 S.t4355 6.541
R32220 S.n18029 S.n18028 6.541
R32221 S.n17285 S.n17284 6.541
R32222 S.n17289 S.t438 6.541
R32223 S.n17292 S.t3277 6.541
R32224 S.n17282 S.n17281 6.541
R32225 S.n17123 S.n17122 6.541
R32226 S.n17131 S.t1201 6.541
R32227 S.n17128 S.t3560 6.541
R32228 S.n17120 S.n17119 6.541
R32229 S.n16383 S.n16382 6.541
R32230 S.n16387 S.t4092 6.541
R32231 S.n16390 S.t2244 6.541
R32232 S.n16380 S.n16379 6.541
R32233 S.n16205 S.n16204 6.541
R32234 S.n16213 S.t188 6.541
R32235 S.n16210 S.t2494 6.541
R32236 S.n16202 S.n16201 6.541
R32237 S.n15459 S.n15458 6.541
R32238 S.n15463 S.t3112 6.541
R32239 S.n15466 S.t1152 6.541
R32240 S.n15456 S.n15455 6.541
R32241 S.n15261 S.n15260 6.541
R32242 S.n15269 S.t3674 6.541
R32243 S.n15266 S.t1481 6.541
R32244 S.n15258 S.n15257 6.541
R32245 S.n14522 S.n14521 6.541
R32246 S.n14526 S.t2060 6.541
R32247 S.n14529 S.t3783 6.541
R32248 S.n14519 S.n14518 6.541
R32249 S.n14308 S.n14307 6.541
R32250 S.n14316 S.t1747 6.541
R32251 S.n14313 S.t4585 6.541
R32252 S.n14305 S.n14304 6.541
R32253 S.n13563 S.n13562 6.541
R32254 S.n13567 S.t649 6.541
R32255 S.n13570 S.t2703 6.541
R32256 S.n13560 S.n13559 6.541
R32257 S.n13329 S.n13328 6.541
R32258 S.n13337 S.t705 6.541
R32259 S.n13334 S.t3524 6.541
R32260 S.n13326 S.n13325 6.541
R32261 S.n12591 S.n12590 6.541
R32262 S.n12595 S.t4070 6.541
R32263 S.n12598 S.t1706 6.541
R32264 S.n12588 S.n12587 6.541
R32265 S.n12341 S.n12340 6.541
R32266 S.n12349 S.t4379 6.541
R32267 S.n12346 S.t2476 6.541
R32268 S.n12338 S.n12337 6.541
R32269 S.n11597 S.n11596 6.541
R32270 S.n11601 S.t3077 6.541
R32271 S.n11604 S.t4560 6.541
R32272 S.n11594 S.n11593 6.541
R32273 S.n11327 S.n11326 6.541
R32274 S.n11335 S.t2478 6.541
R32275 S.n11332 S.t1408 6.541
R32276 S.n11324 S.n11323 6.541
R32277 S.n10590 S.n10589 6.541
R32278 S.n10594 S.t3831 6.541
R32279 S.n10597 S.t4509 6.541
R32280 S.n10587 S.n10586 6.541
R32281 S.n10304 S.n10303 6.541
R32282 S.n10312 S.t2440 6.541
R32283 S.n10309 S.t1353 6.541
R32284 S.n10301 S.n10300 6.541
R32285 S.n9561 S.n9560 6.541
R32286 S.n9565 S.t3785 6.541
R32287 S.n9568 S.t4454 6.541
R32288 S.n9558 S.n9557 6.541
R32289 S.n9255 S.n9254 6.541
R32290 S.n9263 S.t875 6.541
R32291 S.n9260 S.t1296 6.541
R32292 S.n9252 S.n9251 6.541
R32293 S.n8519 S.n8518 6.541
R32294 S.n8523 S.t3742 6.541
R32295 S.n8526 S.t2870 6.541
R32296 S.n8516 S.n8515 6.541
R32297 S.n8197 S.n8196 6.541
R32298 S.n8205 S.t830 6.541
R32299 S.n8202 S.t1246 6.541
R32300 S.n8194 S.n8193 6.541
R32301 S.n7455 S.n7454 6.541
R32302 S.n7459 S.t3698 6.541
R32303 S.n7462 S.t2818 6.541
R32304 S.n7452 S.n7451 6.541
R32305 S.n7113 S.n7112 6.541
R32306 S.n7121 S.t794 6.541
R32307 S.n7118 S.t1456 6.541
R32308 S.n7110 S.n7109 6.541
R32309 S.n6378 S.n6377 6.541
R32310 S.n6382 S.t3868 6.541
R32311 S.n6385 S.t2762 6.541
R32312 S.n6375 S.n6374 6.541
R32313 S.n6020 S.n6019 6.541
R32314 S.n6028 S.t743 6.541
R32315 S.n6025 S.t1401 6.541
R32316 S.n6017 S.n6016 6.541
R32317 S.n5278 S.n5277 6.541
R32318 S.n5282 S.t3824 6.541
R32319 S.n5285 S.t3264 6.541
R32320 S.n5275 S.n5274 6.541
R32321 S.n4900 S.n4899 6.541
R32322 S.n4908 S.t1164 6.541
R32323 S.n4905 S.t1879 6.541
R32324 S.n4897 S.n4896 6.541
R32325 S.n4165 S.n4164 6.541
R32326 S.n4169 S.t4249 6.541
R32327 S.n4172 S.t3220 6.541
R32328 S.n4162 S.n4161 6.541
R32329 S.n3772 S.n3771 6.541
R32330 S.n3780 S.t1115 6.541
R32331 S.n3777 S.t298 6.541
R32332 S.n3769 S.n3768 6.541
R32333 S.n3039 S.n3038 6.541
R32334 S.n3043 S.t2676 6.541
R32335 S.n3046 S.t3175 6.541
R32336 S.n3036 S.n3035 6.541
R32337 S.n2595 S.t3421 6.541
R32338 S.n22816 S.t3926 6.541
R32339 S.n22815 S.t703 6.541
R32340 S.n22773 S.t3467 6.541
R32341 S.n22720 S.t546 6.541
R32342 S.n895 S.n894 6.541
R32343 S.n919 S.t4082 6.541
R32344 S.n916 S.t543 6.541
R32345 S.n898 S.n897 6.541
R32346 S.n1977 S.n1976 6.541
R32347 S.n1987 S.t4126 6.541
R32348 S.n1990 S.t3320 6.541
R32349 S.n1974 S.n1973 6.541
R32350 S.n22292 S.t63 6.541
R32351 S.n22728 S.n22727 6.541
R32352 S.n22746 S.t2558 6.541
R32353 S.n22743 S.t1221 6.541
R32354 S.n22725 S.n22724 6.541
R32355 S.n21308 S.n21307 6.541
R32356 S.n21319 S.t1843 6.541
R32357 S.n21316 S.t3914 6.541
R32358 S.n21305 S.n21304 6.541
R32359 S.n21207 S.n21206 6.541
R32360 S.n21222 S.t1894 6.541
R32361 S.n21219 S.t205 6.541
R32362 S.n21204 S.n21203 6.541
R32363 S.n20485 S.n20484 6.541
R32364 S.n20496 S.t802 6.541
R32365 S.n20493 S.t2876 6.541
R32366 S.n20482 S.n20481 6.541
R32367 S.n20388 S.n20387 6.541
R32368 S.n20403 S.t851 6.541
R32369 S.n20400 S.t3687 6.541
R32370 S.n20385 S.n20384 6.541
R32371 S.n19874 S.n19873 6.541
R32372 S.n19885 S.t4223 6.541
R32373 S.n19882 S.t1851 6.541
R32374 S.n19871 S.n19870 6.541
R32375 S.n20261 S.n20260 6.541
R32376 S.n20273 S.t4557 6.541
R32377 S.n20276 S.t2602 6.541
R32378 S.n20258 S.n20257 6.541
R32379 S.n19020 S.n19019 6.541
R32380 S.n19031 S.t3232 6.541
R32381 S.n19028 S.t1002 6.541
R32382 S.n19017 S.n19016 6.541
R32383 S.n19393 S.n19392 6.541
R32384 S.n19405 S.t3992 6.541
R32385 S.n19408 S.t1613 6.541
R32386 S.n19390 S.n19389 6.541
R32387 S.n18154 S.n18153 6.541
R32388 S.n18165 S.t2195 6.541
R32389 S.n18162 S.t2902 6.541
R32390 S.n18151 S.n18150 6.541
R32391 S.n18506 S.n18505 6.541
R32392 S.n18518 S.t872 6.541
R32393 S.n18521 S.t2974 6.541
R32394 S.n18503 S.n18502 6.541
R32395 S.n17265 S.n17264 6.541
R32396 S.n17276 S.t3543 6.541
R32397 S.n17273 S.t1871 6.541
R32398 S.n17262 S.n17261 6.541
R32399 S.n17606 S.n17605 6.541
R32400 S.n17618 S.t4319 6.541
R32401 S.n17621 S.t1927 6.541
R32402 S.n17603 S.n17602 6.541
R32403 S.n16363 S.n16362 6.541
R32404 S.n16374 S.t2484 6.541
R32405 S.n16371 S.t826 6.541
R32406 S.n16360 S.n16359 6.541
R32407 S.n16683 S.n16682 6.541
R32408 S.n16695 S.t3308 6.541
R32409 S.n16698 S.t884 6.541
R32410 S.n16680 S.n16679 6.541
R32411 S.n15439 S.n15438 6.541
R32412 S.n15450 S.t1462 6.541
R32413 S.n15447 S.t4263 6.541
R32414 S.n15436 S.n15435 6.541
R32415 S.n15748 S.n15747 6.541
R32416 S.n15760 S.t2277 6.541
R32417 S.n15763 S.t4593 6.541
R32418 S.n15745 S.n15744 6.541
R32419 S.n14502 S.n14501 6.541
R32420 S.n14513 S.t662 6.541
R32421 S.n14510 S.t2375 6.541
R32422 S.n14499 S.n14498 6.541
R32423 S.n14790 S.n14789 6.541
R32424 S.n14802 S.t327 6.541
R32425 S.n14805 S.t3182 6.541
R32426 S.n14787 S.n14786 6.541
R32427 S.n13543 S.n13542 6.541
R32428 S.n13554 S.t3753 6.541
R32429 S.n13551 S.t1305 6.541
R32430 S.n13540 S.n13539 6.541
R32431 S.n13820 S.n13819 6.541
R32432 S.n13832 S.t3810 6.541
R32433 S.n13835 S.t2138 6.541
R32434 S.n13817 S.n13816 6.541
R32435 S.n12571 S.n12570 6.541
R32436 S.n12582 S.t2667 6.541
R32437 S.n12579 S.t287 6.541
R32438 S.n12568 S.n12567 6.541
R32439 S.n12827 S.n12826 6.541
R32440 S.n12839 S.t2731 6.541
R32441 S.n12842 S.t1043 6.541
R32442 S.n12824 S.n12823 6.541
R32443 S.n11577 S.n11576 6.541
R32444 S.n11588 S.t1677 6.541
R32445 S.n11585 S.t3769 6.541
R32446 S.n11574 S.n11573 6.541
R32447 S.n11822 S.n11821 6.541
R32448 S.n11834 S.t1730 6.541
R32449 S.n11837 S.t4568 6.541
R32450 S.n11819 S.n11818 6.541
R32451 S.n10570 S.n10569 6.541
R32452 S.n10581 S.t630 6.541
R32453 S.n10578 S.t2682 6.541
R32454 S.n10567 S.n10566 6.541
R32455 S.n10794 S.n10793 6.541
R32456 S.n10806 S.t899 6.541
R32457 S.n10809 S.t3508 6.541
R32458 S.n10791 S.n10790 6.541
R32459 S.n9541 S.n9540 6.541
R32460 S.n9552 S.t4054 6.541
R32461 S.n9549 S.t3060 6.541
R32462 S.n9538 S.n9537 6.541
R32463 S.n9754 S.n9753 6.541
R32464 S.n9766 S.t3961 6.541
R32465 S.n9769 S.t4420 6.541
R32466 S.n9751 S.n9750 6.541
R32467 S.n8499 S.n8498 6.541
R32468 S.n8510 S.t2346 6.541
R32469 S.n8507 S.t1474 6.541
R32470 S.n8496 S.n8495 6.541
R32471 S.n8691 S.n8690 6.541
R32472 S.n8703 S.t3927 6.541
R32473 S.n8706 S.t4364 6.541
R32474 S.n8688 S.n8687 6.541
R32475 S.n7435 S.n7434 6.541
R32476 S.n7446 S.t2303 6.541
R32477 S.n7443 S.t1425 6.541
R32478 S.n7432 S.n7431 6.541
R32479 S.n7616 S.n7615 6.541
R32480 S.n7628 S.t3887 6.541
R32481 S.n7631 S.t4311 6.541
R32482 S.n7613 S.n7612 6.541
R32483 S.n6358 S.n6357 6.541
R32484 S.n6369 S.t2252 6.541
R32485 S.n6366 S.t1373 6.541
R32486 S.n6355 S.n6354 6.541
R32487 S.n6518 S.n6517 6.541
R32488 S.n6530 S.t3843 6.541
R32489 S.n6533 S.t4258 6.541
R32490 S.n6515 S.n6514 6.541
R32491 S.n5258 S.n5257 6.541
R32492 S.n5269 S.t2209 6.541
R32493 S.n5266 S.t1853 6.541
R32494 S.n5255 S.n5254 6.541
R32495 S.n5407 S.n5406 6.541
R32496 S.n5419 S.t4274 6.541
R32497 S.n5422 S.t464 6.541
R32498 S.n5404 S.n5403 6.541
R32499 S.n4145 S.n4144 6.541
R32500 S.n4156 S.t2868 6.541
R32501 S.n4153 S.t1807 6.541
R32502 S.n4142 S.n4141 6.541
R32503 S.n4273 S.n4272 6.541
R32504 S.n4285 S.t4222 6.541
R32505 S.n4288 S.t3404 6.541
R32506 S.n4270 S.n4269 6.541
R32507 S.n3019 S.n3018 6.541
R32508 S.n3030 S.t1278 6.541
R32509 S.n3027 S.t1763 6.541
R32510 S.n3016 S.n3015 6.541
R32511 S.n3137 S.n3136 6.541
R32512 S.n3148 S.t4172 6.541
R32513 S.n3151 S.t3363 6.541
R32514 S.n3134 S.n3133 6.541
R32515 S.n1858 S.n1857 6.541
R32516 S.n1870 S.t1227 6.541
R32517 S.n1867 S.t1718 6.541
R32518 S.n1855 S.n1854 6.541
R32519 S.n873 S.n872 6.541
R32520 S.n876 S.t1175 6.541
R32521 S.n879 S.t1676 6.541
R32522 S.n882 S.n881 6.541
R32523 S.n797 S.n796 6.541
R32524 S.n808 S.t1510 6.541
R32525 S.n811 S.t2766 6.541
R32526 S.n800 S.n799 6.541
R32527 S.n976 S.t2471 6.541
R32528 S.n978 S.t415 6.541
R32529 S.n22820 S.t258 6.541
R32530 S.n22818 S.t986 6.541
R32531 S.n22345 S.n22344 6.541
R32532 S.n22353 S.t3838 6.541
R32533 S.n22356 S.t3081 6.541
R32534 S.n22348 S.n22347 6.541
R32535 S.n22707 S.n22706 6.541
R32536 S.n22718 S.t1010 6.541
R32537 S.n22715 S.t4171 6.541
R32538 S.n22710 S.n22709 6.541
R32539 S.n21339 S.n21338 6.541
R32540 S.n21347 S.t279 6.541
R32541 S.n21350 S.t2378 6.541
R32542 S.n21342 S.n21341 6.541
R32543 S.n21255 S.n21254 6.541
R32544 S.n21263 S.t335 6.541
R32545 S.n21266 S.t3184 6.541
R32546 S.n21258 S.n21257 6.541
R32547 S.n20433 S.n20432 6.541
R32548 S.n20826 S.t3756 6.541
R32549 S.n20829 S.t1309 6.541
R32550 S.n20832 S.n20831 6.541
R32551 S.n20839 S.n20838 6.541
R32552 S.n20847 S.t4005 6.541
R32553 S.n20850 S.t2142 6.541
R32554 S.n20842 S.n20841 6.541
R32555 S.n19799 S.n19798 6.541
R32556 S.n20191 S.t2672 6.541
R32557 S.n20194 S.t513 6.541
R32558 S.n20197 S.n20196 6.541
R32559 S.n20204 S.n20203 6.541
R32560 S.n20215 S.t2999 6.541
R32561 S.n20212 S.t1048 6.541
R32562 S.n20207 S.n20206 6.541
R32563 S.n18927 S.n18926 6.541
R32564 S.n19321 S.t1681 6.541
R32565 S.n19324 S.t1890 6.541
R32566 S.n19327 S.n19326 6.541
R32567 S.n19334 S.n19333 6.541
R32568 S.n19345 S.t360 6.541
R32569 S.n19342 S.t2444 6.541
R32570 S.n19337 S.n19336 6.541
R32571 S.n18044 S.n18043 6.541
R32572 S.n18439 S.t3046 6.541
R32573 S.n18442 S.t1335 6.541
R32574 S.n18445 S.n18444 6.541
R32575 S.n18452 S.n18451 6.541
R32576 S.n18463 S.t3834 6.541
R32577 S.n18460 S.t1406 6.541
R32578 S.n18455 S.n18454 6.541
R32579 S.n17135 S.n17134 6.541
R32580 S.n17534 S.t1994 6.541
R32581 S.n17537 S.t310 6.541
R32582 S.n17540 S.n17539 6.541
R32583 S.n17547 S.n17546 6.541
R32584 S.n17558 S.t2763 6.541
R32585 S.n17555 S.t371 6.541
R32586 S.n17550 S.n17549 6.541
R32587 S.n16217 S.n16216 6.541
R32588 S.n16616 S.t938 6.541
R32589 S.n16619 S.t3788 6.541
R32590 S.n16622 S.n16621 6.541
R32591 S.n16629 S.n16628 6.541
R32592 S.n16640 S.t1757 6.541
R32593 S.n16637 S.t4039 6.541
R32594 S.n16632 S.n16631 6.541
R32595 S.n15273 S.n15272 6.541
R32596 S.n15676 S.t107 6.541
R32597 S.n15679 S.t2708 6.541
R32598 S.n15682 S.n15681 6.541
R32599 S.n15689 S.n15688 6.541
R32600 S.n15700 S.t711 6.541
R32601 S.n15697 S.t3039 6.541
R32602 S.n15692 S.n15691 6.541
R32603 S.n14320 S.n14319 6.541
R32604 S.n14723 S.t3618 6.541
R32605 S.n14726 S.t821 6.541
R32606 S.n14729 S.n14728 6.541
R32607 S.n14736 S.n14735 6.541
R32608 S.n14747 S.t3299 6.541
R32609 S.n14744 S.t1631 6.541
R32610 S.n14739 S.n14738 6.541
R32611 S.n13341 S.n13340 6.541
R32612 S.n13748 S.t2211 6.541
R32613 S.n13751 S.t4253 6.541
R32614 S.n13754 S.n13753 6.541
R32615 S.n13761 S.n13760 6.541
R32616 S.n13772 S.t2267 6.541
R32617 S.n13769 S.t573 6.541
R32618 S.n13764 S.n13763 6.541
R32619 S.n12353 S.n12352 6.541
R32620 S.n12760 S.t1109 6.541
R32621 S.n12763 S.t3257 6.541
R32622 S.n12766 S.n12765 6.541
R32623 S.n12773 S.n12772 6.541
R32624 S.n12784 S.t1171 6.541
R32625 S.n12781 S.t4013 6.541
R32626 S.n12776 S.n12775 6.541
R32627 S.n11339 S.n11338 6.541
R32628 S.n11750 S.t55 6.541
R32629 S.n11753 S.t2225 6.541
R32630 S.n11756 S.n11755 6.541
R32631 S.n11763 S.n11762 6.541
R32632 S.n11774 S.t390 6.541
R32633 S.n11771 S.t3010 6.541
R32634 S.n11766 S.n11765 6.541
R32635 S.n10316 S.n10315 6.541
R32636 S.n10727 S.t3580 6.541
R32637 S.n10730 S.t1561 6.541
R32638 S.n10733 S.n10732 6.541
R32639 S.n10740 S.n10739 6.541
R32640 S.n10751 S.t3980 6.541
R32641 S.n10748 S.t2918 6.541
R32642 S.n10743 S.n10742 6.541
R32643 S.n9267 S.n9266 6.541
R32644 S.n9682 S.t824 6.541
R32645 S.n9685 S.t1511 6.541
R32646 S.n9688 S.n9687 6.541
R32647 S.n9695 S.n9694 6.541
R32648 S.n9706 S.t2421 6.541
R32649 S.n9703 S.t2865 6.541
R32650 S.n9698 S.n9697 6.541
R32651 S.n8209 S.n8208 6.541
R32652 S.n8624 S.t790 6.541
R32653 S.n8627 S.t4425 6.541
R32654 S.n8630 S.n8629 6.541
R32655 S.n8637 S.n8636 6.541
R32656 S.n8648 S.t2386 6.541
R32657 S.n8645 S.t2811 6.541
R32658 S.n8640 S.n8639 6.541
R32659 S.n7125 S.n7124 6.541
R32660 S.n7544 S.t738 6.541
R32661 S.n7547 S.t4371 6.541
R32662 S.n7550 S.n7549 6.541
R32663 S.n7557 S.n7556 6.541
R32664 S.n7568 S.t2351 6.541
R32665 S.n7565 S.t2753 6.541
R32666 S.n7560 S.n7559 6.541
R32667 S.n6032 S.n6031 6.541
R32668 S.n6451 S.t689 6.541
R32669 S.n6454 S.t4320 6.541
R32670 S.n6457 S.n6456 6.541
R32671 S.n6464 S.n6463 6.541
R32672 S.n6475 S.t2305 6.541
R32673 S.n6472 S.t2969 6.541
R32674 S.n6467 S.n6466 6.541
R32675 S.n4912 S.n4911 6.541
R32676 S.n5335 S.t865 6.541
R32677 S.n5338 S.t292 6.541
R32678 S.n5341 S.n5340 6.541
R32679 S.n5348 S.n5347 6.541
R32680 S.n5359 S.t2720 6.541
R32681 S.n5356 S.t3425 6.541
R32682 S.n5351 S.n5350 6.541
R32683 S.n3784 S.n3783 6.541
R32684 S.n4206 S.t1300 6.541
R32685 S.n4209 S.t241 6.541
R32686 S.n4212 S.n4211 6.541
R32687 S.n4219 S.n4218 6.541
R32688 S.n4230 S.t2670 6.541
R32689 S.n4227 S.t1858 6.541
R32690 S.n4222 S.n4221 6.541
R32691 S.n2637 S.n2636 6.541
R32692 S.n3065 S.t4228 6.541
R32693 S.n3068 S.t194 6.541
R32694 S.n3071 S.n3070 6.541
R32695 S.n3078 S.n3077 6.541
R32696 S.n3089 S.t2623 6.541
R32697 S.n3086 S.t1816 6.541
R32698 S.n3081 S.n3080 6.541
R32699 S.n1876 S.n1875 6.541
R32700 S.n1884 S.t4178 6.541
R32701 S.n1887 S.t129 6.541
R32702 S.n1879 S.n1878 6.541
R32703 S.n1921 S.n1920 6.541
R32704 S.n1936 S.t2583 6.541
R32705 S.n1933 S.t2580 6.541
R32706 S.n1924 S.n1923 6.541
R32707 S.n1294 S.t4150 6.541
R32708 S.n400 S.n399 6.541
R32709 S.n411 S.t2849 6.541
R32710 S.n408 S.t1788 6.541
R32711 S.n403 S.n402 6.541
R32712 S.n2129 S.n2128 6.541
R32713 S.n2139 S.t2904 6.541
R32714 S.n2142 S.t1839 6.541
R32715 S.n2126 S.n2125 6.541
R32716 S.n18063 S.t3519 6.541
R32717 S.n18471 S.n18470 6.541
R32718 S.n18488 S.t1495 6.541
R32719 S.n18485 S.t3815 6.541
R32720 S.n18468 S.n18467 6.541
R32721 S.n17163 S.n17162 6.541
R32722 S.n17174 S.t4370 6.541
R32723 S.n17171 S.t2466 6.541
R32724 S.n17160 S.n17159 6.541
R32725 S.n17755 S.n17754 6.541
R32726 S.n17767 S.t445 6.541
R32727 S.n17770 S.t2737 6.541
R32728 S.n17752 S.n17751 6.541
R32729 S.n16263 S.n16262 6.541
R32730 S.n16274 S.t3346 6.541
R32731 S.n16271 S.t1438 6.541
R32732 S.n16260 S.n16259 6.541
R32733 S.n16828 S.n16827 6.541
R32734 S.n16840 S.t3906 6.541
R32735 S.n16843 S.t1738 6.541
R32736 S.n16825 S.n16824 6.541
R32737 S.n15339 S.n15338 6.541
R32738 S.n15350 S.t2322 6.541
R32739 S.n15347 S.t399 6.541
R32740 S.n15336 S.n15335 6.541
R32741 S.n15893 S.n15892 6.541
R32742 S.n15905 S.t3117 6.541
R32743 S.n15908 S.t696 6.541
R32744 S.n15890 S.n15889 6.541
R32745 S.n14402 S.n14401 6.541
R32746 S.n14413 S.t1232 6.541
R32747 S.n14410 S.t3224 6.541
R32748 S.n14399 S.n14398 6.541
R32749 S.n14935 S.n14934 6.541
R32750 S.n14947 S.t1134 6.541
R32751 S.n14950 S.t3787 6.541
R32752 S.n14932 S.n14931 6.541
R32753 S.n13443 S.n13442 6.541
R32754 S.n13454 S.t4338 6.541
R32755 S.n13451 S.t4594 6.541
R32756 S.n13440 S.n13439 6.541
R32757 S.n13965 S.n13964 6.541
R32758 S.n13977 S.t2520 6.541
R32759 S.n13980 S.t651 6.541
R32760 S.n13962 S.n13961 6.541
R32761 S.n12471 S.n12470 6.541
R32762 S.n12482 S.t1180 6.541
R32763 S.n12479 S.t3534 6.541
R32764 S.n12468 S.n12467 6.541
R32765 S.n12972 S.n12971 6.541
R32766 S.n12984 S.t1516 6.541
R32767 S.n12987 S.t4071 6.541
R32768 S.n12969 S.n12968 6.541
R32769 S.n11477 S.n11476 6.541
R32770 S.n11488 S.t162 6.541
R32771 S.n11485 S.t2480 6.541
R32772 S.n11474 S.n11473 6.541
R32773 S.n11967 S.n11966 6.541
R32774 S.n11979 S.t460 6.541
R32775 S.n11982 S.t3080 6.541
R32776 S.n11964 S.n11963 6.541
R32777 S.n10470 S.n10469 6.541
R32778 S.n10481 S.t3657 6.541
R32779 S.n10478 S.t1454 6.541
R32780 S.n10467 S.n10466 6.541
R32781 S.n10939 S.n10938 6.541
R32782 S.n10951 S.t3923 6.541
R32783 S.n10954 S.t2268 6.541
R32784 S.n10936 S.n10935 6.541
R32785 S.n9441 S.n9440 6.541
R32786 S.n9452 S.t2809 6.541
R32787 S.n9449 S.t413 6.541
R32788 S.n9438 S.n9437 6.541
R32789 S.n9899 S.n9898 6.541
R32790 S.n9911 S.t3399 6.541
R32791 S.n9914 S.t1176 6.541
R32792 S.n9896 S.n9895 6.541
R32793 S.n8399 S.n8398 6.541
R32794 S.n8410 S.t1798 6.541
R32795 S.n8407 S.t4380 6.541
R32796 S.n8396 S.n8395 6.541
R32797 S.n8836 S.n8835 6.541
R32798 S.n8848 S.t2371 6.541
R32799 S.n8851 S.t154 6.541
R32800 S.n8833 S.n8832 6.541
R32801 S.n7335 S.n7334 6.541
R32802 S.n7346 S.t759 6.541
R32803 S.n7343 S.t3354 6.541
R32804 S.n7332 S.n7331 6.541
R32805 S.n7761 S.n7760 6.541
R32806 S.n7773 S.t1293 6.541
R32807 S.n7776 S.t3648 6.541
R32808 S.n7758 S.n7757 6.541
R32809 S.n6258 S.n6257 6.541
R32810 S.n6269 S.t4180 6.541
R32811 S.n6266 S.t2328 6.541
R32812 S.n6255 S.n6254 6.541
R32813 S.n6663 S.n6662 6.541
R32814 S.n6675 S.t280 6.541
R32815 S.n6678 S.t2567 6.541
R32816 S.n6660 S.n6659 6.541
R32817 S.n5158 S.n5157 6.541
R32818 S.n5169 S.t3196 6.541
R32819 S.n5166 S.t3855 6.541
R32820 S.n5155 S.n5154 6.541
R32821 S.n5553 S.n5552 6.541
R32822 S.n5565 S.t2047 6.541
R32823 S.n5568 S.t4097 6.541
R32824 S.n5550 S.n5549 6.541
R32825 S.n4046 S.n4045 6.541
R32826 S.n4057 S.t197 6.541
R32827 S.n4054 S.t535 6.541
R32828 S.n4043 S.n4042 6.541
R32829 S.n4418 S.n4417 6.541
R32830 S.n4430 S.t3005 6.541
R32831 S.n4433 S.t1921 6.541
R32832 S.n4415 S.n4414 6.541
R32833 S.n2919 S.n2918 6.541
R32834 S.n2930 S.t4304 6.541
R32835 S.n2927 S.t489 6.541
R32836 S.n2916 S.n2915 6.541
R32837 S.n3281 S.n3280 6.541
R32838 S.n3292 S.t2955 6.541
R32839 S.n3295 S.t1877 6.541
R32840 S.n3278 S.n3277 6.541
R32841 S.n1750 S.n1749 6.541
R32842 S.n1762 S.t4247 6.541
R32843 S.n1759 S.t446 6.541
R32844 S.n1747 S.n1746 6.541
R32845 S.n1416 S.t2851 6.541
R32846 S.n12 S.n11 6.541
R32847 S.n15 S.t1281 6.541
R32848 S.n18 S.t452 6.541
R32849 S.n21 S.n20 6.541
R32850 S.n18947 S.t2483 6.541
R32851 S.n19357 S.n19356 6.541
R32852 S.n19375 S.t956 6.541
R32853 S.n19372 S.t3305 6.541
R32854 S.n19360 S.n19359 6.541
R32855 S.n18071 S.n18070 6.541
R32856 S.n18082 S.t3876 6.541
R32857 S.n18079 S.t1970 6.541
R32858 S.n18074 S.n18073 6.541
R32859 S.n18618 S.n18617 6.541
R32860 S.n18635 S.t4445 6.541
R32861 S.n18638 S.t2274 6.541
R32862 S.n18621 S.n18620 6.541
R32863 S.n17182 S.n17181 6.541
R32864 S.n17193 S.t2817 6.541
R32865 S.n17190 S.t921 6.541
R32866 S.n17185 S.n17184 6.541
R32867 S.n17718 S.n17717 6.541
R32868 S.n17735 S.t3401 6.541
R32869 S.n17738 S.t1178 6.541
R32870 S.n17721 S.n17720 6.541
R32871 S.n16280 S.n16279 6.541
R32872 S.n16291 S.t1800 6.541
R32873 S.n16288 S.t4386 6.541
R32874 S.n16283 S.n16282 6.541
R32875 S.n16791 S.n16790 6.541
R32876 S.n16808 S.t2559 6.541
R32877 S.n16811 S.t166 6.541
R32878 S.n16794 S.n16793 6.541
R32879 S.n15356 S.n15355 6.541
R32880 S.n15367 S.t765 6.541
R32881 S.n15364 S.t3590 6.541
R32882 S.n15359 S.n15358 6.541
R32883 S.n15856 S.n15855 6.541
R32884 S.n15873 S.t1565 6.541
R32885 S.n15876 S.t3653 6.541
R32886 S.n15859 S.n15858 6.541
R32887 S.n14419 S.n14418 6.541
R32888 S.n14430 S.t4185 6.541
R32889 S.n14427 S.t4040 6.541
R32890 S.n14422 S.n14421 6.541
R32891 S.n14898 S.n14897 6.541
R32892 S.n14915 S.t2039 6.541
R32893 S.n14918 S.t98 6.541
R32894 S.n14901 S.n14900 6.541
R32895 S.n13460 S.n13459 6.541
R32896 S.n13471 S.t713 6.541
R32897 S.n13468 S.t3034 6.541
R32898 S.n13463 S.n13462 6.541
R32899 S.n13928 S.n13927 6.541
R32900 S.n13945 S.t972 6.541
R32901 S.n13948 S.t3605 6.541
R32902 S.n13931 S.n13930 6.541
R32903 S.n12488 S.n12487 6.541
R32904 S.n12499 S.t4135 6.541
R32905 S.n12496 S.t1984 6.541
R32906 S.n12491 S.n12490 6.541
R32907 S.n12935 S.n12934 6.541
R32908 S.n12952 S.t4460 6.541
R32909 S.n12955 S.t2531 6.541
R32910 S.n12938 S.n12937 6.541
R32911 S.n11494 S.n11493 6.541
R32912 S.n11505 S.t3152 6.541
R32913 S.n11502 S.t930 6.541
R32914 S.n11497 S.n11496 6.541
R32915 S.n11930 S.n11929 6.541
R32916 S.n11947 S.t3419 6.541
R32917 S.n11950 S.t1748 6.541
R32918 S.n11933 S.n11932 6.541
R32919 S.n10487 S.n10486 6.541
R32920 S.n10498 S.t2333 6.541
R32921 S.n10495 S.t4403 6.541
R32922 S.n10490 S.n10489 6.541
R32923 S.n10902 S.n10901 6.541
R32924 S.n10919 S.t2382 6.541
R32925 S.n10922 S.t707 6.541
R32926 S.n10905 S.n10904 6.541
R32927 S.n9458 S.n9457 6.541
R32928 S.n9469 S.t1247 6.541
R32929 S.n9466 S.t3376 6.541
R32930 S.n9461 S.n9460 6.541
R32931 S.n9862 S.n9861 6.541
R32932 S.n9879 S.t1856 6.541
R32933 S.n9882 S.t4130 6.541
R32934 S.n9865 S.n9864 6.541
R32935 S.n8416 S.n8415 6.541
R32936 S.n8427 S.t233 6.541
R32937 S.n8424 S.t2828 6.541
R32938 S.n8419 S.n8418 6.541
R32939 S.n8799 S.n8798 6.541
R32940 S.n8816 S.t815 6.541
R32941 S.n8819 S.t3146 6.541
R32942 S.n8802 S.n8801 6.541
R32943 S.n7352 S.n7351 6.541
R32944 S.n7363 S.t3714 6.541
R32945 S.n7360 S.t1809 6.541
R32946 S.n7355 S.n7354 6.541
R32947 S.n7724 S.n7723 6.541
R32948 S.n7741 S.t4242 6.541
R32949 S.n7744 S.t2097 6.541
R32950 S.n7727 S.n7726 6.541
R32951 S.n6275 S.n6274 6.541
R32952 S.n6286 S.t2630 6.541
R32953 S.n6283 S.t773 6.541
R32954 S.n6278 S.n6277 6.541
R32955 S.n6626 S.n6625 6.541
R32956 S.n6643 S.t3457 6.541
R32957 S.n6646 S.t1018 6.541
R32958 S.n6629 S.n6628 6.541
R32959 S.n5175 S.n5174 6.541
R32960 S.n5186 S.t1643 6.541
R32961 S.n5183 S.t3542 6.541
R32962 S.n5178 S.n5177 6.541
R32963 S.n5516 S.n5515 6.541
R32964 S.n5533 S.t1500 6.541
R32965 S.n5536 S.t1940 6.541
R32966 S.n5519 S.n5518 6.541
R32967 S.n4063 S.n4062 6.541
R32968 S.n4074 S.t4330 6.541
R32969 S.n4071 S.t3491 6.541
R32970 S.n4066 S.n4065 6.541
R32971 S.n4381 S.n4380 6.541
R32972 S.n4398 S.t1447 6.541
R32973 S.n4401 S.t364 6.541
R32974 S.n4384 S.n4383 6.541
R32975 S.n2936 S.n2935 6.541
R32976 S.n2947 S.t2745 6.541
R32977 S.n2944 S.t3447 6.541
R32978 S.n2939 S.n2938 6.541
R32979 S.n3244 S.n3243 6.541
R32980 S.n3261 S.t1392 6.541
R32981 S.n3264 S.t315 6.541
R32982 S.n3247 S.n3246 6.541
R32983 S.n1768 S.n1767 6.541
R32984 S.n1781 S.t2697 6.541
R32985 S.n1778 S.t3403 6.541
R32986 S.n1771 S.n1770 6.541
R32987 S.n1790 S.n1789 6.541
R32988 S.n1804 S.t1138 6.541
R32989 S.n1801 S.t1861 6.541
R32990 S.n1793 S.n1792 6.541
R32991 S.n2060 S.n2059 6.541
R32992 S.n2081 S.t4284 6.541
R32993 S.n2084 S.t3451 6.541
R32994 S.n2063 S.n2062 6.541
R32995 S.n415 S.n414 6.541
R32996 S.n814 S.t1344 6.541
R32997 S.n817 S.t1820 6.541
R32998 S.n820 S.n819 6.541
R32999 S.n828 S.n827 6.541
R33000 S.n843 S.t4232 6.541
R33001 S.n840 S.t3407 6.541
R33002 S.n831 S.n830 6.541
R33003 S.n1308 S.t1287 6.541
R33004 S.n3221 S.n3220 6.541
R33005 S.n3232 S.t4340 6.541
R33006 S.n3235 S.t3285 6.541
R33007 S.n3218 S.n3217 6.541
R33008 S.n4357 S.n4356 6.541
R33009 S.n4369 S.t4394 6.541
R33010 S.n4372 S.t3330 6.541
R33011 S.n4354 S.n4353 6.541
R33012 S.n5492 S.n5491 6.541
R33013 S.n5504 S.t4449 6.541
R33014 S.n5507 S.t381 6.541
R33015 S.n5489 S.n5488 6.541
R33016 S.n6602 S.n6601 6.541
R33017 S.n6614 S.t3965 6.541
R33018 S.n6617 S.t4436 6.541
R33019 S.n6599 S.n6598 6.541
R33020 S.n7700 S.n7699 6.541
R33021 S.n7712 S.t2951 6.541
R33022 S.n7715 S.t530 6.541
R33023 S.n7697 S.n7696 6.541
R33024 S.n8775 S.n8774 6.541
R33025 S.n8787 S.t3776 6.541
R33026 S.n8790 S.t1590 6.541
R33027 S.n8772 S.n8771 6.541
R33028 S.n9838 S.n9837 6.541
R33029 S.n9850 S.t296 6.541
R33030 S.n9853 S.t2586 6.541
R33031 S.n9835 S.n9834 6.541
R33032 S.n10878 S.n10877 6.541
R33033 S.n10890 S.t827 6.541
R33034 S.n10893 S.t3665 6.541
R33035 S.n10875 S.n10874 6.541
R33036 S.n11906 S.n11905 6.541
R33037 S.n11918 S.t1874 6.541
R33038 S.n11921 S.t179 6.541
R33039 S.n11903 S.n11902 6.541
R33040 S.n12911 S.n12910 6.541
R33041 S.n12923 S.t2907 6.541
R33042 S.n12926 S.t1193 6.541
R33043 S.n12908 S.n12907 6.541
R33044 S.n13904 S.n13903 6.541
R33045 S.n13916 S.t3938 6.541
R33046 S.n13919 S.t2050 6.541
R33047 S.n13901 S.n13900 6.541
R33048 S.n14874 S.n14873 6.541
R33049 S.n14886 S.t477 6.541
R33050 S.n14889 S.t3103 6.541
R33051 S.n14871 S.n14870 6.541
R33052 S.n15832 S.n15831 6.541
R33053 S.n15844 S.t2408 6.541
R33054 S.n15847 S.t4510 6.541
R33055 S.n15829 S.n15828 6.541
R33056 S.n16767 S.n16766 6.541
R33057 S.n16779 S.t1012 6.541
R33058 S.n16782 S.t3154 6.541
R33059 S.n16764 S.n16763 6.541
R33060 S.n17690 S.n17689 6.541
R33061 S.n17702 S.t2089 6.541
R33062 S.n17705 S.t4133 6.541
R33063 S.n17687 S.n17686 6.541
R33064 S.n18590 S.n18589 6.541
R33065 S.n18602 S.t2888 6.541
R33066 S.n18605 S.t709 6.541
R33067 S.n18587 S.n18586 6.541
R33068 S.n19480 S.n19479 6.541
R33069 S.n19492 S.t3925 6.541
R33070 S.n19495 S.t1755 6.541
R33071 S.n19477 S.n19476 6.541
R33072 S.n20226 S.n20225 6.541
R33073 S.n20243 S.t4466 6.541
R33074 S.n20240 S.t2754 6.541
R33075 S.n20223 S.n20222 6.541
R33076 S.n19818 S.t1990 6.541
R33077 S.n18955 S.n18954 6.541
R33078 S.n18966 S.t3368 6.541
R33079 S.n18963 S.t935 6.541
R33080 S.n18952 S.n18951 6.541
R33081 S.n18090 S.n18089 6.541
R33082 S.n18101 S.t2341 6.541
R33083 S.n18098 S.t414 6.541
R33084 S.n18087 S.n18086 6.541
R33085 S.n17201 S.n17200 6.541
R33086 S.n17212 S.t1252 6.541
R33087 S.n17209 S.t3886 6.541
R33088 S.n17198 S.n17197 6.541
R33089 S.n16299 S.n16298 6.541
R33090 S.n16310 S.t238 6.541
R33091 S.n16307 S.t3085 6.541
R33092 S.n16296 S.n16295 6.541
R33093 S.n15375 S.n15374 6.541
R33094 S.n15386 S.t3721 6.541
R33095 S.n15383 S.t4441 6.541
R33096 S.n15372 S.n15371 6.541
R33097 S.n14438 S.n14437 6.541
R33098 S.n14449 S.t571 6.541
R33099 S.n14446 S.t2495 6.541
R33100 S.n14435 S.n14434 6.541
R33101 S.n13479 S.n13478 6.541
R33102 S.n13490 S.t3671 6.541
R33103 S.n13487 S.t1476 6.541
R33104 S.n13476 S.n13475 6.541
R33105 S.n12507 S.n12506 6.541
R33106 S.n12518 S.t2589 6.541
R33107 S.n12515 S.t429 6.541
R33108 S.n12504 S.n12503 6.541
R33109 S.n11513 S.n11512 6.541
R33110 S.n11524 S.t1818 6.541
R33111 S.n11521 S.t3898 6.541
R33112 S.n11510 S.n11509 6.541
R33113 S.n10506 S.n10505 6.541
R33114 S.n10517 S.t780 6.541
R33115 S.n10514 S.t2850 6.541
R33116 S.n10503 S.n10502 6.541
R33117 S.n9477 S.n9476 6.541
R33118 S.n9488 S.t4201 6.541
R33119 S.n9485 S.t1831 6.541
R33120 S.n9474 S.n9473 6.541
R33121 S.n8435 S.n8434 6.541
R33122 S.n8446 S.t3209 6.541
R33123 S.n8443 S.t1260 6.541
R33124 S.n8432 S.n8431 6.541
R33125 S.n7371 S.n7370 6.541
R33126 S.n7382 S.t2171 6.541
R33127 S.n7379 S.t243 6.541
R33128 S.n7368 S.n7367 6.541
R33129 S.n6294 S.n6293 6.541
R33130 S.n6305 S.t1074 6.541
R33131 S.n6302 S.t1543 6.541
R33132 S.n6291 S.n6290 6.541
R33133 S.n5194 S.n5193 6.541
R33134 S.n5205 S.t2354 6.541
R33135 S.n5202 S.t1992 6.541
R33136 S.n5191 S.n5190 6.541
R33137 S.n4082 S.n4081 6.541
R33138 S.n4093 S.t2772 6.541
R33139 S.n4090 S.t1943 6.541
R33140 S.n4079 S.n4078 6.541
R33141 S.n2955 S.n2954 6.541
R33142 S.n2966 S.t1186 6.541
R33143 S.n2963 S.t1904 6.541
R33144 S.n2952 S.n2951 6.541
R33145 S.n2032 S.n2031 6.541
R33146 S.n2047 S.t2727 6.541
R33147 S.n2050 S.t1907 6.541
R33148 S.n2035 S.n2034 6.541
R33149 S.n753 S.n752 6.541
R33150 S.n772 S.t4293 6.541
R33151 S.n769 S.t252 6.541
R33152 S.n756 S.n755 6.541
R33153 S.n1324 S.n1323 6.541
R33154 S.n1327 S.t2679 6.541
R33155 S.n1330 S.t1868 6.541
R33156 S.n1333 S.n1332 6.541
R33157 S.n1319 S.t4237 6.541
R33158 S.n20455 S.t1485 6.541
R33159 S.n20418 S.n20417 6.541
R33160 S.n20426 S.t3942 6.541
R33161 S.n20429 S.t2292 6.541
R33162 S.n20415 S.n20414 6.541
R33163 S.n19835 S.n19834 6.541
R33164 S.n19844 S.t2839 6.541
R33165 S.n19841 S.t433 6.541
R33166 S.n19832 S.n19831 6.541
R33167 S.n20314 S.n20313 6.541
R33168 S.n20332 S.t2911 6.541
R33169 S.n20335 S.t1198 6.541
R33170 S.n20311 S.n20310 6.541
R33171 S.n18983 S.n18982 6.541
R33172 S.n18992 S.t1823 6.541
R33173 S.n18989 S.t3902 6.541
R33174 S.n18980 S.n18979 6.541
R33175 S.n19442 S.n19441 6.541
R33176 S.n19460 S.t2387 6.541
R33177 S.n19463 S.t184 6.541
R33178 S.n19439 S.n19438 6.541
R33179 S.n18118 S.n18117 6.541
R33180 S.n18126 S.t786 6.541
R33181 S.n18123 S.t3379 6.541
R33182 S.n18115 S.n18114 6.541
R33183 S.n18555 S.n18554 6.541
R33184 S.n18570 S.t1583 6.541
R33185 S.n18573 S.t3667 6.541
R33186 S.n18552 S.n18551 6.541
R33187 S.n17229 S.n17228 6.541
R33188 S.n17237 S.t4205 6.541
R33189 S.n17234 S.t2535 6.541
R33190 S.n17226 S.n17225 6.541
R33191 S.n17655 S.n17654 6.541
R33192 S.n17670 S.t523 6.541
R33193 S.n17673 S.t2591 6.541
R33194 S.n17652 S.n17651 6.541
R33195 S.n16327 S.n16326 6.541
R33196 S.n16335 S.t3216 6.541
R33197 S.n16332 S.t3918 6.541
R33198 S.n16324 S.n16323 6.541
R33199 S.n16732 S.n16731 6.541
R33200 S.n16747 S.t1899 6.541
R33201 S.n16750 S.t3970 6.541
R33202 S.n16729 S.n16728 6.541
R33203 S.n15403 S.n15402 6.541
R33204 S.n15411 S.t4579 6.541
R33205 S.n15408 S.t2883 6.541
R33206 S.n15400 S.n15399 6.541
R33207 S.n15797 S.n15796 6.541
R33208 S.n15812 S.t857 6.541
R33209 S.n15815 S.t2952 6.541
R33210 S.n15794 S.n15793 6.541
R33211 S.n14466 S.n14465 6.541
R33212 S.n14474 S.t3521 6.541
R33213 S.n14471 S.t944 6.541
R33214 S.n14463 S.n14462 6.541
R33215 S.n14839 S.n14838 6.541
R33216 S.n14854 S.t3436 6.541
R33217 S.n14857 S.t1550 6.541
R33218 S.n14836 S.n14835 6.541
R33219 S.n13507 S.n13506 6.541
R33220 S.n13515 S.t2125 6.541
R33221 S.n13512 S.t4424 6.541
R33222 S.n13504 S.n13503 6.541
R33223 S.n13869 S.n13868 6.541
R33224 S.n13884 S.t2400 6.541
R33225 S.n13887 S.t728 6.541
R33226 S.n13866 S.n13865 6.541
R33227 S.n12535 S.n12534 6.541
R33228 S.n12543 S.t1267 6.541
R33229 S.n12540 S.t3390 6.541
R33230 S.n12532 S.n12531 6.541
R33231 S.n12876 S.n12875 6.541
R33232 S.n12891 S.t1341 6.541
R33233 S.n12894 S.t4148 6.541
R33234 S.n12873 S.n12872 6.541
R33235 S.n11541 S.n11540 6.541
R33236 S.n11549 S.t250 6.541
R33237 S.n11546 S.t2363 6.541
R33238 S.n11538 S.n11537 6.541
R33239 S.n11871 S.n11870 6.541
R33240 S.n11886 S.t311 6.541
R33241 S.n11889 S.t3163 6.541
R33242 S.n11868 S.n11867 6.541
R33243 S.n10534 S.n10533 6.541
R33244 S.n10542 S.t3736 6.541
R33245 S.n10539 S.t1284 6.541
R33246 S.n10531 S.n10530 6.541
R33247 S.n10843 S.n10842 6.541
R33248 S.n10858 S.t3791 6.541
R33249 S.n10861 S.t2117 6.541
R33250 S.n10840 S.n10839 6.541
R33251 S.n9505 S.n9504 6.541
R33252 S.n9513 S.t2651 6.541
R33253 S.n9510 S.t267 6.541
R33254 S.n9502 S.n9501 6.541
R33255 S.n9803 S.n9802 6.541
R33256 S.n9818 S.t3267 6.541
R33257 S.n9821 S.t1033 6.541
R33258 S.n9800 S.n9799 6.541
R33259 S.n8463 S.n8462 6.541
R33260 S.n8471 S.t1660 6.541
R33261 S.n8468 S.t4212 6.541
R33262 S.n8460 S.n8459 6.541
R33263 S.n8740 S.n8739 6.541
R33264 S.n8755 S.t2431 6.541
R33265 S.n8758 S.t4547 6.541
R33266 S.n8737 S.n8736 6.541
R33267 S.n7399 S.n7398 6.541
R33268 S.n7407 S.t607 6.541
R33269 S.n7404 S.t4545 6.541
R33270 S.n7396 S.n7395 6.541
R33271 S.n7665 S.n7664 6.541
R33272 S.n7680 S.t2468 6.541
R33273 S.n7683 S.t2930 6.541
R33274 S.n7662 S.n7661 6.541
R33275 S.n6322 S.n6321 6.541
R33276 S.n6330 S.t833 6.541
R33277 S.n6327 S.t4489 6.541
R33278 S.n6319 S.n6318 6.541
R33279 S.n6567 S.n6566 6.541
R33280 S.n6582 S.t2427 6.541
R33281 S.n6585 S.t2877 6.541
R33282 S.n6564 S.n6563 6.541
R33283 S.n5222 S.n5221 6.541
R33284 S.n5230 S.t797 6.541
R33285 S.n5227 S.t434 6.541
R33286 S.n5219 S.n5218 6.541
R33287 S.n5457 S.n5456 6.541
R33288 S.n5472 S.t2890 6.541
R33289 S.n5475 S.t3348 6.541
R33290 S.n5454 S.n5453 6.541
R33291 S.n4110 S.n4109 6.541
R33292 S.n4118 S.t1211 6.541
R33293 S.n4115 S.t387 6.541
R33294 S.n4107 S.n4106 6.541
R33295 S.n4322 S.n4321 6.541
R33296 S.n4337 S.t2840 6.541
R33297 S.n4340 S.t1781 6.541
R33298 S.n4319 S.n4318 6.541
R33299 S.n2983 S.n2982 6.541
R33300 S.n2991 S.t4141 6.541
R33301 S.n2988 S.t346 6.541
R33302 S.n2980 S.n2979 6.541
R33303 S.n3185 S.n3184 6.541
R33304 S.n3200 S.t2782 6.541
R33305 S.n3203 S.t1953 6.541
R33306 S.n3182 S.n3181 6.541
R33307 S.n1820 S.n1819 6.541
R33308 S.n1828 S.t4344 6.541
R33309 S.n1825 S.t301 6.541
R33310 S.n1817 S.n1816 6.541
R33311 S.n1999 S.n1998 6.541
R33312 S.n2014 S.t1168 6.541
R33313 S.n2017 S.t352 6.541
R33314 S.n2002 S.n2001 6.541
R33315 S.n777 S.n776 6.541
R33316 S.n791 S.t2735 6.541
R33317 S.n788 S.t3230 6.541
R33318 S.n780 S.n779 6.541
R33319 S.n1841 S.n1840 6.541
R33320 S.n1850 S.t2787 6.541
R33321 S.n1847 S.t3271 6.541
R33322 S.n1838 S.n1837 6.541
R33323 S.n3160 S.n3159 6.541
R33324 S.n3168 S.t1222 6.541
R33325 S.n3171 S.t402 6.541
R33326 S.n3163 S.n3162 6.541
R33327 S.n2997 S.n2996 6.541
R33328 S.n3011 S.t2846 6.541
R33329 S.n3008 S.t3313 6.541
R33330 S.n3000 S.n2999 6.541
R33331 S.n4297 S.n4296 6.541
R33332 S.n4305 S.t1272 6.541
R33333 S.n4308 S.t442 6.541
R33334 S.n4300 S.n4299 6.541
R33335 S.n4124 S.n4123 6.541
R33336 S.n4137 S.t4164 6.541
R33337 S.n4134 S.t3353 6.541
R33338 S.n4127 S.n4126 6.541
R33339 S.n5431 S.n5430 6.541
R33340 S.n5440 S.t1325 6.541
R33341 S.n5443 S.t1803 6.541
R33342 S.n5434 S.n5433 6.541
R33343 S.n5236 S.n5235 6.541
R33344 S.n5250 S.t3749 6.541
R33345 S.n5247 S.t3397 6.541
R33346 S.n5239 S.n5238 6.541
R33347 S.n6542 S.n6541 6.541
R33348 S.n6550 S.t880 6.541
R33349 S.n6553 S.t1310 6.541
R33350 S.n6545 S.n6544 6.541
R33351 S.n6336 S.n6335 6.541
R33352 S.n6350 S.t3794 6.541
R33353 S.n6347 S.t2933 6.541
R33354 S.n6339 S.n6338 6.541
R33355 S.n7640 S.n7639 6.541
R33356 S.n7648 S.t922 6.541
R33357 S.n7651 S.t1362 6.541
R33358 S.n7643 S.n7642 6.541
R33359 S.n7413 S.n7412 6.541
R33360 S.n7427 S.t3840 6.541
R33361 S.n7424 S.t2985 6.541
R33362 S.n7416 S.n7415 6.541
R33363 S.n8715 S.n8714 6.541
R33364 S.n8723 S.t959 6.541
R33365 S.n8726 S.t1421 6.541
R33366 S.n8718 S.n8717 6.541
R33367 S.n8477 S.n8476 6.541
R33368 S.n8491 S.t20 6.541
R33369 S.n8488 S.t3033 6.541
R33370 S.n8480 S.n8479 6.541
R33371 S.n9778 S.n9777 6.541
R33372 S.n9786 S.t1931 6.541
R33373 S.n9789 S.t3998 6.541
R33374 S.n9781 S.n9780 6.541
R33375 S.n9519 S.n9518 6.541
R33376 S.n9533 S.t1090 6.541
R33377 S.n9530 S.t3242 6.541
R33378 S.n9522 S.n9521 6.541
R33379 S.n10818 S.n10817 6.541
R33380 S.n10826 S.t2248 6.541
R33381 S.n10829 S.t552 6.541
R33382 S.n10821 S.n10820 6.541
R33383 S.n10548 S.n10547 6.541
R33384 S.n10562 S.t2189 6.541
R33385 S.n10559 S.t4234 6.541
R33386 S.n10551 S.n10550 6.541
R33387 S.n11846 S.n11845 6.541
R33388 S.n11854 S.t3280 6.541
R33389 S.n11857 S.t1608 6.541
R33390 S.n11849 S.n11848 6.541
R33391 S.n11555 S.n11554 6.541
R33392 S.n11569 S.t3228 6.541
R33393 S.n11566 S.t809 6.541
R33394 S.n11558 S.n11557 6.541
R33395 S.n12851 S.n12850 6.541
R33396 S.n12859 S.t4290 6.541
R33397 S.n12862 S.t2598 6.541
R33398 S.n12854 S.n12853 6.541
R33399 S.n12549 S.n12548 6.541
R33400 S.n12563 S.t4218 6.541
R33401 S.n12560 S.t1847 6.541
R33402 S.n12552 S.n12551 6.541
R33403 S.n13844 S.n13843 6.541
R33404 S.n13852 S.t849 6.541
R33405 S.n13855 S.t3684 6.541
R33406 S.n13847 S.n13846 6.541
R33407 S.n13521 S.n13520 6.541
R33408 S.n13535 S.t799 6.541
R33409 S.n13532 S.t2872 6.541
R33410 S.n13524 S.n13523 6.541
R33411 S.n14814 S.n14813 6.541
R33412 S.n14822 S.t1889 6.541
R33413 S.n14825 S.t203 6.541
R33414 S.n14817 S.n14816 6.541
R33415 S.n14480 S.n14479 6.541
R33416 S.n14494 S.t1973 6.541
R33417 S.n14491 S.t3908 6.541
R33418 S.n14483 S.n14482 6.541
R33419 S.n15772 S.n15771 6.541
R33420 S.n15780 S.t3817 6.541
R33421 S.n15783 S.t1386 6.541
R33422 S.n15775 S.n15774 6.541
R33423 S.n15417 S.n15416 6.541
R33424 S.n15431 S.t3024 6.541
R33425 S.n15428 S.t1315 6.541
R33426 S.n15420 S.n15419 6.541
R33427 S.n16707 S.n16706 6.541
R33428 S.n16715 S.t341 6.541
R33429 S.n16718 S.t2432 6.541
R33430 S.n16710 S.n16709 6.541
R33431 S.n16341 S.n16340 6.541
R33432 S.n16355 S.t4026 6.541
R33433 S.n16352 S.t2381 6.541
R33434 S.n16344 S.n16343 6.541
R33435 S.n17630 S.n17629 6.541
R33436 S.n17638 S.t1370 6.541
R33437 S.n17641 S.t3475 6.541
R33438 S.n17633 S.n17632 6.541
R33439 S.n17243 S.n17242 6.541
R33440 S.n17257 S.t2659 6.541
R33441 S.n17254 S.t3415 6.541
R33442 S.n17246 S.n17245 6.541
R33443 S.n18530 S.n18529 6.541
R33444 S.n18538 S.t4540 6.541
R33445 S.n18541 S.t2121 6.541
R33446 S.n18533 S.n18532 6.541
R33447 S.n18132 S.n18131 6.541
R33448 S.n18146 S.t3740 6.541
R33449 S.n18143 S.t2055 6.541
R33450 S.n18135 S.n18134 6.541
R33451 S.n19417 S.n19416 6.541
R33452 S.n19425 S.t1027 6.541
R33453 S.n19428 S.t3167 6.541
R33454 S.n19420 S.n19419 6.541
R33455 S.n18998 S.n18997 6.541
R33456 S.n19012 S.t255 6.541
R33457 S.n19009 S.t2368 6.541
R33458 S.n19001 S.n19000 6.541
R33459 S.n20289 S.n20288 6.541
R33460 S.n20297 S.t1346 6.541
R33461 S.n20300 S.t4152 6.541
R33462 S.n20292 S.n20291 6.541
R33463 S.n19852 S.n19851 6.541
R33464 S.n19866 S.t1271 6.541
R33465 S.n19863 S.t3393 6.541
R33466 S.n19855 S.n19854 6.541
R33467 S.n20360 S.n20359 6.541
R33468 S.n20371 S.t2403 6.541
R33469 S.n20368 S.t730 6.541
R33470 S.n20363 S.n20362 6.541
R33471 S.n20463 S.n20462 6.541
R33472 S.n20477 S.t2357 6.541
R33473 S.n20474 S.t4433 6.541
R33474 S.n20466 S.n20465 6.541
R33475 S.n21236 S.n21235 6.541
R33476 S.n21244 S.t3440 6.541
R33477 S.n21247 S.t1771 6.541
R33478 S.n21239 S.n21238 6.541
R33479 S.n21300 S.t951 6.541
R33480 S.n1367 S.t2686 6.541
R33481 S.n852 S.n851 6.541
R33482 S.n869 S.t1122 6.541
R33483 S.n866 S.t306 6.541
R33484 S.n855 S.n854 6.541
R33485 S.n2093 S.n2092 6.541
R33486 S.n2109 S.t1336 6.541
R33487 S.n2112 S.t276 6.541
R33488 S.n2096 S.n2095 6.541
R33489 S.n737 S.n736 6.541
R33490 S.n748 S.t2653 6.541
R33491 S.n745 S.t3365 6.541
R33492 S.n740 S.n739 6.541
R33493 S.n720 S.n719 6.541
R33494 S.n731 S.t4203 6.541
R33495 S.n728 S.t401 6.541
R33496 S.n723 S.n722 6.541
R33497 S.n1282 S.t2755 6.541
R33498 S.n368 S.n367 6.541
R33499 S.n379 S.t1452 6.541
R33500 S.n376 S.t370 6.541
R33501 S.n371 S.n370 6.541
R33502 S.n2188 S.n2187 6.541
R33503 S.n2198 S.t1513 6.541
R33504 S.n2201 S.t419 6.541
R33505 S.n2185 S.n2184 6.541
R33506 S.n16236 S.t4558 6.541
R33507 S.n16648 S.n16647 6.541
R33508 S.n16665 S.t2491 6.541
R33509 S.n16662 S.t314 6.541
R33510 S.n16645 S.n16644 6.541
R33511 S.n15301 S.n15300 6.541
R33512 S.n15312 S.t894 6.541
R33513 S.n15309 S.t3499 6.541
R33514 S.n15298 S.n15297 6.541
R33515 S.n15958 S.n15957 6.541
R33516 S.n15970 S.t1470 6.541
R33517 S.n15973 S.t3799 6.541
R33518 S.n15955 S.n15954 6.541
R33519 S.n14366 S.n14365 6.541
R33520 S.n14377 S.t4350 6.541
R33521 S.n14374 S.t1593 6.541
R33522 S.n14363 S.n14362 6.541
R33523 S.n14996 S.n14995 6.541
R33524 S.n15008 S.t4025 6.541
R33525 S.n15011 S.t2380 6.541
R33526 S.n14993 S.n14992 6.541
R33527 S.n13407 S.n13406 6.541
R33528 S.n13418 S.t2958 6.541
R33529 S.n13415 S.t532 6.541
R33530 S.n13404 S.n13403 6.541
R33531 S.n14026 S.n14025 6.541
R33532 S.n14038 S.t3255 6.541
R33533 S.n14041 S.t1313 6.541
R33534 S.n14023 S.n14022 6.541
R33535 S.n12435 S.n12434 6.541
R33536 S.n12446 S.t1915 6.541
R33537 S.n12443 S.t4199 6.541
R33538 S.n12432 S.n12431 6.541
R33539 S.n13033 S.n13032 6.541
R33540 S.n13045 S.t2220 6.541
R33541 S.n13048 S.t294 6.541
R33542 S.n13030 S.n13029 6.541
R33543 S.n11441 S.n11440 6.541
R33544 S.n11452 S.t873 6.541
R33545 S.n11449 S.t1052 6.541
R33546 S.n11438 S.n11437 6.541
R33547 S.n12028 S.n12027 6.541
R33548 S.n12040 S.t3570 6.541
R33549 S.n12043 S.t1678 6.541
R33550 S.n12025 S.n12024 6.541
R33551 S.n10434 S.n10433 6.541
R33552 S.n10445 S.t2254 6.541
R33553 S.n10442 S.t4575 6.541
R33554 S.n10431 S.n10430 6.541
R33555 S.n11000 S.n10999 6.541
R33556 S.n11012 S.t2505 6.541
R33557 S.n11015 S.t634 6.541
R33558 S.n10997 S.n10996 6.541
R33559 S.n9405 S.n9404 6.541
R33560 S.n9416 S.t1160 6.541
R33561 S.n9413 S.t3517 6.541
R33562 S.n9402 S.n9401 6.541
R33563 S.n9960 S.n9959 6.541
R33564 S.n9972 S.t1998 6.541
R33565 S.n9975 S.t4058 6.541
R33566 S.n9957 S.n9956 6.541
R33567 S.n8363 S.n8362 6.541
R33568 S.n8374 S.t133 6.541
R33569 S.n8371 S.t2993 6.541
R33570 S.n8360 S.n8359 6.541
R33571 S.n8897 S.n8896 6.541
R33572 S.n8909 S.t937 6.541
R33573 S.n8912 S.t3282 6.541
R33574 S.n8894 S.n8893 6.541
R33575 S.n7299 S.n7298 6.541
R33576 S.n7310 S.t3856 6.541
R33577 S.n7307 S.t1949 6.541
R33578 S.n7296 S.n7295 6.541
R33579 S.n7822 S.n7821 6.541
R33580 S.n7834 S.t4414 6.541
R33581 S.n7837 S.t2249 6.541
R33582 S.n7819 S.n7818 6.541
R33583 S.n6222 S.n6221 6.541
R33584 S.n6233 S.t2788 6.541
R33585 S.n6230 S.t902 6.541
R33586 S.n6219 S.n6218 6.541
R33587 S.n6724 S.n6723 6.541
R33588 S.n6736 S.t3386 6.541
R33589 S.n6739 S.t1156 6.541
R33590 S.n6721 S.n6720 6.541
R33591 S.n5122 S.n5121 6.541
R33592 S.n5133 S.t1780 6.541
R33593 S.n5130 S.t2438 6.541
R33594 S.n5119 S.n5118 6.541
R33595 S.n5614 S.n5613 6.541
R33596 S.n5626 S.t410 6.541
R33597 S.n5629 S.t2704 6.541
R33598 S.n5611 S.n5610 6.541
R33599 S.n4010 S.n4009 6.541
R33600 S.n4021 S.t3318 6.541
R33601 S.n4018 S.t1397 6.541
R33602 S.n4007 S.n4006 6.541
R33603 S.n4479 S.n4478 6.541
R33604 S.n4491 S.t3881 6.541
R33605 S.n4494 S.t2223 6.541
R33606 S.n4476 S.n4475 6.541
R33607 S.n2883 S.n2882 6.541
R33608 S.n2894 S.t2748 6.541
R33609 S.n2891 S.t361 6.541
R33610 S.n2880 S.n2879 6.541
R33611 S.n3341 S.n3340 6.541
R33612 S.n3352 S.t3078 6.541
R33613 S.n3355 S.t1124 6.541
R33614 S.n3338 S.n3337 6.541
R33615 S.n1713 S.n1712 6.541
R33616 S.n1725 S.t1744 6.541
R33617 S.n1722 S.t3553 6.541
R33618 S.n1710 S.n1709 6.541
R33619 S.n1412 S.t1196 6.541
R33620 S.n59 S.n58 6.541
R33621 S.n62 S.t4402 6.541
R33622 S.n65 S.t3335 6.541
R33623 S.n68 S.n67 6.541
R33624 S.n17155 S.t4007 6.541
R33625 S.n17570 S.n17569 6.541
R33626 S.n17588 S.t2000 6.541
R33627 S.n17585 S.t4296 6.541
R33628 S.n17573 S.n17572 6.541
R33629 S.n16244 S.n16243 6.541
R33630 S.n16255 S.t379 6.541
R33631 S.n16252 S.t3000 6.541
R33632 S.n16247 S.n16246 6.541
R33633 S.n16856 S.n16855 6.541
R33634 S.n16873 S.t942 6.541
R33635 S.n16876 S.t3284 6.541
R33636 S.n16859 S.n16858 6.541
R33637 S.n15320 S.n15319 6.541
R33638 S.n15331 S.t3858 6.541
R33639 S.n15328 S.t1951 6.541
R33640 S.n15323 S.n15322 6.541
R33641 S.n15921 S.n15920 6.541
R33642 S.n15938 S.t4417 6.541
R33643 S.n15941 S.t2256 6.541
R33644 S.n15924 S.n15923 6.541
R33645 S.n14383 S.n14382 6.541
R33646 S.n14394 S.t2792 6.541
R33647 S.n14391 S.t4549 6.541
R33648 S.n14386 S.n14385 6.541
R33649 S.n14959 S.n14958 6.541
R33650 S.n14976 S.t2694 6.541
R33651 S.n14979 S.t825 6.541
R33652 S.n14962 S.n14961 6.541
R33653 S.n13424 S.n13423 6.541
R33654 S.n13435 S.t1390 6.541
R33655 S.n13432 S.t3729 6.541
R33656 S.n13427 S.n13426 6.541
R33657 S.n13989 S.n13988 6.541
R33658 S.n14006 S.t1701 6.541
R33659 S.n14009 S.t4260 6.541
R33660 S.n13992 S.n13991 6.541
R33661 S.n12452 S.n12451 6.541
R33662 S.n12463 S.t358 6.541
R33663 S.n12460 S.t582 6.541
R33664 S.n12455 S.n12454 6.541
R33665 S.n12996 S.n12995 6.541
R33666 S.n13013 S.t3066 6.541
R33667 S.n13016 S.t1111 6.541
R33668 S.n12999 S.n12998 6.541
R33669 S.n11458 S.n11457 6.541
R33670 S.n11469 S.t1736 6.541
R33671 S.n11466 S.t4019 6.541
R33672 S.n11461 S.n11460 6.541
R33673 S.n11991 S.n11990 6.541
R33674 S.n12008 S.t2020 6.541
R33675 S.n12011 S.t57 6.541
R33676 S.n11994 S.n11993 6.541
R33677 S.n10451 S.n10450 6.541
R33678 S.n10462 S.t699 6.541
R33679 S.n10459 S.t3016 6.541
R33680 S.n10454 S.n10453 6.541
R33681 S.n10963 S.n10962 6.541
R33682 S.n10980 S.t954 6.541
R33683 S.n10983 S.t3585 6.541
R33684 S.n10966 S.n10965 6.541
R33685 S.n9422 S.n9421 6.541
R33686 S.n9433 S.t4114 6.541
R33687 S.n9430 S.t1967 6.541
R33688 S.n9425 S.n9424 6.541
R33689 S.n9923 S.n9922 6.541
R33690 S.n9940 S.t441 6.541
R33691 S.n9943 S.t2736 6.541
R33692 S.n9926 S.n9925 6.541
R33693 S.n8380 S.n8379 6.541
R33694 S.n8391 S.t3344 6.541
R33695 S.n8388 S.t1435 6.541
R33696 S.n8383 S.n8382 6.541
R33697 S.n8860 S.n8859 6.541
R33698 S.n8877 S.t3903 6.541
R33699 S.n8880 S.t1731 6.541
R33700 S.n8863 S.n8862 6.541
R33701 S.n7316 S.n7315 6.541
R33702 S.n7327 S.t2319 6.541
R33703 S.n7324 S.t391 6.541
R33704 S.n7319 S.n7318 6.541
R33705 S.n7785 S.n7784 6.541
R33706 S.n7802 S.t2861 6.541
R33707 S.n7805 S.t688 6.541
R33708 S.n7788 S.n7787 6.541
R33709 S.n6239 S.n6238 6.541
R33710 S.n6250 S.t1228 6.541
R33711 S.n6247 S.t3865 6.541
R33712 S.n6242 S.n6241 6.541
R33713 S.n6687 S.n6686 6.541
R33714 S.n6704 S.t1841 6.541
R33715 S.n6707 S.t4109 6.541
R33716 S.n6690 S.n6689 6.541
R33717 S.n5139 S.n5138 6.541
R33718 S.n5150 S.t215 6.541
R33719 S.n5147 S.t892 6.541
R33720 S.n5142 S.n5141 6.541
R33721 S.n5577 S.n5576 6.541
R33722 S.n5594 S.t3373 6.541
R33723 S.n5597 S.t1144 6.541
R33724 S.n5580 S.n5579 6.541
R33725 S.n4027 S.n4026 6.541
R33726 S.n4038 S.t1767 6.541
R33727 S.n4035 S.t4346 6.541
R33728 S.n4030 S.n4029 6.541
R33729 S.n4442 S.n4441 6.541
R33730 S.n4459 S.t2530 6.541
R33731 S.n4462 S.t665 6.541
R33732 S.n4445 S.n4444 6.541
R33733 S.n2900 S.n2899 6.541
R33734 S.n2911 S.t1189 6.541
R33735 S.n2908 S.t2053 6.541
R33736 S.n2903 S.n2902 6.541
R33737 S.n3304 S.n3303 6.541
R33738 S.n3321 S.t4512 6.541
R33739 S.n3324 S.t3423 6.541
R33740 S.n3307 S.n3306 6.541
R33741 S.n1731 S.n1730 6.541
R33742 S.n1742 S.t1297 6.541
R33743 S.n1739 S.t2003 6.541
R33744 S.n1734 S.n1733 6.541
R33745 S.n2151 S.n2150 6.541
R33746 S.n2168 S.t4458 6.541
R33747 S.n2171 S.t3382 6.541
R33748 S.n2154 S.n2153 6.541
R33749 S.n702 S.n701 6.541
R33750 S.n713 S.t1248 6.541
R33751 S.n710 S.t1955 6.541
R33752 S.n705 S.n704 6.541
R33753 S.n685 S.n684 6.541
R33754 S.n696 S.t2815 6.541
R33755 S.n693 S.t3502 6.541
R33756 S.n688 S.n687 6.541
R33757 S.n1269 S.t2729 6.541
R33758 S.n336 S.n335 6.541
R33759 S.n347 S.t4055 6.541
R33760 S.n344 S.t2205 6.541
R33761 S.n339 S.n338 6.541
R33762 S.n2247 S.n2246 6.541
R33763 S.n2257 S.t385 6.541
R33764 S.n2260 S.t3239 6.541
R33765 S.n2244 S.n2243 6.541
R33766 S.n14339 S.t156 6.541
R33767 S.n14755 S.n14754 6.541
R33768 S.n14772 S.t2613 6.541
R33769 S.n14769 S.t950 6.541
R33770 S.n14752 S.n14751 6.541
R33771 S.n13369 S.n13368 6.541
R33772 S.n13380 S.t1566 6.541
R33773 S.n13377 S.t3650 6.541
R33774 S.n13366 S.n13365 6.541
R33775 S.n14091 S.n14090 6.541
R33776 S.n14103 S.t1623 6.541
R33777 S.n14106 S.t4438 6.541
R33778 S.n14088 S.n14087 6.541
R33779 S.n12399 S.n12398 6.541
R33780 S.n12410 S.t502 6.541
R33781 S.n12407 S.t2570 6.541
R33782 S.n12396 S.n12395 6.541
R33783 S.n13094 S.n13093 6.541
R33784 S.n13106 S.t568 6.541
R33785 S.n13109 S.t3395 6.541
R33786 S.n13091 S.n13090 6.541
R33787 S.n11405 S.n11404 6.541
R33788 S.n11416 S.t3956 6.541
R33789 S.n11413 S.t1579 6.541
R33790 S.n11402 S.n11401 6.541
R33791 S.n12089 S.n12088 6.541
R33792 S.n12101 S.t4229 6.541
R33793 S.n12104 S.t2370 6.541
R33794 S.n12086 S.n12085 6.541
R33795 S.n10398 S.n10397 6.541
R33796 S.n10409 S.t2936 6.541
R33797 S.n10406 S.t756 6.541
R33798 S.n10395 S.n10394 6.541
R33799 S.n11061 S.n11060 6.541
R33800 S.n11073 S.t3237 6.541
R33801 S.n11076 S.t1291 6.541
R33802 S.n11058 S.n11057 6.541
R33803 S.n9369 S.n9368 6.541
R33804 S.n9380 S.t1900 6.541
R33805 S.n9377 S.t2131 6.541
R33806 S.n9366 S.n9365 6.541
R33807 S.n10021 S.n10020 6.541
R33808 S.n10033 S.t593 6.541
R33809 S.n10036 S.t2656 6.541
R33810 S.n10018 S.n10017 6.541
R33811 S.n8327 S.n8326 6.541
R33812 S.n8338 S.t3273 6.541
R33813 S.n8335 S.t1599 6.541
R33814 S.n8324 S.n8323 6.541
R33815 S.n8958 S.n8957 6.541
R33816 S.n8970 S.t4028 6.541
R33817 S.n8973 S.t1663 6.541
R33818 S.n8955 S.n8954 6.541
R33819 S.n7263 S.n7262 6.541
R33820 S.n7274 S.t2237 6.541
R33821 S.n7271 S.t537 6.541
R33822 S.n7260 S.n7259 6.541
R33823 S.n7883 S.n7882 6.541
R33824 S.n7895 S.t3023 6.541
R33825 S.n7898 S.t609 6.541
R33826 S.n7880 S.n7879 6.541
R33827 S.n6186 S.n6185 6.541
R33828 S.n6197 S.t1145 6.541
R33829 S.n6194 S.t3990 6.541
R33830 S.n6183 S.n6182 6.541
R33831 S.n6785 S.n6784 6.541
R33832 S.n6797 S.t1978 6.541
R33833 S.n6800 S.t4266 6.541
R33834 S.n6782 S.n6781 6.541
R33835 S.n5086 S.n5085 6.541
R33836 S.n5097 S.t362 6.541
R33837 S.n5094 S.t1014 6.541
R33838 S.n5083 S.n5082 6.541
R33839 S.n5675 S.n5674 6.541
R33840 S.n5687 S.t3513 6.541
R33841 S.n5690 S.t1306 6.541
R33842 S.n5672 S.n5671 6.541
R33843 S.n3974 S.n3973 6.541
R33844 S.n3985 S.t1909 6.541
R33845 S.n3982 S.t4523 6.541
R33846 S.n3971 S.n3970 6.541
R33847 S.n4540 S.n4539 6.541
R33848 S.n4552 S.t2462 6.541
R33849 S.n4555 S.t807 6.541
R33850 S.n4537 S.n4536 6.541
R33851 S.n2847 S.n2846 6.541
R33852 S.n2858 S.t1358 6.541
R33853 S.n2855 S.t3468 6.541
R33854 S.n2844 S.n2843 6.541
R33855 S.n3401 S.n3400 6.541
R33856 S.n3412 S.t1431 6.541
R33857 S.n3415 S.t4231 6.541
R33858 S.n3398 S.n3397 6.541
R33859 S.n1676 S.n1675 6.541
R33860 S.n1688 S.t326 6.541
R33861 S.n1685 S.t2422 6.541
R33862 S.n1673 S.n1672 6.541
R33863 S.n1408 S.t4314 6.541
R33864 S.n91 S.n90 6.541
R33865 S.n94 S.t3015 6.541
R33866 S.n97 S.t1930 6.541
R33867 S.n100 S.n99 6.541
R33868 S.n15293 S.t541 6.541
R33869 S.n15712 S.n15711 6.541
R33870 S.n15730 S.t3027 6.541
R33871 S.n15727 S.t835 6.541
R33872 S.n15715 S.n15714 6.541
R33873 S.n14347 S.n14346 6.541
R33874 S.n14358 S.t1400 6.541
R33875 S.n14355 S.t3148 6.541
R33876 S.n14350 S.n14349 6.541
R33877 S.n15024 S.n15023 6.541
R33878 S.n15041 S.t1056 6.541
R33879 S.n15044 S.t3920 6.541
R33880 S.n15027 S.n15026 6.541
R33881 S.n13388 S.n13387 6.541
R33882 S.n13399 S.t4516 6.541
R33883 S.n13396 S.t2101 6.541
R33884 S.n13391 S.n13390 6.541
R33885 S.n14054 S.n14053 6.541
R33886 S.n14071 S.t4580 6.541
R33887 S.n14074 S.t2881 6.541
R33888 S.n14057 S.n14056 6.541
R33889 S.n12416 S.n12415 6.541
R33890 S.n12427 S.t3462 6.541
R33891 S.n12424 S.t1021 6.541
R33892 S.n12419 S.n12418 6.541
R33893 S.n13057 S.n13056 6.541
R33894 S.n13074 S.t3759 6.541
R33895 S.n13077 S.t1850 6.541
R33896 S.n13060 S.n13059 6.541
R33897 S.n11422 S.n11421 6.541
R33898 S.n11433 S.t2418 6.541
R33899 S.n11430 S.t230 6.541
R33900 S.n11425 S.n11424 6.541
R33901 S.n12052 S.n12051 6.541
R33902 S.n12069 S.t2677 6.541
R33903 S.n12072 S.t814 6.541
R33904 S.n12055 S.n12054 6.541
R33905 S.n10415 S.n10414 6.541
R33906 S.n10426 S.t1371 6.541
R33907 S.n10423 S.t1619 6.541
R33908 S.n10418 S.n10417 6.541
R33909 S.n11024 S.n11023 6.541
R33910 S.n11041 S.t4047 6.541
R33911 S.n11044 S.t2191 6.541
R33912 S.n11027 S.n11026 6.541
R33913 S.n9386 S.n9385 6.541
R33914 S.n9397 S.t2721 6.541
R33915 S.n9394 S.t564 6.541
R33916 S.n9389 S.n9388 6.541
R33917 S.n9984 S.n9983 6.541
R33918 S.n10001 S.t3547 6.541
R33919 S.n10004 S.t1094 6.541
R33920 S.n9987 S.n9986 6.541
R33921 S.n8344 S.n8343 6.541
R33922 S.n8355 S.t1721 6.541
R33923 S.n8352 S.t4555 6.541
R33924 S.n8347 S.n8346 6.541
R33925 S.n8921 S.n8920 6.541
R33926 S.n8938 S.t2487 6.541
R33927 S.n8941 S.t24 6.541
R33928 S.n8924 S.n8923 6.541
R33929 S.n7280 S.n7279 6.541
R33930 S.n7291 S.t676 6.541
R33931 S.n7288 S.t3497 6.541
R33932 S.n7283 S.n7282 6.541
R33933 S.n7846 S.n7845 6.541
R33934 S.n7863 S.t1467 6.541
R33935 S.n7866 S.t3792 6.541
R33936 S.n7849 S.n7848 6.541
R33937 S.n6203 S.n6202 6.541
R33938 S.n6214 S.t4347 6.541
R33939 S.n6211 S.t2449 6.541
R33940 S.n6206 S.n6205 6.541
R33941 S.n6748 S.n6747 6.541
R33942 S.n6765 S.t422 6.541
R33943 S.n6768 S.t2712 6.541
R33944 S.n6751 S.n6750 6.541
R33945 S.n5103 S.n5102 6.541
R33946 S.n5114 S.t3328 6.541
R33947 S.n5111 S.t3978 6.541
R33948 S.n5106 S.n5105 6.541
R33949 S.n5638 S.n5637 6.541
R33950 S.n5655 S.t1964 6.541
R33951 S.n5658 S.t4254 6.541
R33952 S.n5641 S.n5640 6.541
R33953 S.n3991 S.n3990 6.541
R33954 S.n4002 S.t349 6.541
R33955 S.n3999 S.t2964 6.541
R33956 S.n3994 S.n3993 6.541
R33957 S.n4503 S.n4502 6.541
R33958 S.n4520 S.t918 6.541
R33959 S.n4523 S.t3766 6.541
R33960 S.n4506 S.n4505 6.541
R33961 S.n2864 S.n2863 6.541
R33962 S.n2875 S.t4307 6.541
R33963 S.n2872 S.t1920 6.541
R33964 S.n2867 S.n2866 6.541
R33965 S.n3364 S.n3363 6.541
R33966 S.n3381 S.t4377 6.541
R33967 S.n3384 S.t2680 6.541
R33968 S.n3367 S.n3366 6.541
R33969 S.n1694 S.n1693 6.541
R33970 S.n1705 S.t3294 6.541
R33971 S.n1702 S.t877 6.541
R33972 S.n1697 S.n1696 6.541
R33973 S.n2210 S.n2209 6.541
R33974 S.n2227 S.t3581 6.541
R33975 S.n2230 S.t1688 6.541
R33976 S.n2213 S.n2212 6.541
R33977 S.n667 S.n666 6.541
R33978 S.n678 S.t2265 6.541
R33979 S.n675 S.t547 6.541
R33980 S.n670 S.n669 6.541
R33981 S.n650 S.n649 6.541
R33982 S.n661 S.t3807 6.541
R33983 S.n658 S.t1377 6.541
R33984 S.n653 S.n652 6.541
R33985 S.n1256 S.t1338 6.541
R33986 S.n304 S.n303 6.541
R33987 S.n315 S.t2447 6.541
R33988 S.n312 S.t792 6.541
R33989 S.n307 S.n306 6.541
R33990 S.n2306 S.n2305 6.541
R33991 S.n2316 S.t3493 6.541
R33992 S.n2319 S.t1827 6.541
R33993 S.n2303 S.n2302 6.541
R33994 S.n12372 S.t1157 6.541
R33995 S.n12792 S.n12791 6.541
R33996 S.n12809 S.t3682 6.541
R33997 S.n12806 S.t1995 6.541
R33998 S.n12789 S.n12788 6.541
R33999 S.n11367 S.n11366 6.541
R34000 S.n11378 S.t2540 6.541
R34001 S.n11375 S.t132 6.541
R34002 S.n11364 S.n11363 6.541
R34003 S.n12154 S.n12153 6.541
R34004 S.n12166 S.t2596 6.541
R34005 S.n12169 S.t936 6.541
R34006 S.n12151 S.n12150 6.541
R34007 S.n10362 S.n10361 6.541
R34008 S.n10373 S.t1540 6.541
R34009 S.n10370 S.t3635 6.541
R34010 S.n10359 S.n10358 6.541
R34011 S.n11122 S.n11121 6.541
R34012 S.n11134 S.t1602 6.541
R34013 S.n11137 S.t4411 6.541
R34014 S.n11119 S.n11118 6.541
R34015 S.n9333 S.n9332 6.541
R34016 S.n9344 S.t483 6.541
R34017 S.n9341 S.t2555 6.541
R34018 S.n9330 S.n9329 6.541
R34019 S.n10082 S.n10081 6.541
R34020 S.n10094 S.t1255 6.541
R34021 S.n10097 S.t3385 6.541
R34022 S.n10079 S.n10078 6.541
R34023 S.n8291 S.n8290 6.541
R34024 S.n8302 S.t3944 6.541
R34025 S.n8299 S.t2298 6.541
R34026 S.n8288 S.n8287 6.541
R34027 S.n9019 S.n9018 6.541
R34028 S.n9031 S.t237 6.541
R34029 S.n9034 S.t2355 6.541
R34030 S.n9016 S.n9015 6.541
R34031 S.n7227 S.n7226 6.541
R34032 S.n7238 S.t2913 6.541
R34033 S.n7235 S.t3659 6.541
R34034 S.n7224 S.n7223 6.541
R34035 S.n7944 S.n7943 6.541
R34036 S.n7956 S.t1629 6.541
R34037 S.n7959 S.t3717 6.541
R34038 S.n7941 S.n7940 6.541
R34039 S.n6150 S.n6149 6.541
R34040 S.n6161 S.t4251 6.541
R34041 S.n6158 S.t2573 6.541
R34042 S.n6147 S.n6146 6.541
R34043 S.n6846 S.n6845 6.541
R34044 S.n6858 S.t574 6.541
R34045 S.n6861 S.t2631 6.541
R34046 S.n6843 S.n6842 6.541
R34047 S.n5050 S.n5049 6.541
R34048 S.n5061 S.t3258 6.541
R34049 S.n5058 S.t4104 6.541
R34050 S.n5047 S.n5046 6.541
R34051 S.n5736 S.n5735 6.541
R34052 S.n5748 S.t2126 6.541
R34053 S.n5751 S.t4168 6.541
R34054 S.n5733 S.n5732 6.541
R34055 S.n3938 S.n3937 6.541
R34056 S.n3949 S.t273 6.541
R34057 S.n3946 S.t3120 6.541
R34058 S.n3935 S.n3934 6.541
R34059 S.n4601 S.n4600 6.541
R34060 S.n4613 S.t1038 6.541
R34061 S.n4616 S.t3897 6.541
R34062 S.n4598 S.n4597 6.541
R34063 S.n2811 S.n2810 6.541
R34064 S.n2822 S.t4479 6.541
R34065 S.n2819 S.t2073 6.541
R34066 S.n2808 S.n2807 6.541
R34067 S.n3461 S.n3460 6.541
R34068 S.n3472 S.t4554 6.541
R34069 S.n3475 S.t2848 6.541
R34070 S.n3458 S.n3457 6.541
R34071 S.n1639 S.n1638 6.541
R34072 S.n1651 S.t3434 6.541
R34073 S.n1648 S.t998 6.541
R34074 S.n1636 S.n1635 6.541
R34075 S.n1404 S.t4287 6.541
R34076 S.n123 S.n122 6.541
R34077 S.n981 S.t900 6.541
R34078 S.n984 S.t3744 6.541
R34079 S.n987 S.n986 6.541
R34080 S.n13361 S.t693 6.541
R34081 S.n13784 S.n13783 6.541
R34082 S.n13802 S.t3177 6.541
R34083 S.n13799 S.t1489 6.541
R34084 S.n13787 S.n13786 6.541
R34085 S.n12380 S.n12379 6.541
R34086 S.n12391 S.t2067 6.541
R34087 S.n12388 S.t4113 6.541
R34088 S.n12383 S.n12382 6.541
R34089 S.n13122 S.n13121 6.541
R34090 S.n13139 S.t2134 6.541
R34091 S.n13142 S.t439 6.541
R34092 S.n13125 S.n13124 6.541
R34093 S.n11386 S.n11385 6.541
R34094 S.n11397 S.t993 6.541
R34095 S.n11394 S.t3134 6.541
R34096 S.n11389 S.n11388 6.541
R34097 S.n12117 S.n12116 6.541
R34098 S.n12134 S.t1042 6.541
R34099 S.n12137 S.t3901 6.541
R34100 S.n12120 S.n12119 6.541
R34101 S.n10379 S.n10378 6.541
R34102 S.n10390 S.t4493 6.541
R34103 S.n10387 S.t2082 6.541
R34104 S.n10382 S.n10381 6.541
R34105 S.n11085 S.n11084 6.541
R34106 S.n11102 S.t259 6.541
R34107 S.n11105 S.t2859 6.541
R34108 S.n11088 S.n11087 6.541
R34109 S.n9350 S.n9349 6.541
R34110 S.n9361 S.t3444 6.541
R34111 S.n9358 S.t1224 6.541
R34112 S.n9353 S.n9352 6.541
R34113 S.n10045 S.n10044 6.541
R34114 S.n10062 S.t4207 6.541
R34115 S.n10065 S.t1838 6.541
R34116 S.n10048 S.n10047 6.541
R34117 S.n8308 S.n8307 6.541
R34118 S.n8319 S.t2406 6.541
R34119 S.n8316 S.t3156 6.541
R34120 S.n8311 S.n8310 6.541
R34121 S.n8982 S.n8981 6.541
R34122 S.n8999 S.t1061 6.541
R34123 S.n9002 S.t3212 6.541
R34124 S.n8985 S.n8984 6.541
R34125 S.n7244 S.n7243 6.541
R34126 S.n7255 S.t3781 6.541
R34127 S.n7252 S.t2105 6.541
R34128 S.n7247 S.n7246 6.541
R34129 S.n7907 S.n7906 6.541
R34130 S.n7924 S.t4583 6.541
R34131 S.n7927 S.t2172 6.541
R34132 S.n7910 S.n7909 6.541
R34133 S.n6167 S.n6166 6.541
R34134 S.n6178 S.t2700 6.541
R34135 S.n6175 S.t1026 6.541
R34136 S.n6170 S.n6169 6.541
R34137 S.n6809 S.n6808 6.541
R34138 S.n6826 S.t3526 6.541
R34139 S.n6829 S.t1078 6.541
R34140 S.n6812 S.n6811 6.541
R34141 S.n5067 S.n5066 6.541
R34142 S.n5078 S.t1703 6.541
R34143 S.n5075 S.t2561 6.541
R34144 S.n5070 S.n5069 6.541
R34145 S.n5699 S.n5698 6.541
R34146 S.n5716 S.t558 6.541
R34147 S.n5719 S.t2869 6.541
R34148 S.n5702 S.n5701 6.541
R34149 S.n3955 S.n3954 6.541
R34150 S.n3966 S.t3453 6.541
R34151 S.n3963 S.t1570 6.541
R34152 S.n3958 S.n3957 6.541
R34153 S.n4564 S.n4563 6.541
R34154 S.n4581 S.t4003 6.541
R34155 S.n4584 S.t2361 6.541
R34156 S.n4567 S.n4566 6.541
R34157 S.n2828 S.n2827 6.541
R34158 S.n2839 S.t2924 6.541
R34159 S.n2836 S.t508 6.541
R34160 S.n2831 S.n2830 6.541
R34161 S.n3424 S.n3423 6.541
R34162 S.n3441 S.t2992 6.541
R34163 S.n3444 S.t1280 6.541
R34164 S.n3427 S.n3426 6.541
R34165 S.n1657 S.n1656 6.541
R34166 S.n1668 S.t1888 6.541
R34167 S.n1665 S.t3962 6.541
R34168 S.n1660 S.n1659 6.541
R34169 S.n2269 S.n2268 6.541
R34170 S.n2286 S.t1946 6.541
R34171 S.n2289 S.t264 6.541
R34172 S.n2272 S.n2271 6.541
R34173 S.n632 S.n631 6.541
R34174 S.n643 S.t845 6.541
R34175 S.n640 S.t2942 6.541
R34176 S.n635 S.n634 6.541
R34177 S.n615 S.n614 6.541
R34178 S.n626 S.t2399 6.541
R34179 S.n623 S.t4496 6.541
R34180 S.n618 S.n617 6.541
R34181 S.n1243 S.t4459 6.541
R34182 S.n272 S.n271 6.541
R34183 S.n283 S.t1022 6.541
R34184 S.n280 S.t3882 6.541
R34185 S.n275 S.n274 6.541
R34186 S.n2365 S.n2364 6.541
R34187 S.n2375 S.t2104 6.541
R34188 S.n2378 S.t411 6.541
R34189 S.n2362 S.n2361 6.541
R34190 S.n10335 S.t2235 6.541
R34191 S.n10759 S.n10758 6.541
R34192 S.n10776 S.t173 6.541
R34193 S.n10773 S.t3020 6.541
R34194 S.n10756 S.n10755 6.541
R34195 S.n9295 S.n9294 6.541
R34196 S.n9306 S.t3597 6.541
R34197 S.n9303 S.t1136 6.541
R34198 S.n9292 S.n9291 6.541
R34199 S.n10147 S.n10146 6.541
R34200 S.n10159 S.t4121 6.541
R34201 S.n10162 S.t1974 6.541
R34202 S.n10144 S.n10143 6.541
R34203 S.n8255 S.n8254 6.541
R34204 S.n8266 S.t2526 6.541
R34205 S.n8263 S.t660 6.541
R34206 S.n8252 S.n8251 6.541
R34207 S.n9080 S.n9079 6.541
R34208 S.n9092 S.t3141 6.541
R34209 S.n9095 S.t926 6.541
R34210 S.n9077 S.n9076 6.541
R34211 S.n7191 S.n7190 6.541
R34212 S.n7202 S.t1521 6.541
R34213 S.n7199 S.t4079 6.541
R34214 S.n7188 S.n7187 6.541
R34215 S.n8005 S.n8004 6.541
R34216 S.n8017 S.t2321 6.541
R34217 S.n8020 S.t4392 6.541
R34218 S.n8002 S.n8001 6.541
R34219 S.n6114 S.n6113 6.541
R34220 S.n6125 S.t465 6.541
R34221 S.n6122 S.t3309 6.541
R34222 S.n6111 S.n6110 6.541
R34223 S.n6907 S.n6906 6.541
R34224 S.n6919 S.t1234 6.541
R34225 S.n6922 S.t3367 6.541
R34226 S.n6904 S.n6903 6.541
R34227 S.n5014 S.n5013 6.541
R34228 S.n5025 S.t3930 6.541
R34229 S.n5022 S.t2710 6.541
R34230 S.n5011 S.n5010 6.541
R34231 S.n5797 S.n5796 6.541
R34232 S.n5809 S.t714 6.541
R34233 S.n5812 S.t2779 6.541
R34234 S.n5794 S.n5793 6.541
R34235 S.n3902 S.n3901 6.541
R34236 S.n3913 S.t3383 6.541
R34237 S.n3910 S.t1713 6.541
R34238 S.n3899 S.n3898 6.541
R34239 S.n4662 S.n4661 6.541
R34240 S.n4674 S.t4136 6.541
R34241 S.n4677 S.t2289 6.541
R34242 S.n4659 S.n4658 6.541
R34243 S.n2775 S.n2774 6.541
R34244 S.n2786 S.t2831 6.541
R34245 S.n2783 S.t667 6.541
R34246 S.n2772 S.n2771 6.541
R34247 S.n3521 S.n3520 6.541
R34248 S.n3532 S.t3153 6.541
R34249 S.n3535 S.t1191 6.541
R34250 S.n3518 S.n3517 6.541
R34251 S.n1602 S.n1601 6.541
R34252 S.n1614 S.t1814 6.541
R34253 S.n1611 S.t4089 6.541
R34254 S.n1599 S.n1598 6.541
R34255 S.n1400 S.t2905 6.541
R34256 S.n1010 S.n1009 6.541
R34257 S.n1013 S.t3986 6.541
R34258 S.n1016 S.t2347 6.541
R34259 S.n1019 S.n1018 6.541
R34260 S.n11359 S.t1720 6.541
R34261 S.n11786 S.n11785 6.541
R34262 S.n11804 S.t4144 6.541
R34263 S.n11801 S.t2485 6.541
R34264 S.n11789 S.n11788 6.541
R34265 S.n10343 S.n10342 6.541
R34266 S.n10354 S.t3095 6.541
R34267 S.n10351 S.t673 6.541
R34268 S.n10346 S.n10345 6.541
R34269 S.n11150 S.n11149 6.541
R34270 S.n11167 S.t3159 6.541
R34271 S.n11170 S.t1461 6.541
R34272 S.n11153 S.n11152 6.541
R34273 S.n9314 S.n9313 6.541
R34274 S.n9325 S.t2046 6.541
R34275 S.n9322 S.t4093 6.541
R34276 S.n9317 S.n9316 6.541
R34277 S.n10110 S.n10109 6.541
R34278 S.n10127 S.t2578 6.541
R34279 S.n10130 S.t420 6.541
R34280 S.n10113 S.n10112 6.541
R34281 S.n8272 S.n8271 6.541
R34282 S.n8283 S.t977 6.541
R34283 S.n8280 S.t3616 6.541
R34284 S.n8275 S.n8274 6.541
R34285 S.n9043 S.n9042 6.541
R34286 S.n9060 S.t1802 6.541
R34287 S.n9063 S.t3892 6.541
R34288 S.n9046 S.n9045 6.541
R34289 S.n7208 S.n7207 6.541
R34290 S.n7219 S.t4467 6.541
R34291 S.n7216 S.t2764 6.541
R34292 S.n7211 S.n7210 6.541
R34293 S.n7968 S.n7967 6.541
R34294 S.n7985 S.t767 6.541
R34295 S.n7988 S.t2838 6.541
R34296 S.n7971 S.n7970 6.541
R34297 S.n6131 S.n6130 6.541
R34298 S.n6142 S.t3426 6.541
R34299 S.n6139 S.t4116 6.541
R34300 S.n6134 S.n6133 6.541
R34301 S.n6870 S.n6869 6.541
R34302 S.n6887 S.t2137 6.541
R34303 S.n6890 S.t4181 6.541
R34304 S.n6873 S.n6872 6.541
R34305 S.n5031 S.n5030 6.541
R34306 S.n5042 S.t284 6.541
R34307 S.n5039 S.t1151 6.541
R34308 S.n5034 S.n5033 6.541
R34309 S.n5760 S.n5759 6.541
R34310 S.n5777 S.t3672 6.541
R34311 S.n5780 S.t1217 6.541
R34312 S.n5763 S.n5762 6.541
R34313 S.n3919 S.n3918 6.541
R34314 S.n3930 S.t1837 6.541
R34315 S.n3927 S.t117 6.541
R34316 S.n3922 S.n3921 6.541
R34317 S.n4625 S.n4624 6.541
R34318 S.n4642 S.t2590 6.541
R34319 S.n4645 S.t725 6.541
R34320 S.n4628 S.n4627 6.541
R34321 S.n2792 S.n2791 6.541
R34322 S.n2803 S.t1263 6.541
R34323 S.n2800 S.t3628 6.541
R34324 S.n2795 S.n2794 6.541
R34325 S.n3484 S.n3483 6.541
R34326 S.n3501 S.t1598 6.541
R34327 S.n3504 S.t4401 6.541
R34328 S.n3487 S.n3486 6.541
R34329 S.n1620 S.n1619 6.541
R34330 S.n1631 S.t473 6.541
R34331 S.n1628 S.t2546 6.541
R34332 S.n1623 S.n1622 6.541
R34333 S.n2328 S.n2327 6.541
R34334 S.n2345 S.t536 6.541
R34335 S.n2348 S.t3374 6.541
R34336 S.n2331 S.n2330 6.541
R34337 S.n597 S.n596 6.541
R34338 S.n608 S.t3937 6.541
R34339 S.n605 S.t1549 6.541
R34340 S.n600 S.n599 6.541
R34341 S.n580 S.n579 6.541
R34342 S.n591 S.t970 6.541
R34343 S.n588 S.t3102 6.541
R34344 S.n583 S.n582 6.541
R34345 S.n1230 S.t2810 6.541
R34346 S.n243 S.n242 6.541
R34347 S.n251 S.t4115 6.541
R34348 S.n222 S.t2269 6.541
R34349 S.n246 S.n245 6.541
R34350 S.n2424 S.n2423 6.541
R34351 S.n2434 S.t695 6.541
R34352 S.n2437 S.t3296 6.541
R34353 S.n2421 S.n2420 6.541
R34354 S.n8228 S.t3761 6.541
R34355 S.n8656 S.n8655 6.541
R34356 S.n8673 S.t1724 6.541
R34357 S.n8670 S.t4010 6.541
R34358 S.n8653 S.n8652 6.541
R34359 S.n7153 S.n7152 6.541
R34360 S.n7164 S.t48 6.541
R34361 S.n7161 S.t2678 6.541
R34362 S.n7150 S.n7149 6.541
R34363 S.n8070 S.n8069 6.541
R34364 S.n8082 S.t684 6.541
R34365 S.n8085 S.t3004 6.541
R34366 S.n8067 S.n8066 6.541
R34367 S.n6078 S.n6077 6.541
R34368 S.n6089 S.t3574 6.541
R34369 S.n6086 S.t1685 6.541
R34370 S.n6075 S.n6074 6.541
R34371 S.n6968 S.n6967 6.541
R34372 S.n6980 S.t4100 6.541
R34373 S.n6983 S.t1958 6.541
R34374 S.n6965 S.n6964 6.541
R34375 S.n4978 S.n4977 6.541
R34376 S.n4989 S.t2511 6.541
R34377 S.n4986 S.t3225 6.541
R34378 S.n4975 S.n4974 6.541
R34379 S.n5858 S.n5857 6.541
R34380 S.n5870 S.t1391 6.541
R34381 S.n5873 S.t3489 6.541
R34382 S.n5855 S.n5854 6.541
R34383 S.n3866 S.n3865 6.541
R34384 S.n3877 S.t4044 6.541
R34385 S.n3874 S.t2397 6.541
R34386 S.n3863 S.n3862 6.541
R34387 S.n4723 S.n4722 6.541
R34388 S.n4735 S.t359 6.541
R34389 S.n4738 S.t2968 6.541
R34390 S.n4720 S.n4719 6.541
R34391 S.n2739 S.n2738 6.541
R34392 S.n2750 S.t3537 6.541
R34393 S.n2747 S.t3774 6.541
R34394 S.n2736 S.n2735 6.541
R34395 S.n3581 S.n3580 6.541
R34396 S.n3592 S.t1737 6.541
R34397 S.n3595 S.t4310 6.541
R34398 S.n3578 S.n3577 6.541
R34399 S.n1565 S.n1564 6.541
R34400 S.n1577 S.t396 6.541
R34401 S.n1574 S.t2689 6.541
R34402 S.n1562 S.n1561 6.541
R34403 S.n1396 S.t1514 6.541
R34404 S.n1042 S.n1041 6.541
R34405 S.n1045 S.t2572 6.541
R34406 S.n1048 S.t919 6.541
R34407 S.n1051 S.n1050 6.541
R34408 S.n9287 S.t2695 6.541
R34409 S.n9718 S.n9717 6.541
R34410 S.n9736 S.t1166 6.541
R34411 S.n9733 S.t3520 6.541
R34412 S.n9721 S.n9720 6.541
R34413 S.n8236 S.n8235 6.541
R34414 S.n8247 S.t4067 6.541
R34415 S.n8244 S.t2221 6.541
R34416 S.n8239 S.n8238 6.541
R34417 S.n9108 S.n9107 6.541
R34418 S.n9125 S.t142 6.541
R34419 S.n9128 S.t2470 6.541
R34420 S.n9111 S.n9110 6.541
R34421 S.n7172 S.n7171 6.541
R34422 S.n7183 S.t3072 6.541
R34423 S.n7180 S.t1121 6.541
R34424 S.n7175 S.n7174 6.541
R34425 S.n8033 S.n8032 6.541
R34426 S.n8050 S.t3642 6.541
R34427 S.n8053 S.t1444 6.541
R34428 S.n8036 S.n8035 6.541
R34429 S.n6095 S.n6094 6.541
R34430 S.n6106 S.t2023 6.541
R34431 S.n6103 S.t72 6.541
R34432 S.n6098 S.n6097 6.541
R34433 S.n6931 S.n6930 6.541
R34434 S.n6948 S.t2796 6.541
R34435 S.n6951 S.t404 6.541
R34436 S.n6934 S.n6933 6.541
R34437 S.n4995 S.n4994 6.541
R34438 S.n5006 S.t963 6.541
R34439 S.n5003 S.t1886 6.541
R34440 S.n4998 S.n4997 6.541
R34441 S.n5821 S.n5820 6.541
R34442 S.n5838 S.t4339 6.541
R34443 S.n5841 S.t1942 6.541
R34444 S.n5824 S.n5823 6.541
R34445 S.n3883 S.n3882 6.541
R34446 S.n3894 S.t2502 6.541
R34447 S.n3891 S.t3266 6.541
R34448 S.n3886 S.n3885 6.541
R34449 S.n4686 S.n4685 6.541
R34450 S.n4703 S.t1181 6.541
R34451 S.n4706 S.t3827 6.541
R34452 S.n4689 S.n4688 6.541
R34453 S.n2756 S.n2755 6.541
R34454 S.n2767 S.t4388 6.541
R34455 S.n2764 S.t2230 6.541
R34456 S.n2759 S.n2758 6.541
R34457 S.n3544 S.n3543 6.541
R34458 S.n3561 S.t164 6.541
R34459 S.n3564 S.t2750 6.541
R34460 S.n3547 S.n3546 6.541
R34461 S.n1583 S.n1582 6.541
R34462 S.n1594 S.t3360 6.541
R34463 S.n1591 S.t1132 6.541
R34464 S.n1586 S.n1585 6.541
R34465 S.n2387 S.n2386 6.541
R34466 S.n2404 S.t3658 6.541
R34467 S.n2407 S.t1749 6.541
R34468 S.n2390 S.n2389 6.541
R34469 S.n562 S.n561 6.541
R34470 S.n573 S.t2334 6.541
R34471 S.n570 S.t96 6.541
R34472 S.n565 S.n564 6.541
R34473 S.n545 S.n544 6.541
R34474 S.n556 S.t3869 6.541
R34475 S.n553 S.t1697 6.541
R34476 S.n548 S.n547 6.541
R34477 S.n1217 S.t1415 6.541
R34478 S.n208 S.n207 6.541
R34479 S.n219 S.t2719 6.541
R34480 S.n216 S.t846 6.541
R34481 S.n211 S.n210 6.541
R34482 S.n2483 S.n2482 6.541
R34483 S.n2493 S.t1372 6.541
R34484 S.n2496 S.t3967 6.541
R34485 S.n2480 S.n2479 6.541
R34486 S.n6051 S.t260 6.541
R34487 S.n6483 S.n6482 6.541
R34488 S.n6500 S.t2705 6.541
R34489 S.n6497 S.t548 6.541
R34490 S.n6480 S.n6479 6.541
R34491 S.n4940 S.n4939 6.541
R34492 S.n4951 S.t1086 6.541
R34493 S.n4948 S.t1813 6.541
R34494 S.n4937 S.n4936 6.541
R34495 S.n5923 S.n5922 6.541
R34496 S.n5935 S.t4244 6.541
R34497 S.n5938 S.t2102 6.541
R34498 S.n5920 S.n5919 6.541
R34499 S.n3830 S.n3829 6.541
R34500 S.n3841 S.t2634 6.541
R34501 S.n3838 S.t777 6.541
R34502 S.n3827 S.n3826 6.541
R34503 S.n4784 S.n4783 6.541
R34504 S.n4796 S.t3256 6.541
R34505 S.n4799 S.t1576 6.541
R34506 S.n4781 S.n4780 6.541
R34507 S.n2703 S.n2702 6.541
R34508 S.n2714 S.t2151 6.541
R34509 S.n2711 S.t4195 6.541
R34510 S.n2700 S.n2699 6.541
R34511 S.n3641 S.n3640 6.541
R34512 S.n3652 S.t2419 6.541
R34513 S.n3655 S.t514 6.541
R34514 S.n3638 S.n3637 6.541
R34515 S.n1528 S.n1527 6.541
R34516 S.n1540 S.t1054 6.541
R34517 S.n1537 S.t3416 6.541
R34518 S.n1525 S.n1524 6.541
R34519 S.n1392 S.t4363 6.541
R34520 S.n1074 S.n1073 6.541
R34521 S.n1077 S.t1161 6.541
R34522 S.n1080 S.t3811 6.541
R34523 S.n1083 S.n1082 6.541
R34524 S.n7145 S.t4230 6.541
R34525 S.n7580 S.n7579 6.541
R34526 S.n7598 S.t2243 6.541
R34527 S.n7595 S.t4561 6.541
R34528 S.n7583 S.n7582 6.541
R34529 S.n6059 S.n6058 6.541
R34530 S.n6070 S.t624 6.541
R34531 S.n6067 S.t3238 6.541
R34532 S.n6062 S.n6061 6.541
R34533 S.n6996 S.n6995 6.541
R34534 S.n7013 S.t1147 6.541
R34535 S.n7016 S.t3504 6.541
R34536 S.n6999 S.n6998 6.541
R34537 S.n4959 S.n4958 6.541
R34538 S.n4970 S.t4050 6.541
R34539 S.n4967 S.t245 6.541
R34540 S.n4962 S.n4961 6.541
R34541 S.n5886 S.n5885 6.541
R34542 S.n5903 S.t2692 6.541
R34543 S.n5906 S.t533 6.541
R34544 S.n5889 S.n5888 6.541
R34545 S.n3847 S.n3846 6.541
R34546 S.n3858 S.t1079 6.541
R34547 S.n3855 S.t3730 6.541
R34548 S.n3850 S.n3849 6.541
R34549 S.n4747 S.n4746 6.541
R34550 S.n4764 S.t1916 6.541
R34551 S.n4767 S.t4530 6.541
R34552 S.n4750 S.n4749 6.541
R34553 S.n2720 S.n2719 6.541
R34554 S.n2731 S.t586 6.541
R34555 S.n2728 S.t2903 6.541
R34556 S.n2723 S.n2722 6.541
R34557 S.n3604 S.n3603 6.541
R34558 S.n3621 S.t874 6.541
R34559 S.n3624 S.t3472 6.541
R34560 S.n3607 S.n3606 6.541
R34561 S.n1546 S.n1545 6.541
R34562 S.n1557 S.t4024 6.541
R34563 S.n1554 S.t4240 6.541
R34564 S.n1549 S.n1548 6.541
R34565 S.n2446 S.n2445 6.541
R34566 S.n2463 S.t2255 6.541
R34567 S.n2466 S.t329 6.541
R34568 S.n2449 S.n2448 6.541
R34569 S.n527 S.n526 6.541
R34570 S.n538 S.t906 6.541
R34571 S.n535 S.t3252 6.541
R34572 S.n530 S.n529 6.541
R34573 S.n510 S.n509 6.541
R34574 S.n521 S.t4578 6.541
R34575 S.n518 S.t274 6.541
R34576 S.n513 S.n512 6.541
R34577 S.n1204 S.t2132 6.541
R34578 S.n176 S.n175 6.541
R34579 S.n187 S.t3445 6.541
R34580 S.n184 S.t1558 6.541
R34581 S.n179 S.n178 6.541
R34582 S.n2542 S.n2541 6.541
R34583 S.n2552 S.t4225 6.541
R34584 S.n2555 S.t2550 6.541
R34585 S.n2539 S.n2538 6.541
R34586 S.n3803 S.t3867 6.541
R34587 S.n4238 S.n4237 6.541
R34588 S.n4255 S.t1844 6.541
R34589 S.n4252 S.t125 6.541
R34590 S.n4235 S.n4234 6.541
R34591 S.n2665 S.n2664 6.541
R34592 S.n2676 S.t741 6.541
R34593 S.n2673 S.t2806 6.541
R34594 S.n2662 S.n2661 6.541
R34595 S.n3705 S.n3704 6.541
R34596 S.n3716 S.t805 6.541
R34597 S.n3719 S.t3633 6.541
R34598 S.n3702 S.n3701 6.541
R34599 S.n1491 S.n1490 6.541
R34600 S.n1503 S.t4159 6.541
R34601 S.n1500 S.t1792 6.541
R34602 S.n1488 S.n1487 6.541
R34603 S.n1388 S.t565 6.541
R34604 S.n1106 S.n1105 6.541
R34605 S.n1109 S.t1901 6.541
R34606 S.n1112 S.t4503 6.541
R34607 S.n1115 S.n1114 6.541
R34608 S.n4932 S.t3359 6.541
R34609 S.n5371 S.n5370 6.541
R34610 S.n5389 S.t1295 6.541
R34611 S.n5386 S.t3651 6.541
R34612 S.n5374 S.n5373 6.541
R34613 S.n3811 S.n3810 6.541
R34614 S.n3822 S.t4182 6.541
R34615 S.n3819 S.t2329 6.541
R34616 S.n3814 S.n3813 6.541
R34617 S.n4812 S.n4811 6.541
R34618 S.n4829 S.t281 6.541
R34619 S.n4832 S.t3129 6.541
R34620 S.n4815 S.n4814 6.541
R34621 S.n2684 S.n2683 6.541
R34622 S.n2695 S.t3697 6.541
R34623 S.n2692 S.t1242 6.541
R34624 S.n2687 S.n2686 6.541
R34625 S.n3668 S.n3667 6.541
R34626 S.n3685 S.t3760 6.541
R34627 S.n3688 S.t2079 6.541
R34628 S.n3671 S.n3670 6.541
R34629 S.n1509 S.n1508 6.541
R34630 S.n1520 S.t2609 6.541
R34631 S.n1517 S.t227 6.541
R34632 S.n1512 S.n1511 6.541
R34633 S.n2505 S.n2504 6.541
R34634 S.n2522 S.t2937 6.541
R34635 S.n2525 S.t1004 6.541
R34636 S.n2508 S.n2507 6.541
R34637 S.n492 S.n491 6.541
R34638 S.n503 S.t1622 6.541
R34639 S.n500 S.t3919 6.541
R34640 S.n495 S.n494 6.541
R34641 S.n475 S.n474 6.541
R34642 S.n486 S.t3172 6.541
R34643 S.n483 S.t754 6.541
R34644 S.n478 S.n477 6.541
R34645 S.n1191 S.t719 6.541
R34646 S.n144 S.n143 6.541
R34647 S.n155 S.t1825 6.541
R34648 S.n152 S.t104 6.541
R34649 S.n147 S.n146 6.541
R34650 S.n1944 S.n1943 6.541
R34651 S.n1959 S.t2845 6.541
R34652 S.n1956 S.t1135 6.541
R34653 S.n1941 S.n1940 6.541
R34654 S.n1464 S.t375 6.541
R34655 S.n1384 S.t3679 6.541
R34656 S.n1144 S.n1143 6.541
R34657 S.n1147 S.t257 6.541
R34658 S.n1150 S.t3110 6.541
R34659 S.n1153 S.n1152 6.541
R34660 S.n2657 S.t4360 6.541
R34661 S.n3101 S.n3100 6.541
R34662 S.n3119 S.t2359 6.541
R34663 S.n3116 S.t672 6.541
R34664 S.n3104 S.n3103 6.541
R34665 S.n1472 S.n1471 6.541
R34666 S.n1483 S.t1206 6.541
R34667 S.n1480 S.t3341 6.541
R34668 S.n1475 S.n1474 6.541
R34669 S.n2568 S.n2567 6.541
R34670 S.n2585 S.t1276 6.541
R34671 S.n2588 S.t4091 6.541
R34672 S.n2571 S.n2570 6.541
R34673 S.n457 S.n456 6.541
R34674 S.n468 S.t191 6.541
R34675 S.n465 S.t2315 6.541
R34676 S.n460 S.n459 6.541
R34677 S.n441 S.n440 6.541
R34678 S.n452 S.t1761 6.541
R34679 S.n449 S.t3851 6.541
R34680 S.n444 S.n443 6.541
R34681 S.n1380 S.t2283 6.541
R34682 S.n931 S.n930 6.541
R34683 S.n944 S.t3370 6.541
R34684 S.n947 S.t1702 6.541
R34685 S.n934 S.n933 6.541
R34686 S.n436 S.t890 6.541
R34687 S.n1430 S.t3934 6.541
R34688 S.n22309 S.n22308 6.541
R34689 S.n22312 S.t1170 6.541
R34690 S.n21970 S.t4382 6.541
R34691 S.n21972 S.t2063 6.541
R34692 S.n22995 S.t1693 6.541
R34693 S.n22993 S.t958 6.541
R34694 S.n22759 S.n22758 6.541
R34695 S.n22767 S.t2566 6.541
R34696 S.n22770 S.t4535 6.541
R34697 S.n22762 S.n22761 6.541
R34698 S.n21322 S.n21321 6.541
R34699 S.n21333 S.t3406 6.541
R34700 S.n21330 S.t1418 6.541
R34701 S.n21325 S.n21324 6.541
R34702 S.n22302 S.n22301 6.541
R34703 S.n22305 S.t111 6.541
R34704 S.n22335 S.n22334 6.541
R34705 S.n22338 S.t853 6.541
R34706 S.n22330 S.n22329 6.541
R34707 S.n22315 S.t1808 6.541
R34708 S.n20177 S.t2439 6.105
R34709 S.n20185 S.n20184 6.105
R34710 S.n20188 S.n20187 6.105
R34711 S.n20180 S.t157 6.105
R34712 S.n21131 S.t3681 6.105
R34713 S.n21135 S.n21134 6.105
R34714 S.n21138 S.n21137 6.105
R34715 S.n21128 S.t1443 6.105
R34716 S.n22958 S.t3945 6.105
R34717 S.n22637 S.t2874 6.105
R34718 S.n22642 S.n22641 6.105
R34719 S.n22645 S.n22644 6.105
R34720 S.n22634 S.t4430 6.105
R34721 S.n22008 S.t1039 6.105
R34722 S.n22015 S.n22014 6.105
R34723 S.n22012 S.n22011 6.105
R34724 S.n22005 S.t2044 6.105
R34725 S.n21614 S.t2979 6.105
R34726 S.n21619 S.n21618 6.105
R34727 S.n21622 S.n21621 6.105
R34728 S.n21611 S.t1665 6.105
R34729 S.n21940 S.t2645 6.105
R34730 S.n21944 S.n21943 6.105
R34731 S.n21947 S.n21946 6.105
R34732 S.n21937 S.t3654 6.105
R34733 S.n20791 S.t2923 6.105
R34734 S.n20796 S.n20795 6.105
R34735 S.n20799 S.n20798 6.105
R34736 S.n20788 S.t1616 6.105
R34737 S.n21145 S.t763 6.105
R34738 S.n22965 S.t2409 6.105
R34739 S.n22650 S.t1307 6.105
R34740 S.n22658 S.n22657 6.105
R34741 S.n22661 S.n22660 6.105
R34742 S.n22653 S.t2875 6.105
R34743 S.n21989 S.t4004 6.105
R34744 S.n22000 S.n21999 6.105
R34745 S.n21997 S.n21996 6.105
R34746 S.n21992 S.t484 6.105
R34747 S.n21632 S.t1413 6.105
R34748 S.n21640 S.n21639 6.105
R34749 S.n21643 S.n21642 6.105
R34750 S.n21635 S.t28 6.105
R34751 S.n21955 S.t1188 6.105
R34752 S.n21964 S.n21963 6.105
R34753 S.n21967 S.n21966 6.105
R34754 S.n21958 S.t3506 6.105
R34755 S.n20809 S.t4526 6.105
R34756 S.n20820 S.n20819 6.105
R34757 S.n20823 S.n20822 6.105
R34758 S.n20812 S.t2202 6.105
R34759 S.n20340 S.t2275 6.105
R34760 S.n19307 S.t378 6.105
R34761 S.n19315 S.n19314 6.105
R34762 S.n19318 S.n19317 6.105
R34763 S.n19310 S.t2643 6.105
R34764 S.n19531 S.t1621 6.105
R34765 S.n19538 S.n19537 6.105
R34766 S.n19535 S.n19534 6.105
R34767 S.n19528 S.t3891 6.105
R34768 S.n22951 S.t978 6.105
R34769 S.n22621 S.t4429 6.105
R34770 S.n22626 S.n22625 6.105
R34771 S.n22629 S.n22628 6.105
R34772 S.n22618 S.t1482 6.105
R34773 S.n22023 S.t2592 6.105
R34774 S.n22030 S.n22029 6.105
R34775 S.n22027 S.n22026 6.105
R34776 S.n22020 S.t3599 6.105
R34777 S.n21598 S.t4539 6.105
R34778 S.n21603 S.n21602 6.105
R34779 S.n21606 S.n21605 6.105
R34780 S.n21595 S.t3211 6.105
R34781 S.n21925 S.t4193 6.105
R34782 S.n21929 S.n21928 6.105
R34783 S.n21932 S.n21931 6.105
R34784 S.n21922 S.t697 6.105
R34785 S.n20775 S.t4477 6.105
R34786 S.n20780 S.n20779 6.105
R34787 S.n20783 S.n20782 6.105
R34788 S.n20772 S.t3169 6.105
R34789 S.n21115 S.t4145 6.105
R34790 S.n21119 S.n21118 6.105
R34791 S.n21122 S.n21121 6.105
R34792 S.n21112 S.t654 6.105
R34793 S.n20164 S.t4423 6.105
R34794 S.n20169 S.n20168 6.105
R34795 S.n20172 S.n20171 6.105
R34796 S.n20161 S.t3122 6.105
R34797 S.n19500 S.t3775 6.105
R34798 S.n18425 S.t2814 6.105
R34799 S.n18433 S.n18432 6.105
R34800 S.n18436 S.n18435 6.105
R34801 S.n18428 S.t678 6.105
R34802 S.n18674 S.t682 6.105
R34803 S.n18681 S.n18680 6.105
R34804 S.n18678 S.n18677 6.105
R34805 S.n18671 S.t1834 6.105
R34806 S.n22944 S.t2344 6.105
R34807 S.n22605 S.t1479 6.105
R34808 S.n22610 S.n22609 6.105
R34809 S.n22613 S.n22612 6.105
R34810 S.n22602 S.t3037 6.105
R34811 S.n22038 S.t4137 6.105
R34812 S.n22045 S.n22044 6.105
R34813 S.n22042 S.n22041 6.105
R34814 S.n22035 S.t644 6.105
R34815 S.n21582 S.t1584 6.105
R34816 S.n21587 S.n21586 6.105
R34817 S.n21590 S.n21589 6.105
R34818 S.n21579 S.t235 6.105
R34819 S.n21910 S.t1238 6.105
R34820 S.n21914 S.n21913 6.105
R34821 S.n21917 S.n21916 6.105
R34822 S.n21907 S.t2257 6.105
R34823 S.n20759 S.t1532 6.105
R34824 S.n20764 S.n20763 6.105
R34825 S.n20767 S.n20766 6.105
R34826 S.n20756 S.t182 6.105
R34827 S.n21100 S.t1187 6.105
R34828 S.n21104 S.n21103 6.105
R34829 S.n21107 S.n21106 6.105
R34830 S.n21097 S.t2215 6.105
R34831 S.n20148 S.t1473 6.105
R34832 S.n20153 S.n20152 6.105
R34833 S.n20156 S.n20155 6.105
R34834 S.n20145 S.t115 6.105
R34835 S.n19546 S.t1142 6.105
R34836 S.n19553 S.n19552 6.105
R34837 S.n19550 S.n19549 6.105
R34838 S.n19543 S.t2161 6.105
R34839 S.n19294 S.t1423 6.105
R34840 S.n19299 S.n19298 6.105
R34841 S.n19302 S.n19301 6.105
R34842 S.n19291 S.t40 6.105
R34843 S.n18643 S.t3750 6.105
R34844 S.n17520 S.t782 6.105
R34845 S.n17528 S.n17527 6.105
R34846 S.n17531 S.n17530 6.105
R34847 S.n17523 S.t3191 6.105
R34848 S.n17806 S.t3139 6.105
R34849 S.n17813 S.n17812 6.105
R34850 S.n17810 S.n17809 6.105
R34851 S.n17803 S.t891 6.105
R34852 S.n22937 S.t3877 6.105
R34853 S.n22589 S.t3036 6.105
R34854 S.n22594 S.n22593 6.105
R34855 S.n22597 S.n22596 6.105
R34856 S.n22586 S.t4597 6.105
R34857 S.n22053 S.t974 6.105
R34858 S.n22060 S.n22059 6.105
R34859 S.n22057 S.n22056 6.105
R34860 S.n22050 S.t1961 6.105
R34861 S.n21566 S.t3137 6.105
R34862 S.n21571 S.n21570 6.105
R34863 S.n21574 S.n21573 6.105
R34864 S.n21563 S.t1799 6.105
R34865 S.n21895 S.t2803 6.105
R34866 S.n21899 S.n21898 6.105
R34867 S.n21902 S.n21901 6.105
R34868 S.n21892 S.t3800 6.105
R34869 S.n20743 S.t3086 6.105
R34870 S.n20748 S.n20747 6.105
R34871 S.n20751 S.n20750 6.105
R34872 S.n20740 S.t1752 6.105
R34873 S.n21085 S.t2746 6.105
R34874 S.n21089 S.n21088 6.105
R34875 S.n21092 S.n21091 6.105
R34876 S.n21082 S.t3758 6.105
R34877 S.n20132 S.t3032 6.105
R34878 S.n20137 S.n20136 6.105
R34879 S.n20140 S.n20139 6.105
R34880 S.n20129 S.t1709 6.105
R34881 S.n19561 S.t2698 6.105
R34882 S.n19568 S.n19567 6.105
R34883 S.n19565 S.n19564 6.105
R34884 S.n19558 S.t3707 6.105
R34885 S.n19278 S.t2984 6.105
R34886 S.n19283 S.n19282 6.105
R34887 S.n19286 S.n19285 6.105
R34888 S.n19275 S.t1669 6.105
R34889 S.n18689 S.t1119 6.105
R34890 S.n18696 S.n18695 6.105
R34891 S.n18693 S.n18692 6.105
R34892 S.n18686 S.t3663 6.105
R34893 S.n18412 S.t2934 6.105
R34894 S.n18417 S.n18416 6.105
R34895 S.n18420 S.n18419 6.105
R34896 S.n18409 S.t1625 6.105
R34897 S.n17775 S.t746 6.105
R34898 S.n16602 S.t3227 6.105
R34899 S.n16610 S.n16609 6.105
R34900 S.n16613 S.n16612 6.105
R34901 S.n16605 S.t1128 6.105
R34902 S.n16912 S.t1029 6.105
R34903 S.n16919 S.n16918 6.105
R34904 S.n16916 S.n16915 6.105
R34905 S.n16909 S.t3338 6.105
R34906 S.n22930 S.t915 6.105
R34907 S.n22573 S.t4596 6.105
R34908 S.n22578 S.n22577 6.105
R34909 S.n22581 S.n22580 6.105
R34910 S.n22570 S.t1641 6.105
R34911 S.n22068 S.t2522 6.105
R34912 S.n22075 S.n22074 6.105
R34913 S.n22072 S.n22071 6.105
R34914 S.n22065 S.t3510 6.105
R34915 S.n21550 S.t136 6.105
R34916 S.n21555 S.n21554 6.105
R34917 S.n21558 S.n21557 6.105
R34918 S.n21547 S.t3345 6.105
R34919 S.n21880 S.t4106 6.105
R34920 S.n21884 S.n21883 6.105
R34921 S.n21887 S.n21886 6.105
R34922 S.n21877 S.t618 6.105
R34923 S.n20727 S.t65 6.105
R34924 S.n20732 S.n20731 6.105
R34925 S.n20735 S.n20734 6.105
R34926 S.n20724 S.t3301 6.105
R34927 S.n21070 S.t4303 6.105
R34928 S.n21074 S.n21073 6.105
R34929 S.n21077 S.n21076 6.105
R34930 S.n21067 S.t804 6.105
R34931 S.n20116 S.t4589 6.105
R34932 S.n20121 S.n20120 6.105
R34933 S.n20124 S.n20123 6.105
R34934 S.n20113 S.t3263 6.105
R34935 S.n19576 S.t4248 6.105
R34936 S.n19583 S.n19582 6.105
R34937 S.n19580 S.n19579 6.105
R34938 S.n19573 S.t751 6.105
R34939 S.n19262 S.t4544 6.105
R34940 S.n19267 S.n19266 6.105
R34941 S.n19270 S.n19269 6.105
R34942 S.n19259 S.t3219 6.105
R34943 S.n18704 S.t2675 6.105
R34944 S.n18711 S.n18710 6.105
R34945 S.n18708 S.n18707 6.105
R34946 S.n18701 S.t702 6.105
R34947 S.n18396 S.t4486 6.105
R34948 S.n18401 S.n18400 6.105
R34949 S.n18404 S.n18403 6.105
R34950 S.n18393 S.t3174 6.105
R34951 S.n17821 S.t2628 6.105
R34952 S.n17828 S.n17827 6.105
R34953 S.n17825 S.n17824 6.105
R34954 S.n17818 S.t3639 6.105
R34955 S.n17507 S.t4440 6.105
R34956 S.n17512 S.n17511 6.105
R34957 S.n17515 S.n17514 6.105
R34958 S.n17504 S.t3131 6.105
R34959 S.n16881 S.t2260 6.105
R34960 S.n15662 S.t1108 6.105
R34961 S.n15670 S.n15669 6.105
R34962 S.n15673 S.n15672 6.105
R34963 S.n15665 S.t3677 6.105
R34964 S.n16009 S.t3496 6.105
R34965 S.n16016 S.n16015 6.105
R34966 S.n16013 S.n16012 6.105
R34967 S.n16006 S.t1240 6.105
R34968 S.n22923 S.t2460 6.105
R34969 S.n22557 S.t1642 6.105
R34970 S.n22562 S.n22561 6.105
R34971 S.n22565 S.n22564 6.105
R34972 S.n22554 S.t3194 6.105
R34973 S.n22083 S.t4060 6.105
R34974 S.n22090 S.n22089 6.105
R34975 S.n22087 S.n22086 6.105
R34976 S.n22080 S.t553 6.105
R34977 S.n21534 S.t1723 6.105
R34978 S.n21539 S.n21538 6.105
R34979 S.n21542 S.n21541 6.105
R34980 S.n21531 S.t377 6.105
R34981 S.n21865 S.t1153 6.105
R34982 S.n21869 S.n21868 6.105
R34983 S.n21872 S.n21871 6.105
R34984 S.n21862 S.t2179 6.105
R34985 S.n20711 S.t1682 6.105
R34986 S.n20716 S.n20715 6.105
R34987 S.n20719 S.n20718 6.105
R34988 S.n20708 S.t336 6.105
R34989 S.n21055 S.t1106 6.105
R34990 S.n21059 S.n21058 6.105
R34991 S.n21062 S.n21061 6.105
R34992 S.n21052 S.t2129 6.105
R34993 S.n20100 S.t1636 6.105
R34994 S.n20105 S.n20104 6.105
R34995 S.n20108 S.n20107 6.105
R34996 S.n20097 S.t291 6.105
R34997 S.n19591 S.t1299 6.105
R34998 S.n19598 S.n19597 6.105
R34999 S.n19595 S.n19594 6.105
R35000 S.n19588 S.t2314 6.105
R35001 S.n19246 S.t1587 6.105
R35002 S.n19251 S.n19250 6.105
R35003 S.n19254 S.n19253 6.105
R35004 S.n19243 S.t240 6.105
R35005 S.n18719 S.t4227 6.105
R35006 S.n18726 S.n18725 6.105
R35007 S.n18723 S.n18722 6.105
R35008 S.n18716 S.t2264 6.105
R35009 S.n18380 S.t1541 6.105
R35010 S.n18385 S.n18384 6.105
R35011 S.n18388 S.n18387 6.105
R35012 S.n18377 S.t192 6.105
R35013 S.n17836 S.t4177 6.105
R35014 S.n17843 S.n17842 6.105
R35015 S.n17840 S.n17839 6.105
R35016 S.n17833 S.t681 6.105
R35017 S.n17491 S.t1490 6.105
R35018 S.n17496 S.n17495 6.105
R35019 S.n17499 S.n17498 6.105
R35020 S.n17488 S.t127 6.105
R35021 S.n16927 S.t4129 6.105
R35022 S.n16934 S.n16933 6.105
R35023 S.n16931 S.n16930 6.105
R35024 S.n16924 S.t638 6.105
R35025 S.n16589 S.t1434 6.105
R35026 S.n16594 S.n16593 6.105
R35027 S.n16597 S.n16596 6.105
R35028 S.n16586 S.t53 6.105
R35029 S.n15978 S.t3763 6.105
R35030 S.n14709 S.t3600 6.105
R35031 S.n14717 S.n14716 6.105
R35032 S.n14720 S.n14719 6.105
R35033 S.n14712 S.t1679 6.105
R35034 S.n15080 S.t1433 6.105
R35035 S.n15087 S.n15086 6.105
R35036 S.n15084 S.n15083 6.105
R35037 S.n15077 S.t3726 6.105
R35038 S.n22916 S.t1374 6.105
R35039 S.n22541 S.t3195 6.105
R35040 S.n22546 S.n22545 6.105
R35041 S.n22549 S.n22548 6.105
R35042 S.n22538 S.t213 6.105
R35043 S.n22098 S.t1100 6.105
R35044 S.n22105 S.n22104 6.105
R35045 S.n22102 S.n22101 6.105
R35046 S.n22095 S.t2119 6.105
R35047 S.n21518 S.t3275 6.105
R35048 S.n21523 S.n21522 6.105
R35049 S.n21526 S.n21525 6.105
R35050 S.n21515 S.t1937 6.105
R35051 S.n21850 S.t2711 6.105
R35052 S.n21854 S.n21853 6.105
R35053 S.n21857 S.n21856 6.105
R35054 S.n21847 S.t3723 6.105
R35055 S.n20695 S.t3233 6.105
R35056 S.n20700 S.n20699 6.105
R35057 S.n20703 S.n20702 6.105
R35058 S.n20692 S.t1895 6.105
R35059 S.n21040 S.t2663 6.105
R35060 S.n21044 S.n21043 6.105
R35061 S.n21047 S.n21046 6.105
R35062 S.n21037 S.t3676 6.105
R35063 S.n20084 S.t3188 6.105
R35064 S.n20089 S.n20088 6.105
R35065 S.n20092 S.n20091 6.105
R35066 S.n20081 S.t1852 6.105
R35067 S.n19606 S.t2615 6.105
R35068 S.n19613 S.n19612 6.105
R35069 S.n19610 S.n19609 6.105
R35070 S.n19603 S.t3631 6.105
R35071 S.n19230 S.t3145 6.105
R35072 S.n19235 S.n19234 6.105
R35073 S.n19238 S.n19237 6.105
R35074 S.n19227 S.t1806 6.105
R35075 S.n18734 S.t1277 6.105
R35076 S.n18741 S.n18740 6.105
R35077 S.n18738 S.n18737 6.105
R35078 S.n18731 S.t3806 6.105
R35079 S.n18364 S.t3092 6.105
R35080 S.n18369 S.n18368 6.105
R35081 S.n18372 S.n18371 6.105
R35082 S.n18361 S.t1762 6.105
R35083 S.n17851 S.t1226 6.105
R35084 S.n17858 S.n17857 6.105
R35085 S.n17855 S.n17854 6.105
R35086 S.n17848 S.t2242 6.105
R35087 S.n17475 S.t3045 6.105
R35088 S.n17480 S.n17479 6.105
R35089 S.n17483 S.n17482 6.105
R35090 S.n17472 S.t1717 6.105
R35091 S.n16942 S.t1174 6.105
R35092 S.n16949 S.n16948 6.105
R35093 S.n16946 S.n16945 6.105
R35094 S.n16939 S.t2201 6.105
R35095 S.n16573 S.t2994 6.105
R35096 S.n16578 S.n16577 6.105
R35097 S.n16581 S.n16580 6.105
R35098 S.n16570 S.t1675 6.105
R35099 S.n16024 S.t1126 6.105
R35100 S.n16031 S.n16030 6.105
R35101 S.n16028 S.n16027 6.105
R35102 S.n16021 S.t2149 6.105
R35103 S.n15649 S.t2943 6.105
R35104 S.n15654 S.n15653 6.105
R35105 S.n15657 S.n15656 6.105
R35106 S.n15646 S.t1632 6.105
R35107 S.n15049 S.t1614 6.105
R35108 S.n13734 S.t2751 6.105
R35109 S.n13742 S.n13741 6.105
R35110 S.n13745 S.n13744 6.105
R35111 S.n13737 S.t2579 6.105
R35112 S.n14142 S.t3981 6.105
R35113 S.n14149 S.n14148 6.105
R35114 S.n14146 S.n14145 6.105
R35115 S.n14139 S.t1782 6.105
R35116 S.n22909 S.t2939 6.105
R35117 S.n22525 S.t147 6.105
R35118 S.n22530 S.n22529 6.105
R35119 S.n22533 S.n22532 6.105
R35120 S.n22522 S.t1963 6.105
R35121 S.n22113 S.t2967 6.105
R35122 S.n22120 S.n22119 6.105
R35123 S.n22117 S.n22116 6.105
R35124 S.n22110 S.t3904 6.105
R35125 S.n21502 S.t304 6.105
R35126 S.n21507 S.n21506 6.105
R35127 S.n21510 S.n21509 6.105
R35128 S.n21499 S.t3485 6.105
R35129 S.n21835 S.t4265 6.105
R35130 S.n21839 S.n21838 6.105
R35131 S.n21842 S.n21841 6.105
R35132 S.n21832 S.t769 6.105
R35133 S.n20679 S.t256 6.105
R35134 S.n20684 S.n20683 6.105
R35135 S.n20687 S.n20686 6.105
R35136 S.n20676 S.t3438 6.105
R35137 S.n21025 S.t4214 6.105
R35138 S.n21029 S.n21028 6.105
R35139 S.n21032 S.n21031 6.105
R35140 S.n21022 S.t718 6.105
R35141 S.n20068 S.t210 6.105
R35142 S.n20073 S.n20072 6.105
R35143 S.n20076 S.n20075 6.105
R35144 S.n20065 S.t3396 6.105
R35145 S.n19621 S.t4163 6.105
R35146 S.n19628 S.n19627 6.105
R35147 S.n19625 S.n19624 6.105
R35148 S.n19618 S.t670 6.105
R35149 S.n19214 S.t151 6.105
R35150 S.n19219 S.n19218 6.105
R35151 S.n19222 S.n19221 6.105
R35152 S.n19211 S.t3352 6.105
R35153 S.n18749 S.t2593 6.105
R35154 S.n18756 S.n18755 6.105
R35155 S.n18753 S.n18752 6.105
R35156 S.n18746 S.t625 6.105
R35157 S.n18348 S.t80 6.105
R35158 S.n18353 S.n18352 6.105
R35159 S.n18356 S.n18355 6.105
R35160 S.n18345 S.t3312 6.105
R35161 S.n17866 S.t2786 6.105
R35162 S.n17873 S.n17872 6.105
R35163 S.n17870 S.n17869 6.105
R35164 S.n17863 S.t3784 6.105
R35165 S.n17459 S.t4604 6.105
R35166 S.n17464 S.n17463 6.105
R35167 S.n17467 S.n17466 6.105
R35168 S.n17456 S.t3270 6.105
R35169 S.n16957 S.t2734 6.105
R35170 S.n16964 S.n16963 6.105
R35171 S.n16961 S.n16960 6.105
R35172 S.n16954 S.t3743 6.105
R35173 S.n16557 S.t4552 6.105
R35174 S.n16562 S.n16561 6.105
R35175 S.n16565 S.n16564 6.105
R35176 S.n16554 S.t3229 6.105
R35177 S.n16039 S.t2685 6.105
R35178 S.n16046 S.n16045 6.105
R35179 S.n16043 S.n16042 6.105
R35180 S.n16036 S.t3696 6.105
R35181 S.n15633 S.t4500 6.105
R35182 S.n15638 S.n15637 6.105
R35183 S.n15641 S.n15640 6.105
R35184 S.n15630 S.t3183 6.105
R35185 S.n15095 S.t2638 6.105
R35186 S.n15102 S.n15101 6.105
R35187 S.n15099 S.n15098 6.105
R35188 S.n15092 S.t3646 6.105
R35189 S.n14696 S.t4447 6.105
R35190 S.n14701 S.n14700 6.105
R35191 S.n14704 S.n14703 6.105
R35192 S.n14693 S.t3140 6.105
R35193 S.n14111 S.t3121 6.105
R35194 S.n12746 S.t726 6.105
R35195 S.n12754 S.n12753 6.105
R35196 S.n12757 S.n12756 6.105
R35197 S.n12749 S.t617 6.105
R35198 S.n13178 S.t1938 6.105
R35199 S.n13185 S.n13184 6.105
R35200 S.n13182 S.n13181 6.105
R35201 S.n13175 S.t4184 6.105
R35202 S.n22902 S.t4495 6.105
R35203 S.n22509 S.t1503 6.105
R35204 S.n22514 S.n22513 6.105
R35205 S.n22517 S.n22516 6.105
R35206 S.n22506 S.t3512 6.105
R35207 S.n22128 S.t4527 6.105
R35208 S.n22135 S.n22134 6.105
R35209 S.n22132 S.n22131 6.105
R35210 S.n22125 S.t940 6.105
R35211 S.n21486 S.t2639 6.105
R35212 S.n21491 S.n21490 6.105
R35213 S.n21494 S.n21493 6.105
R35214 S.n21483 S.t2959 6.105
R35215 S.n21820 S.t3822 6.105
R35216 S.n21824 S.n21823 6.105
R35217 S.n21827 S.n21826 6.105
R35218 S.n21817 S.t253 6.105
R35219 S.n20663 S.t1824 6.105
R35220 S.n20668 S.n20667 6.105
R35221 S.n20671 S.n20670 6.105
R35222 S.n20660 S.t478 6.105
R35223 S.n21010 S.t1262 6.105
R35224 S.n21014 S.n21013 6.105
R35225 S.n21017 S.n21016 6.105
R35226 S.n21007 S.t2282 6.105
R35227 S.n20052 S.t1777 6.105
R35228 S.n20057 S.n20056 6.105
R35229 S.n20060 S.n20059 6.105
R35230 S.n20049 S.t436 6.105
R35231 S.n19636 S.t1210 6.105
R35232 S.n19643 S.n19642 6.105
R35233 S.n19640 S.n19639 6.105
R35234 S.n19633 S.t2233 6.105
R35235 S.n19198 S.t1728 6.105
R35236 S.n19203 S.n19202 6.105
R35237 S.n19206 S.n19205 6.105
R35238 S.n19195 S.t383 6.105
R35239 S.n18764 S.t4140 6.105
R35240 S.n18771 S.n18770 6.105
R35241 S.n18768 S.n18767 6.105
R35242 S.n18761 S.t2185 6.105
R35243 S.n18332 S.t1689 6.105
R35244 S.n18337 S.n18336 6.105
R35245 S.n18340 S.n18339 6.105
R35246 S.n18329 S.t345 6.105
R35247 S.n17881 S.t4094 6.105
R35248 S.n17888 S.n17887 6.105
R35249 S.n17885 S.n17884 6.105
R35250 S.n17878 S.t596 6.105
R35251 S.n17443 S.t1650 6.105
R35252 S.n17448 S.n17447 6.105
R35253 S.n17451 S.n17450 6.105
R35254 S.n17440 S.t300 6.105
R35255 S.n16972 S.t4292 6.105
R35256 S.n16979 S.n16978 6.105
R35257 S.n16976 S.n16975 6.105
R35258 S.n16969 S.t788 6.105
R35259 S.n16541 S.t1597 6.105
R35260 S.n16546 S.n16545 6.105
R35261 S.n16549 S.n16548 6.105
R35262 S.n16538 S.t251 6.105
R35263 S.n16054 S.t4236 6.105
R35264 S.n16061 S.n16060 6.105
R35265 S.n16058 S.n16057 6.105
R35266 S.n16051 S.t740 6.105
R35267 S.n15617 S.t1551 6.105
R35268 S.n15622 S.n15621 6.105
R35269 S.n15625 S.n15624 6.105
R35270 S.n15614 S.t204 6.105
R35271 S.n15110 S.t4188 6.105
R35272 S.n15117 S.n15116 6.105
R35273 S.n15114 S.n15113 6.105
R35274 S.n15107 S.t691 6.105
R35275 S.n14680 S.t1497 6.105
R35276 S.n14685 S.n14684 6.105
R35277 S.n14688 S.n14687 6.105
R35278 S.n14677 S.t140 6.105
R35279 S.n14157 S.t517 6.105
R35280 S.n14164 S.n14163 6.105
R35281 S.n14161 S.n14160 6.105
R35282 S.n14154 S.t1498 6.105
R35283 S.n13721 S.t783 6.105
R35284 S.n13726 S.n13725 6.105
R35285 S.n13729 S.n13728 6.105
R35286 S.n13718 S.t3939 6.105
R35287 S.n13147 S.t38 6.105
R35288 S.n11736 S.t3179 6.105
R35289 S.n11744 S.n11743 6.105
R35290 S.n11747 S.n11746 6.105
R35291 S.n11739 S.t3124 6.105
R35292 S.n12205 S.t4367 6.105
R35293 S.n12212 S.n12211 6.105
R35294 S.n12209 S.n12208 6.105
R35295 S.n12202 S.t2176 6.105
R35296 S.n22895 S.t1546 6.105
R35297 S.n22493 S.t3057 6.105
R35298 S.n22498 S.n22497 6.105
R35299 S.n22501 S.n22500 6.105
R35300 S.n22490 S.t557 6.105
R35301 S.n22143 S.t1574 6.105
R35302 S.n22150 S.n22149 6.105
R35303 S.n22147 S.n22146 6.105
R35304 S.n22140 S.t2489 6.105
R35305 S.n21470 S.t3979 6.105
R35306 S.n21475 S.n21474 6.105
R35307 S.n21478 S.n21477 6.105
R35308 S.n21467 S.t4517 6.105
R35309 S.n21805 S.t862 6.105
R35310 S.n21809 S.n21808 6.105
R35311 S.n21812 S.n21811 6.105
R35312 S.n21802 S.t1822 6.105
R35313 S.n20647 S.t3203 6.105
R35314 S.n20652 S.n20651 6.105
R35315 S.n20655 S.n20654 6.105
R35316 S.n20644 S.t3464 6.105
R35317 S.n20995 S.t4305 6.105
R35318 S.n20999 S.n20998 6.105
R35319 S.n21002 S.n21001 6.105
R35320 S.n20992 S.t787 6.105
R35321 S.n20036 S.t3326 6.105
R35322 S.n20041 S.n20040 6.105
R35323 S.n20044 S.n20043 6.105
R35324 S.n20033 S.t1993 6.105
R35325 S.n19651 S.t2774 6.105
R35326 S.n19658 S.n19657 6.105
R35327 S.n19655 S.n19654 6.105
R35328 S.n19648 S.t3778 6.105
R35329 S.n19182 S.t3279 6.105
R35330 S.n19187 S.n19186 6.105
R35331 S.n19190 S.n19189 6.105
R35332 S.n19179 S.t1945 6.105
R35333 S.n18779 S.t1185 6.105
R35334 S.n18786 S.n18785 6.105
R35335 S.n18783 S.n18782 6.105
R35336 S.n18776 S.t3732 6.105
R35337 S.n18316 S.t3240 6.105
R35338 S.n18321 S.n18320 6.105
R35339 S.n18324 S.n18323 6.105
R35340 S.n18313 S.t1903 6.105
R35341 S.n17896 S.t1137 6.105
R35342 S.n17903 S.n17902 6.105
R35343 S.n17900 S.n17899 6.105
R35344 S.n17893 S.t2158 6.105
R35345 S.n17427 S.t3199 6.105
R35346 S.n17432 S.n17431 6.105
R35347 S.n17435 S.n17434 6.105
R35348 S.n17424 S.t1860 6.105
R35349 S.n16987 S.t1091 6.105
R35350 S.n16994 S.n16993 6.105
R35351 S.n16991 S.n16990 6.105
R35352 S.n16984 S.t2110 6.105
R35353 S.n16525 S.t3155 6.105
R35354 S.n16530 S.n16529 6.105
R35355 S.n16533 S.n16532 6.105
R35356 S.n16522 S.t1819 6.105
R35357 S.n16069 S.t1286 6.105
R35358 S.n16076 S.n16075 6.105
R35359 S.n16073 S.n16072 6.105
R35360 S.n16066 S.t2300 6.105
R35361 S.n15601 S.t3104 6.105
R35362 S.n15606 S.n15605 6.105
R35363 S.n15609 S.n15608 6.105
R35364 S.n15598 S.t1769 6.105
R35365 S.n15125 S.t1235 6.105
R35366 S.n15132 S.n15131 6.105
R35367 S.n15129 S.n15128 6.105
R35368 S.n15122 S.t2247 6.105
R35369 S.n14664 S.t3050 6.105
R35370 S.n14669 S.n14668 6.105
R35371 S.n14672 S.n14671 6.105
R35372 S.n14661 S.t1725 6.105
R35373 S.n14172 S.t2083 6.105
R35374 S.n14179 S.n14178 6.105
R35375 S.n14176 S.n14175 6.105
R35376 S.n14169 S.t3051 6.105
R35377 S.n13705 S.t2335 6.105
R35378 S.n13710 S.n13709 6.105
R35379 S.n13713 S.n13712 6.105
R35380 S.n13702 S.t975 6.105
R35381 S.n13193 S.t2030 6.105
R35382 S.n13200 S.n13199 6.105
R35383 S.n13197 S.n13196 6.105
R35384 S.n13190 S.t3002 6.105
R35385 S.n12733 S.t2291 6.105
R35386 S.n12738 S.n12737 6.105
R35387 S.n12741 S.n12740 6.105
R35388 S.n12730 S.t932 6.105
R35389 S.n12174 S.t1624 6.105
R35390 S.n10713 S.t1057 6.105
R35391 S.n10721 S.n10720 6.105
R35392 S.n10724 S.n10723 6.105
R35393 S.n10716 S.t1063 6.105
R35394 S.n11206 S.t2336 6.105
R35395 S.n11213 S.n11212 6.105
R35396 S.n11210 S.n11209 6.105
R35397 S.n11203 S.t18 6.105
R35398 S.n22888 S.t3099 6.105
R35399 S.n22477 S.t10 6.105
R35400 S.n22482 S.n22481 6.105
R35401 S.n22485 S.n22484 6.105
R35402 S.n22474 S.t2124 6.105
R35403 S.n22158 S.t3127 6.105
R35404 S.n22165 S.n22164 6.105
R35405 S.n22162 S.n22161 6.105
R35406 S.n22155 S.t4032 6.105
R35407 S.n21454 S.t1016 6.105
R35408 S.n21459 S.n21458 6.105
R35409 S.n21462 S.n21461 6.105
R35410 S.n21451 S.t1567 6.105
R35411 S.n21790 S.t2411 6.105
R35412 S.n21794 S.n21793 6.105
R35413 S.n21797 S.n21796 6.105
R35414 S.n21787 S.t3369 6.105
R35415 S.n20631 S.t4522 6.105
R35416 S.n20636 S.n20635 6.105
R35417 S.n20639 S.n20638 6.105
R35418 S.n20628 S.t504 6.105
R35419 S.n20980 S.t1354 6.105
R35420 S.n20984 S.n20983 6.105
R35421 S.n20987 S.n20986 6.105
R35422 S.n20977 S.t2339 6.105
R35423 S.n20020 S.t3704 6.105
R35424 S.n20025 S.n20024 6.105
R35425 S.n20028 S.n20027 6.105
R35426 S.n20017 S.t3958 6.105
R35427 S.n19666 S.t325 6.105
R35428 S.n19673 S.n19672 6.105
R35429 S.n19670 S.n19669 6.105
R35430 S.n19663 S.t1254 6.105
R35431 S.n19166 S.t309 6.105
R35432 S.n19171 S.n19170 6.105
R35433 S.n19174 S.n19173 6.105
R35434 S.n19163 S.t3492 6.105
R35435 S.n18794 S.t2747 6.105
R35436 S.n18801 S.n18800 6.105
R35437 S.n18798 S.n18797 6.105
R35438 S.n18791 S.t779 6.105
R35439 S.n18300 S.t266 6.105
R35440 S.n18305 S.n18304 6.105
R35441 S.n18308 S.n18307 6.105
R35442 S.n18297 S.t3449 6.105
R35443 S.n17911 S.t2696 6.105
R35444 S.n17918 S.n17917 6.105
R35445 S.n17915 S.n17914 6.105
R35446 S.n17908 S.t3708 6.105
R35447 S.n17411 S.t219 6.105
R35448 S.n17416 S.n17415 6.105
R35449 S.n17419 S.n17418 6.105
R35450 S.n17408 S.t3402 6.105
R35451 S.n17002 S.t2652 6.105
R35452 S.n17009 S.n17008 6.105
R35453 S.n17006 S.n17005 6.105
R35454 S.n16999 S.t3661 6.105
R35455 S.n16509 S.t168 6.105
R35456 S.n16514 S.n16513 6.105
R35457 S.n16517 S.n16516 6.105
R35458 S.n16506 S.t3362 6.105
R35459 S.n16084 S.t2600 6.105
R35460 S.n16091 S.n16090 6.105
R35461 S.n16088 S.n16087 6.105
R35462 S.n16081 S.t3619 6.105
R35463 S.n15585 S.t99 6.105
R35464 S.n15590 S.n15589 6.105
R35465 S.n15593 S.n15592 6.105
R35466 S.n15582 S.t3322 6.105
R35467 S.n15140 S.t2797 6.105
R35468 S.n15147 S.n15146 6.105
R35469 S.n15144 S.n15143 6.105
R35470 S.n15137 S.t3790 6.105
R35471 S.n14648 S.t1 6.105
R35472 S.n14653 S.n14652 6.105
R35473 S.n14656 S.n14655 6.105
R35474 S.n14645 S.t3276 6.105
R35475 S.n14187 S.t3636 6.105
R35476 S.n14194 S.n14193 6.105
R35477 S.n14191 S.n14190 6.105
R35478 S.n14184 S.t3 6.105
R35479 S.n13689 S.t3873 6.105
R35480 S.n13694 S.n13693 6.105
R35481 S.n13697 S.n13696 6.105
R35482 S.n13686 S.t2523 6.105
R35483 S.n13208 S.t3582 6.105
R35484 S.n13215 S.n13214 6.105
R35485 S.n13212 S.n13211 6.105
R35486 S.n13205 S.t4559 6.105
R35487 S.n12717 S.t3829 6.105
R35488 S.n12722 S.n12721 6.105
R35489 S.n12725 S.n12724 6.105
R35490 S.n12714 S.t2482 6.105
R35491 S.n12220 S.t3528 6.105
R35492 S.n12227 S.n12226 6.105
R35493 S.n12224 S.n12223 6.105
R35494 S.n12217 S.t4507 6.105
R35495 S.n11723 S.t3786 6.105
R35496 S.n11728 S.n11727 6.105
R35497 S.n11731 S.n11730 6.105
R35498 S.n11720 S.t2441 6.105
R35499 S.n11175 S.t3135 6.105
R35500 S.n9668 S.t3541 6.105
R35501 S.n9676 S.n9675 6.105
R35502 S.n9679 S.n9678 6.105
R35503 S.n9671 S.t3617 6.105
R35504 S.n10198 S.t249 6.105
R35505 S.n10205 S.n10204 6.105
R35506 S.n10202 S.n10201 6.105
R35507 S.n10195 S.t2515 6.105
R35508 S.n22881 S.t90 6.105
R35509 S.n22461 S.t1657 6.105
R35510 S.n22466 S.n22465 6.105
R35511 S.n22469 S.n22468 6.105
R35512 S.n22458 S.t3670 6.105
R35513 S.n22173 S.t121 6.105
R35514 S.n22180 S.n22179 6.105
R35515 S.n22177 S.n22176 6.105
R35516 S.n22170 S.t1064 6.105
R35517 S.n21438 S.t2563 6.105
R35518 S.n21443 S.n21442 6.105
R35519 S.n21446 S.n21445 6.105
R35520 S.n21435 S.t3116 6.105
R35521 S.n21775 S.t3948 6.105
R35522 S.n21779 S.n21778 6.105
R35523 S.n21782 S.n21781 6.105
R35524 S.n21772 S.t405 6.105
R35525 S.n20615 S.t1571 6.105
R35526 S.n20620 S.n20619 6.105
R35527 S.n20623 S.n20622 6.105
R35528 S.n20612 S.t2069 6.105
R35529 S.n20965 S.t2919 6.105
R35530 S.n20969 S.n20968 6.105
R35531 S.n20972 S.n20971 6.105
R35532 S.n20962 S.t3875 6.105
R35533 S.n20004 S.t507 6.105
R35534 S.n20009 S.n20008 6.105
R35535 S.n20012 S.n20011 6.105
R35536 S.n20001 S.t995 6.105
R35537 S.n19681 S.t1887 6.105
R35538 S.n19688 S.n19687 6.105
R35539 S.n19685 S.n19684 6.105
R35540 S.n19678 S.t2819 6.105
R35541 S.n19150 S.t4167 6.105
R35542 S.n19155 S.n19154 6.105
R35543 S.n19158 S.n19157 6.105
R35544 S.n19147 S.t4492 6.105
R35545 S.n18809 S.t1333 6.105
R35546 S.n18816 S.n18815 6.105
R35547 S.n18813 S.n18812 6.105
R35548 S.n18806 S.t1801 6.105
R35549 S.n18284 S.t1829 6.105
R35550 S.n18289 S.n18288 6.105
R35551 S.n18292 S.n18291 6.105
R35552 S.n18281 S.t490 6.105
R35553 S.n17926 S.t4250 6.105
R35554 S.n17933 S.n17932 6.105
R35555 S.n17930 S.n17929 6.105
R35556 S.n17923 S.t747 6.105
R35557 S.n17395 S.t1783 6.105
R35558 S.n17400 S.n17399 6.105
R35559 S.n17403 S.n17402 6.105
R35560 S.n17392 S.t448 6.105
R35561 S.n17017 S.t4202 6.105
R35562 S.n17024 S.n17023 6.105
R35563 S.n17021 S.n17020 6.105
R35564 S.n17014 S.t704 6.105
R35565 S.n16493 S.t1739 6.105
R35566 S.n16498 S.n16497 6.105
R35567 S.n16501 S.n16500 6.105
R35568 S.n16490 S.t400 6.105
R35569 S.n16099 S.t4149 6.105
R35570 S.n16106 S.n16105 6.105
R35571 S.n16103 S.n16102 6.105
R35572 S.n16096 S.t663 6.105
R35573 S.n15569 S.t1699 6.105
R35574 S.n15574 S.n15573 6.105
R35575 S.n15577 S.n15576 6.105
R35576 S.n15566 S.t351 6.105
R35577 S.n15155 S.t4101 6.105
R35578 S.n15162 S.n15161 6.105
R35579 S.n15159 S.n15158 6.105
R35580 S.n15152 S.t610 6.105
R35581 S.n14632 S.t1654 6.105
R35582 S.n14637 S.n14636 6.105
R35583 S.n14640 S.n14639 6.105
R35584 S.n14629 S.t307 6.105
R35585 S.n14202 S.t675 6.105
R35586 S.n14209 S.n14208 6.105
R35587 S.n14206 S.n14205 6.105
R35588 S.n14199 S.t1653 6.105
R35589 S.n13673 S.t910 6.105
R35590 S.n13678 S.n13677 6.105
R35591 S.n13681 S.n13680 6.105
R35592 S.n13670 S.t4063 6.105
R35593 S.n13223 S.t631 6.105
R35594 S.n13230 S.n13229 6.105
R35595 S.n13227 S.n13226 6.105
R35596 S.n13220 S.t1601 6.105
R35597 S.n12701 S.t868 6.105
R35598 S.n12706 S.n12705 6.105
R35599 S.n12709 S.n12708 6.105
R35600 S.n12698 S.t4023 6.105
R35601 S.n12235 S.t576 6.105
R35602 S.n12242 S.n12241 6.105
R35603 S.n12239 S.n12238 6.105
R35604 S.n12232 S.t1560 6.105
R35605 S.n11707 S.t823 6.105
R35606 S.n11712 S.n11711 6.105
R35607 S.n11715 S.n11714 6.105
R35608 S.n11704 S.t3983 6.105
R35609 S.n11221 S.t526 6.105
R35610 S.n11228 S.n11227 6.105
R35611 S.n11225 S.n11224 6.105
R35612 S.n11218 S.t1509 6.105
R35613 S.n10700 S.t791 6.105
R35614 S.n10705 S.n10704 6.105
R35615 S.n10708 S.n10707 6.105
R35616 S.n10697 S.t3947 6.105
R35617 S.n10167 S.t59 6.105
R35618 S.n8610 S.t1483 6.105
R35619 S.n8618 S.n8617 6.105
R35620 S.n8621 S.n8620 6.105
R35621 S.n8613 S.t1615 6.105
R35622 S.n9164 S.t3837 6.105
R35623 S.n9171 S.n9170 6.105
R35624 S.n9168 S.n9167 6.105
R35625 S.n9161 S.t466 6.105
R35626 S.n22874 S.t1453 6.105
R35627 S.n22445 S.t3207 6.105
R35628 S.n22450 S.n22449 6.105
R35629 S.n22453 S.n22452 6.105
R35630 S.n22442 S.t712 6.105
R35631 S.n22188 S.t1714 6.105
R35632 S.n22195 S.n22194 6.105
R35633 S.n22192 S.n22191 6.105
R35634 S.n22185 S.t2617 6.105
R35635 S.n21422 S.t4103 6.105
R35636 S.n21427 S.n21426 6.105
R35637 S.n21430 S.n21429 6.105
R35638 S.n21419 S.t112 6.105
R35639 S.n21760 S.t985 6.105
R35640 S.n21764 S.n21763 6.105
R35641 S.n21767 S.n21766 6.105
R35642 S.n21757 S.t1959 6.105
R35643 S.n20599 S.t3123 6.105
R35644 S.n20604 S.n20603 6.105
R35645 S.n20607 S.n20606 6.105
R35646 S.n20596 S.t3624 6.105
R35647 S.n20950 S.t4473 6.105
R35648 S.n20954 S.n20953 6.105
R35649 S.n20957 S.n20956 6.105
R35650 S.n20947 S.t912 6.105
R35651 S.n19988 S.t2072 6.105
R35652 S.n19993 S.n19992 6.105
R35653 S.n19996 S.n19995 6.105
R35654 S.n19985 S.t2542 6.105
R35655 S.n19696 S.t3431 6.105
R35656 S.n19703 S.n19702 6.105
R35657 S.n19700 S.n19699 6.105
R35658 S.n19693 S.t4369 6.105
R35659 S.n19134 S.t1000 6.105
R35660 S.n19139 S.n19138 6.105
R35661 S.n19142 S.n19141 6.105
R35662 S.n19131 S.t1545 6.105
R35663 S.n18824 S.t2900 6.105
R35664 S.n18831 S.n18830 6.105
R35665 S.n18828 S.n18827 6.105
R35666 S.n18821 S.t3347 6.105
R35667 S.n18268 S.t202 6.105
R35668 S.n18273 S.n18272 6.105
R35669 S.n18276 S.n18275 6.105
R35670 S.n18265 S.t485 6.105
R35671 S.n17941 S.t1869 6.105
R35672 S.n17948 S.n17947 6.105
R35673 S.n17945 S.n17944 6.105
R35674 S.n17938 S.t2789 6.105
R35675 S.n17379 S.t3331 6.105
R35676 S.n17384 S.n17383 6.105
R35677 S.n17387 S.n17386 6.105
R35678 S.n17376 S.t2004 6.105
R35679 S.n17032 S.t1251 6.105
R35680 S.n17039 S.n17038 6.105
R35681 S.n17036 S.n17035 6.105
R35682 S.n17029 S.t2262 6.105
R35683 S.n16477 S.t3286 6.105
R35684 S.n16482 S.n16481 6.105
R35685 S.n16485 S.n16484 6.105
R35686 S.n16474 S.t1957 6.105
R35687 S.n16114 S.t1195 6.105
R35688 S.n16121 S.n16120 6.105
R35689 S.n16118 S.n16117 6.105
R35690 S.n16111 S.t2222 6.105
R35691 S.n15553 S.t3254 6.105
R35692 S.n15558 S.n15557 6.105
R35693 S.n15561 S.n15560 6.105
R35694 S.n15550 S.t1911 6.105
R35695 S.n15170 S.t1148 6.105
R35696 S.n15177 S.n15176 6.105
R35697 S.n15174 S.n15173 6.105
R35698 S.n15167 S.t2174 6.105
R35699 S.n14616 S.t3204 6.105
R35700 S.n14621 S.n14620 6.105
R35701 S.n14624 S.n14623 6.105
R35702 S.n14613 S.t1867 6.105
R35703 S.n14217 S.t1996 6.105
R35704 S.n14224 S.n14223 6.105
R35705 S.n14221 S.n14220 6.105
R35706 S.n14214 S.t2966 6.105
R35707 S.n13657 S.t2455 6.105
R35708 S.n13662 S.n13661 6.105
R35709 S.n13665 S.n13664 6.105
R35710 S.n13654 S.t1099 6.105
R35711 S.n13238 S.t2193 6.105
R35712 S.n13245 S.n13244 6.105
R35713 S.n13242 S.n13241 6.105
R35714 S.n13235 S.t3158 6.105
R35715 S.n12685 S.t2416 6.105
R35716 S.n12690 S.n12689 6.105
R35717 S.n12693 S.n12692 6.105
R35718 S.n12682 S.t1055 6.105
R35719 S.n12250 S.t2140 6.105
R35720 S.n12257 S.n12256 6.105
R35721 S.n12254 S.n12253 6.105
R35722 S.n12247 S.t3111 6.105
R35723 S.n11691 S.t2379 6.105
R35724 S.n11696 S.n11695 6.105
R35725 S.n11699 S.n11698 6.105
R35726 S.n11688 S.t1019 6.105
R35727 S.n11236 S.t2092 6.105
R35728 S.n11243 S.n11242 6.105
R35729 S.n11240 S.n11239 6.105
R35730 S.n11233 S.t3062 6.105
R35731 S.n10684 S.t2345 6.105
R35732 S.n10689 S.n10688 6.105
R35733 S.n10692 S.n10691 6.105
R35734 S.n10681 S.t983 6.105
R35735 S.n10213 S.t2040 6.105
R35736 S.n10220 S.n10219 6.105
R35737 S.n10217 S.n10216 6.105
R35738 S.n10210 S.t3013 6.105
R35739 S.n9655 S.t2304 6.105
R35740 S.n9660 S.n9659 6.105
R35741 S.n9663 S.n9662 6.105
R35742 S.n9652 S.t939 6.105
R35743 S.n9133 S.t6 6.105
R35744 S.n7530 S.t3911 6.105
R35745 S.n7538 S.n7537 6.105
R35746 S.n7541 S.n7540 6.105
R35747 S.n7533 S.t4064 6.105
R35748 S.n8121 S.t1776 6.105
R35749 S.n8128 S.n8127 6.105
R35750 S.n8125 S.n8124 6.105
R35751 S.n8118 S.t4021 6.105
R35752 S.n22867 S.t3014 6.105
R35753 S.n22429 S.t229 6.105
R35754 S.n22434 S.n22433 6.105
R35755 S.n22437 S.n22436 6.105
R35756 S.n22426 S.t2272 6.105
R35757 S.n22203 S.t3042 6.105
R35758 S.n22210 S.n22209 6.105
R35759 S.n22207 S.n22206 6.105
R35760 S.n22200 S.t3964 6.105
R35761 S.n21406 S.t1150 6.105
R35762 S.n21411 S.n21410 6.105
R35763 S.n21414 S.n21413 6.105
R35764 S.n21403 S.t1707 6.105
R35765 S.n21745 S.t2533 6.105
R35766 S.n21749 S.n21748 6.105
R35767 S.n21752 S.n21751 6.105
R35768 S.n21742 S.t3507 6.105
R35769 S.n20583 S.t120 6.105
R35770 S.n20588 S.n20587 6.105
R35771 S.n20591 S.n20590 6.105
R35772 S.n20580 S.t666 6.105
R35773 S.n20935 S.t1529 6.105
R35774 S.n20939 S.n20938 6.105
R35775 S.n20942 S.n20941 6.105
R35776 S.n20932 S.t2456 6.105
R35777 S.n19972 S.t3627 6.105
R35778 S.n19977 S.n19976 6.105
R35779 S.n19980 S.n19979 6.105
R35780 S.n19969 S.t4085 6.105
R35781 S.n19711 S.t470 6.105
R35782 S.n19718 S.n19717 6.105
R35783 S.n19715 S.n19714 6.105
R35784 S.n19708 S.t1424 6.105
R35785 S.n19118 S.t2545 6.105
R35786 S.n19123 S.n19122 6.105
R35787 S.n19126 S.n19125 6.105
R35788 S.n19115 S.t3098 6.105
R35789 S.n18839 S.t4456 6.105
R35790 S.n18846 S.n18845 6.105
R35791 S.n18843 S.n18842 6.105
R35792 S.n18836 S.t380 6.105
R35793 S.n18252 S.t1554 6.105
R35794 S.n18257 S.n18256 6.105
R35795 S.n18260 S.n18259 6.105
R35796 S.n18249 S.t2048 6.105
R35797 S.n17956 S.t3413 6.105
R35798 S.n17963 S.n17962 6.105
R35799 S.n17960 S.n17959 6.105
R35800 S.n17953 S.t4349 6.105
R35801 S.n17363 S.t729 6.105
R35802 S.n17368 S.n17367 6.105
R35803 S.n17371 S.n17370 6.105
R35804 S.n17360 S.t981 6.105
R35805 S.n17047 S.t2377 6.105
R35806 S.n17054 S.n17053 6.105
R35807 S.n17051 S.n17050 6.105
R35808 S.n17044 S.t3329 6.105
R35809 S.n16461 S.t317 6.105
R35810 S.n16466 S.n16465 6.105
R35811 S.n16469 S.n16468 6.105
R35812 S.n16458 S.t3503 6.105
R35813 S.n16129 S.t2758 6.105
R35814 S.n16136 S.n16135 6.105
R35815 S.n16133 S.n16132 6.105
R35816 S.n16126 S.t3765 6.105
R35817 S.n15537 S.t277 6.105
R35818 S.n15542 S.n15541 6.105
R35819 S.n15545 S.n15544 6.105
R35820 S.n15534 S.t3456 6.105
R35821 S.n15185 S.t2706 6.105
R35822 S.n15192 S.n15191 6.105
R35823 S.n15189 S.n15188 6.105
R35824 S.n15182 S.t3716 6.105
R35825 S.n14600 S.t226 6.105
R35826 S.n14605 S.n14604 6.105
R35827 S.n14608 S.n14607 6.105
R35828 S.n14597 S.t3411 6.105
R35829 S.n14232 S.t3545 6.105
R35830 S.n14239 S.n14238 6.105
R35831 S.n14236 S.n14235 6.105
R35832 S.n14229 S.t4525 6.105
R35833 S.n13641 S.t3995 6.105
R35834 S.n13646 S.n13645 6.105
R35835 S.n13649 S.n13648 6.105
R35836 S.n13638 S.t2661 6.105
R35837 S.n13253 S.t3494 6.105
R35838 S.n13260 S.n13259 6.105
R35839 S.n13257 S.n13256 6.105
R35840 S.n13250 S.t4468 6.105
R35841 S.n12669 S.t3954 6.105
R35842 S.n12674 S.n12673 6.105
R35843 S.n12677 S.n12676 6.105
R35844 S.n12666 S.t2608 6.105
R35845 S.n12265 S.t3685 6.105
R35846 S.n12272 S.n12271 6.105
R35847 S.n12269 S.n12268 6.105
R35848 S.n12262 S.t108 6.105
R35849 S.n11675 S.t3915 6.105
R35850 S.n11680 S.n11679 6.105
R35851 S.n11683 S.n11682 6.105
R35852 S.n11672 S.t2565 6.105
R35853 S.n11251 S.t3643 6.105
R35854 S.n11258 S.n11257 6.105
R35855 S.n11255 S.n11254 6.105
R35856 S.n11248 S.t17 6.105
R35857 S.n10668 S.t3880 6.105
R35858 S.n10673 S.n10672 6.105
R35859 S.n10676 S.n10675 6.105
R35860 S.n10665 S.t2528 6.105
R35861 S.n10228 S.t3595 6.105
R35862 S.n10235 S.n10234 6.105
R35863 S.n10232 S.n10231 6.105
R35864 S.n10225 S.t4570 6.105
R35865 S.n9639 S.t3839 6.105
R35866 S.n9644 S.n9643 6.105
R35867 S.n9647 S.n9646 6.105
R35868 S.n9636 S.t2488 6.105
R35869 S.n9179 S.t2018 6.105
R35870 S.n9186 S.n9185 6.105
R35871 S.n9183 S.n9182 6.105
R35872 S.n9176 S.t4521 6.105
R35873 S.n8597 S.t3795 6.105
R35874 S.n8602 S.n8601 6.105
R35875 S.n8605 S.n8604 6.105
R35876 S.n8594 S.t2452 6.105
R35877 S.n8090 S.t1603 6.105
R35878 S.n6437 S.t1865 6.105
R35879 S.n6445 S.n6444 6.105
R35880 S.n6448 S.n6447 6.105
R35881 S.n6440 S.t2108 6.105
R35882 S.n7052 S.t4175 6.105
R35883 S.n7059 S.n7058 6.105
R35884 S.n7056 S.n7055 6.105
R35885 S.n7049 S.t1983 6.105
R35886 S.n22860 S.t4573 6.105
R35887 S.n22413 S.t1795 6.105
R35888 S.n22418 S.n22417 6.105
R35889 S.n22421 S.n22420 6.105
R35890 S.n22410 S.t3813 6.105
R35891 S.n22218 S.t4599 6.105
R35892 S.n22225 S.n22224 6.105
R35893 S.n22222 S.n22221 6.105
R35894 S.n22215 S.t999 6.105
R35895 S.n21390 S.t2709 6.105
R35896 S.n21395 S.n21394 6.105
R35897 S.n21398 S.n21397 6.105
R35898 S.n21387 S.t3261 6.105
R35899 S.n21730 S.t3884 6.105
R35900 S.n21734 S.n21733 6.105
R35901 S.n21737 S.n21736 6.105
R35902 S.n21727 S.t323 6.105
R35903 S.n20567 S.t1712 6.105
R35904 S.n20572 S.n20571 6.105
R35905 S.n20575 S.n20574 6.105
R35906 S.n20564 S.t2226 6.105
R35907 S.n20920 S.t3083 6.105
R35908 S.n20924 S.n20923 6.105
R35909 S.n20927 S.n20926 6.105
R35910 S.n20917 S.t3999 6.105
R35911 S.n19956 S.t668 6.105
R35912 S.n19961 S.n19960 6.105
R35913 S.n19964 S.n19963 6.105
R35914 S.n19953 S.t1127 6.105
R35915 S.n19726 S.t2033 6.105
R35916 S.n19733 S.n19732 6.105
R35917 S.n19730 S.n19729 6.105
R35918 S.n19723 S.t2987 6.105
R35919 S.n19102 S.t4088 6.105
R35920 S.n19107 S.n19106 6.105
R35921 S.n19110 S.n19109 6.105
R35922 S.n19099 S.t87 6.105
R35923 S.n18854 S.t1507 6.105
R35924 S.n18861 S.n18860 6.105
R35925 S.n18858 S.n18857 6.105
R35926 S.n18851 S.t1939 6.105
R35927 S.n18236 S.t3105 6.105
R35928 S.n18241 S.n18240 6.105
R35929 S.n18244 S.n18243 6.105
R35930 S.n18233 S.t3602 6.105
R35931 S.n17971 S.t457 6.105
R35932 S.n17978 S.n17977 6.105
R35933 S.n17975 S.n17974 6.105
R35934 S.n17968 S.t1399 6.105
R35935 S.n17347 S.t2054 6.105
R35936 S.n17352 S.n17351 6.105
R35937 S.n17355 S.n17354 6.105
R35938 S.n17344 S.t2527 6.105
R35939 S.n17062 S.t3913 6.105
R35940 S.n17069 S.n17068 6.105
R35941 S.n17066 S.n17065 6.105
R35942 S.n17059 S.t363 6.105
R35943 S.n16445 S.t1194 6.105
R35944 S.n16450 S.n16449 6.105
R35945 S.n16453 S.n16452 6.105
R35946 S.n16442 S.t1524 6.105
R35947 S.n16144 S.t2880 6.105
R35948 S.n16151 S.n16150 6.105
R35949 S.n16148 S.n16147 6.105
R35950 S.n16141 S.t3841 6.105
R35951 S.n15521 S.t1840 6.105
R35952 S.n15526 S.n15525 6.105
R35953 S.n15529 S.n15528 6.105
R35954 S.n15518 S.t497 6.105
R35955 S.n15200 S.t4259 6.105
R35956 S.n15207 S.n15206 6.105
R35957 S.n15204 S.n15203 6.105
R35958 S.n15197 S.t761 6.105
R35959 S.n14584 S.t1789 6.105
R35960 S.n14589 S.n14588 6.105
R35961 S.n14592 S.n14591 6.105
R35962 S.n14581 S.t456 6.105
R35963 S.n14247 S.t591 6.105
R35964 S.n14254 S.n14253 6.105
R35965 S.n14251 S.n14250 6.105
R35966 S.n14244 S.t1573 6.105
R35967 S.n13625 S.t1030 6.105
R35968 S.n13630 S.n13629 6.105
R35969 S.n13633 S.n13632 6.105
R35970 S.n13622 S.t4208 6.105
R35971 S.n13268 S.t539 6.105
R35972 S.n13275 S.n13274 6.105
R35973 S.n13272 S.n13271 6.105
R35974 S.n13265 S.t1522 6.105
R35975 S.n12653 S.t989 6.105
R35976 S.n12658 S.n12657 6.105
R35977 S.n12661 S.n12660 6.105
R35978 S.n12650 S.t4158 6.105
R35979 S.n12280 S.t491 6.105
R35980 S.n12287 S.n12286 6.105
R35981 S.n12284 S.n12283 6.105
R35982 S.n12277 S.t1463 6.105
R35983 S.n11659 S.t952 6.105
R35984 S.n11664 S.n11663 6.105
R35985 S.n11667 S.n11666 6.105
R35986 S.n11656 S.t4107 6.105
R35987 S.n11266 S.t680 6.105
R35988 S.n11273 S.n11272 6.105
R35989 S.n11270 S.n11269 6.105
R35990 S.n11263 S.t1662 6.105
R35991 S.n10652 S.t917 6.105
R35992 S.n10657 S.n10656 6.105
R35993 S.n10660 S.n10659 6.105
R35994 S.n10649 S.t4068 6.105
R35995 S.n10243 S.t642 6.105
R35996 S.n10250 S.n10249 6.105
R35997 S.n10247 S.n10246 6.105
R35998 S.n10240 S.t1610 6.105
R35999 S.n9623 S.t876 6.105
R36000 S.n9628 S.n9627 6.105
R36001 S.n9631 S.n9630 6.105
R36002 S.n9620 S.t4031 6.105
R36003 S.n9194 S.t3566 6.105
R36004 S.n9201 S.n9200 6.105
R36005 S.n9198 S.n9197 6.105
R36006 S.n9191 S.t1569 6.105
R36007 S.n8581 S.t832 6.105
R36008 S.n8586 S.n8585 6.105
R36009 S.n8589 S.n8588 6.105
R36010 S.n8578 S.t3993 6.105
R36011 S.n8136 S.t3515 6.105
R36012 S.n8143 S.n8142 6.105
R36013 S.n8140 S.n8139 6.105
R36014 S.n8133 S.t4487 6.105
R36015 S.n7517 S.t798 6.105
R36016 S.n7522 S.n7521 6.105
R36017 S.n7525 S.n7524 6.105
R36018 S.n7514 S.t3949 6.105
R36019 S.n7021 S.t3115 6.105
R36020 S.n5321 S.t4275 6.105
R36021 S.n5329 S.n5328 6.105
R36022 S.n5332 S.n5331 6.105
R36023 S.n5324 S.t12 6.105
R36024 S.n5974 S.t2162 6.105
R36025 S.n5981 S.n5980 6.105
R36026 S.n5978 S.n5977 6.105
R36027 S.n5971 S.t4419 6.105
R36028 S.n22853 S.t3710 6.105
R36029 S.n22397 S.t3340 6.105
R36030 S.n22402 S.n22401 6.105
R36031 S.n22405 S.n22404 6.105
R36032 S.n22394 S.t855 6.105
R36033 S.n22233 S.t1645 6.105
R36034 S.n22240 S.n22239 6.105
R36035 S.n22237 S.n22236 6.105
R36036 S.n22230 S.t2547 6.105
R36037 S.n21374 S.t4264 6.105
R36038 S.n21379 S.n21378 6.105
R36039 S.n21382 S.n21381 6.105
R36040 S.n21371 S.t290 6.105
R36041 S.n21715 S.t920 6.105
R36042 S.n21719 S.n21718 6.105
R36043 S.n21722 S.n21721 6.105
R36044 S.n21712 S.t1883 6.105
R36045 S.n20551 S.t3265 6.105
R36046 S.n20556 S.n20555 6.105
R36047 S.n20559 S.n20558 6.105
R36048 S.n20548 S.t3770 6.105
R36049 S.n20905 S.t4383 6.105
R36050 S.n20909 S.n20908 6.105
R36051 S.n20912 S.n20911 6.105
R36052 S.n20902 S.t841 6.105
R36053 S.n19940 S.t2231 6.105
R36054 S.n19945 S.n19944 6.105
R36055 S.n19948 S.n19947 6.105
R36056 S.n19937 S.t2684 6.105
R36057 S.n19741 S.t3589 6.105
R36058 S.n19748 S.n19747 6.105
R36059 S.n19745 S.n19744 6.105
R36060 S.n19738 S.t4546 6.105
R36061 S.n19086 S.t1131 6.105
R36062 S.n19091 S.n19090 6.105
R36063 S.n19094 S.n19093 6.105
R36064 S.n19083 S.t1692 6.105
R36065 S.n18869 S.t3061 6.105
R36066 S.n18876 S.n18875 6.105
R36067 S.n18873 S.n18872 6.105
R36068 S.n18866 S.t3486 6.105
R36069 S.n18220 S.t94 6.105
R36070 S.n18225 S.n18224 6.105
R36071 S.n18228 S.n18227 6.105
R36072 S.n18217 S.t647 6.105
R36073 S.n17986 S.t2015 6.105
R36074 S.n17993 S.n17992 6.105
R36075 S.n17990 S.n17989 6.105
R36076 S.n17983 S.t2965 6.105
R36077 S.n17331 S.t3610 6.105
R36078 S.n17336 S.n17335 6.105
R36079 S.n17339 S.n17338 6.105
R36080 S.n17328 S.t4069 6.105
R36081 S.n17077 S.t949 6.105
R36082 S.n17084 S.n17083 6.105
R36083 S.n17081 S.n17080 6.105
R36084 S.n17074 S.t1922 6.105
R36085 S.n16429 S.t2532 6.105
R36086 S.n16434 S.n16433 6.105
R36087 S.n16437 S.n16436 6.105
R36088 S.n16426 S.t3075 6.105
R36089 S.n16159 S.t4432 6.105
R36090 S.n16166 S.n16165 6.105
R36091 S.n16163 S.n16162 6.105
R36092 S.n16156 S.t878 6.105
R36093 S.n15505 S.t1750 6.105
R36094 S.n15510 S.n15509 6.105
R36095 S.n15513 S.n15512 6.105
R36096 S.n15502 S.t2027 6.105
R36097 S.n15215 S.t3394 6.105
R36098 S.n15222 S.n15221 6.105
R36099 S.n15219 S.n15218 6.105
R36100 S.n15212 S.t4327 6.105
R36101 S.n14568 S.t3336 6.105
R36102 S.n14573 S.n14572 6.105
R36103 S.n14576 S.n14575 6.105
R36104 S.n14565 S.t2014 6.105
R36105 S.n14262 S.t2155 6.105
R36106 S.n14269 S.n14268 6.105
R36107 S.n14266 S.n14265 6.105
R36108 S.n14259 S.t3125 6.105
R36109 S.n13609 S.t2581 6.105
R36110 S.n13614 S.n13613 6.105
R36111 S.n13617 S.n13616 6.105
R36112 S.n13606 S.t1258 6.105
R36113 S.n13283 S.t2106 6.105
R36114 S.n13290 S.n13289 6.105
R36115 S.n13287 S.n13286 6.105
R36116 S.n13280 S.t3071 6.105
R36117 S.n12637 S.t2538 6.105
R36118 S.n12642 S.n12641 6.105
R36119 S.n12645 S.n12644 6.105
R36120 S.n12634 S.t1204 6.105
R36121 S.n12295 S.t2056 6.105
R36122 S.n12302 S.n12301 6.105
R36123 S.n12299 S.n12298 6.105
R36124 S.n12292 S.t3021 6.105
R36125 S.n11643 S.t2500 6.105
R36126 S.n11648 S.n11647 6.105
R36127 S.n11651 S.n11650 6.105
R36128 S.n11640 S.t1154 6.105
R36129 S.n11281 S.t2006 6.105
R36130 S.n11288 S.n11287 6.105
R36131 S.n11285 S.n11284 6.105
R36132 S.n11278 S.t2978 6.105
R36133 S.n10636 S.t2461 6.105
R36134 S.n10641 S.n10640 6.105
R36135 S.n10644 S.n10643 6.105
R36136 S.n10633 S.t1107 6.105
R36137 S.n10258 S.t2200 6.105
R36138 S.n10265 S.n10264 6.105
R36139 S.n10262 S.n10261 6.105
R36140 S.n10255 S.t3166 6.105
R36141 S.n9607 S.t2423 6.105
R36142 S.n9612 S.n9611 6.105
R36143 S.n9615 S.n9614 6.105
R36144 S.n9604 S.t1062 6.105
R36145 S.n9209 S.t616 6.105
R36146 S.n9216 S.n9215 6.105
R36147 S.n9213 S.n9212 6.105
R36148 S.n9206 S.t3118 6.105
R36149 S.n8565 S.t2388 6.105
R36150 S.n8570 S.n8569 6.105
R36151 S.n8573 S.n8572 6.105
R36152 S.n8562 S.t1028 6.105
R36153 S.n8151 S.t559 6.105
R36154 S.n8158 S.n8157 6.105
R36155 S.n8155 S.n8154 6.105
R36156 S.n8148 S.t1542 6.105
R36157 S.n7501 S.t2353 6.105
R36158 S.n7506 S.n7505 6.105
R36159 S.n7509 S.n7508 6.105
R36160 S.n7498 S.t987 6.105
R36161 S.n7067 S.t509 6.105
R36162 S.n7074 S.n7073 6.105
R36163 S.n7071 S.n7070 6.105
R36164 S.n7064 S.t1491 6.105
R36165 S.n6424 S.t2307 6.105
R36166 S.n6429 S.n6428 6.105
R36167 S.n6432 S.n6431 6.105
R36168 S.n6421 S.t946 6.105
R36169 S.n5943 S.t613 6.105
R36170 S.n4192 S.t720 6.105
R36171 S.n4200 S.n4199 6.105
R36172 S.n4203 S.n4202 6.105
R36173 S.n4195 S.t3735 6.105
R36174 S.n4869 S.t3073 6.105
R36175 S.n4876 S.n4875 6.105
R36176 S.n4873 S.n4872 6.105
R36177 S.n4866 S.t840 6.105
R36178 S.n22846 S.t753 6.105
R36179 S.n22381 S.t2465 6.105
R36180 S.n22386 S.n22385 6.105
R36181 S.n22389 S.n22388 6.105
R36182 S.n22378 S.t4515 6.105
R36183 S.n22248 S.t784 6.105
R36184 S.n22255 S.n22254 6.105
R36185 S.n22252 S.n22251 6.105
R36186 S.n22245 S.t1727 6.105
R36187 S.n21358 S.t1316 6.105
R36188 S.n21363 S.n21362 6.105
R36189 S.n21366 S.n21365 6.105
R36190 S.n21355 S.t1848 6.105
R36191 S.n21700 S.t2463 6.105
R36192 S.n21704 S.n21703 6.105
R36193 S.n21707 S.n21706 6.105
R36194 S.n21697 S.t3430 6.105
R36195 S.n20535 S.t293 6.105
R36196 S.n20540 S.n20539 6.105
R36197 S.n20543 S.n20542 6.105
R36198 S.n20532 S.t811 6.105
R36199 S.n20890 S.t1436 6.105
R36200 S.n20894 S.n20893 6.105
R36201 S.n20897 S.n20896 6.105
R36202 S.n20887 S.t2394 6.105
R36203 S.n19924 S.t3773 6.105
R36204 S.n19929 S.n19928 6.105
R36205 S.n19932 S.n19931 6.105
R36206 S.n19921 S.t4235 6.105
R36207 S.n19756 S.t394 6.105
R36208 S.n19763 S.n19762 6.105
R36209 S.n19760 S.n19759 6.105
R36210 S.n19753 S.t1331 6.105
R36211 S.n19070 S.t2691 6.105
R36212 S.n19075 S.n19074 6.105
R36213 S.n19078 S.n19077 6.105
R36214 S.n19067 S.t3246 6.105
R36215 S.n18884 S.t22 6.105
R36216 S.n18891 S.n18890 6.105
R36217 S.n18888 S.n18887 6.105
R36218 S.n18881 S.t528 6.105
R36219 S.n18204 S.t1696 6.105
R36220 S.n18209 S.n18208 6.105
R36221 S.n18212 S.n18211 6.105
R36222 S.n18201 S.t2208 6.105
R36223 S.n18001 S.t3561 6.105
R36224 S.n18008 S.n18007 6.105
R36225 S.n18005 S.n18004 6.105
R36226 S.n17998 S.t4524 6.105
R36227 S.n17315 S.t657 6.105
R36228 S.n17320 S.n17319 6.105
R36229 S.n17323 S.n17322 6.105
R36230 S.n17312 S.t1105 6.105
R36231 S.n17092 S.t2501 6.105
R36232 S.n17099 S.n17098 6.105
R36233 S.n17096 S.n17095 6.105
R36234 S.n17089 S.t3469 6.105
R36235 S.n16413 S.t4073 6.105
R36236 S.n16418 S.n16417 6.105
R36237 S.n16421 S.n16420 6.105
R36238 S.n16410 S.t50 6.105
R36239 S.n16174 S.t1484 6.105
R36240 S.n16181 S.n16180 6.105
R36241 S.n16178 S.n16177 6.105
R36242 S.n16171 S.t2424 6.105
R36243 S.n15489 S.t3079 6.105
R36244 S.n15494 S.n15493 6.105
R36245 S.n15497 S.n15496 6.105
R36246 S.n15486 S.t3578 6.105
R36247 S.n15230 S.t437 6.105
R36248 S.n15237 S.n15236 6.105
R36249 S.n15234 S.n15233 6.105
R36250 S.n15227 S.t1379 6.105
R36251 S.n14552 S.t2271 6.105
R36252 S.n14557 S.n14556 6.105
R36253 S.n14560 S.n14559 6.105
R36254 S.n14549 S.t2512 6.105
R36255 S.n14277 S.t3029 6.105
R36256 S.n14284 S.n14283 6.105
R36257 S.n14281 S.n14280 6.105
R36258 S.n14274 S.t3957 6.105
R36259 S.n13593 S.t4123 6.105
R36260 S.n13598 S.n13597 6.105
R36261 S.n13601 S.n13600 6.105
R36262 S.n13590 S.t2824 6.105
R36263 S.n13298 S.t3656 6.105
R36264 S.n13305 S.n13304 6.105
R36265 S.n13302 S.n13301 6.105
R36266 S.n13295 S.t44 6.105
R36267 S.n12621 S.t4080 6.105
R36268 S.n12626 S.n12625 6.105
R36269 S.n12629 S.n12628 6.105
R36270 S.n12618 S.t2769 6.105
R36271 S.n12310 S.t3611 6.105
R36272 S.n12317 S.n12316 6.105
R36273 S.n12314 S.n12313 6.105
R36274 S.n12307 S.t4581 6.105
R36275 S.n11627 S.t4042 6.105
R36276 S.n11632 S.n11631 6.105
R36277 S.n11635 S.n11634 6.105
R36278 S.n11624 S.t2715 6.105
R36279 S.n11296 S.t3556 6.105
R36280 S.n11303 S.n11302 6.105
R36281 S.n11300 S.n11299 6.105
R36282 S.n11293 S.t4534 6.105
R36283 S.n10620 S.t4002 6.105
R36284 S.n10625 S.n10624 6.105
R36285 S.n10628 S.n10627 6.105
R36286 S.n10617 S.t2666 6.105
R36287 S.n10273 S.t3505 6.105
R36288 S.n10280 S.n10279 6.105
R36289 S.n10277 S.n10276 6.105
R36290 S.n10270 S.t4476 6.105
R36291 S.n9591 S.t3960 6.105
R36292 S.n9596 S.n9595 6.105
R36293 S.n9599 S.n9598 6.105
R36294 S.n9588 S.t2616 6.105
R36295 S.n9227 S.t2177 6.105
R36296 S.n9231 S.n9230 6.105
R36297 S.n9219 S.n9218 6.105
R36298 S.n9224 S.t113 6.105
R36299 S.n8549 S.t3928 6.105
R36300 S.n8554 S.n8553 6.105
R36301 S.n8557 S.n8556 6.105
R36302 S.n8546 S.t2577 6.105
R36303 S.n8166 S.t2127 6.105
R36304 S.n8173 S.n8172 6.105
R36305 S.n8170 S.n8169 6.105
R36306 S.n8163 S.t3096 6.105
R36307 S.n7485 S.t3890 6.105
R36308 S.n7490 S.n7489 6.105
R36309 S.n7493 S.n7492 6.105
R36310 S.n7482 S.t2536 6.105
R36311 S.n7082 S.t2074 6.105
R36312 S.n7089 S.n7088 6.105
R36313 S.n7086 S.n7085 6.105
R36314 S.n7079 S.t3048 6.105
R36315 S.n6408 S.t3844 6.105
R36316 S.n6413 S.n6412 6.105
R36317 S.n6416 S.n6415 6.105
R36318 S.n6405 S.t2497 6.105
R36319 S.n5989 S.t2022 6.105
R36320 S.n5996 S.n5995 6.105
R36321 S.n5993 S.n5992 6.105
R36322 S.n5986 S.t2995 6.105
R36323 S.n5308 S.t3804 6.105
R36324 S.n5313 S.n5312 6.105
R36325 S.n5316 S.n5315 6.105
R36326 S.n5305 S.t2458 6.105
R36327 S.n4837 S.t2122 6.105
R36328 S.n3051 S.t4256 6.105
R36329 S.n3059 S.n3058 6.105
R36330 S.n3062 S.n3061 6.105
R36331 S.n3054 S.t542 6.105
R36332 S.n3756 S.t979 6.105
R36333 S.n3764 S.n3763 6.105
R36334 S.n3761 S.n3760 6.105
R36335 S.n3753 S.t3289 6.105
R36336 S.n22839 S.t2312 6.105
R36337 S.n22670 S.t4006 6.105
R36338 S.n22667 S.n22666 6.105
R36339 S.n22664 S.n22663 6.105
R36340 S.n22268 S.t1294 6.105
R36341 S.n22263 S.t2338 6.105
R36342 S.n22680 S.n22679 6.105
R36343 S.n22677 S.n22676 6.105
R36344 S.n22260 S.t3278 6.105
R36345 S.n21683 S.t471 6.105
R36346 S.n21680 S.n21679 6.105
R36347 S.n21677 S.n21676 6.105
R36348 S.n21674 S.t965 6.105
R36349 S.n21669 S.t1640 6.105
R36350 S.n21689 S.n21688 6.105
R36351 S.n21692 S.n21691 6.105
R36352 S.n21666 S.t2543 6.105
R36353 S.n20520 S.t1854 6.105
R36354 S.n20524 S.n20523 6.105
R36355 S.n20527 S.n20526 6.105
R36356 S.n20517 S.t2367 6.105
R36357 S.n20874 S.t2997 6.105
R36358 S.n20879 S.n20878 6.105
R36359 S.n20882 S.n20881 6.105
R36360 S.n20871 S.t3933 6.105
R36361 S.n19909 S.t813 6.105
R36362 S.n19913 S.n19912 6.105
R36363 S.n19916 S.n19915 6.105
R36364 S.n19906 S.t1285 6.105
R36365 S.n19771 S.t1950 6.105
R36366 S.n19779 S.n19778 6.105
R36367 S.n19776 S.n19775 6.105
R36368 S.n19768 S.t2897 6.105
R36369 S.n19055 S.t4243 6.105
R36370 S.n19059 S.n19058 6.105
R36371 S.n19062 S.n19061 6.105
R36372 S.n19052 S.t268 6.105
R36373 S.n18899 S.t1410 6.105
R36374 S.n18907 S.n18906 6.105
R36375 S.n18904 S.n18903 6.105
R36376 S.n18896 S.t1870 6.105
R36377 S.n18189 S.t3251 6.105
R36378 S.n18193 S.n18192 6.105
R36379 S.n18196 S.n18195 6.105
R36380 S.n18186 S.t3748 6.105
R36381 S.n18016 S.t608 6.105
R36382 S.n18024 S.n18023 6.105
R36383 S.n18021 S.n18020 6.105
R36384 S.n18013 S.t1572 6.105
R36385 S.n17300 S.t2213 6.105
R36386 S.n17304 S.n17303 6.105
R36387 S.n17307 S.n17306 6.105
R36388 S.n17297 S.t2665 6.105
R36389 S.n17107 S.t4043 6.105
R36390 S.n17115 S.n17114 6.105
R36391 S.n17112 S.n17111 6.105
R36392 S.n17104 S.t510 6.105
R36393 S.n16398 S.t1113 6.105
R36394 S.n16402 S.n16401 6.105
R36395 S.n16405 S.n16404 6.105
R36396 S.n16395 S.t1674 6.105
R36397 S.n16189 S.t3041 6.105
R36398 S.n16197 S.n16196 6.105
R36399 S.n16194 S.n16193 6.105
R36400 S.n16186 S.t3963 6.105
R36401 S.n15474 S.t61 6.105
R36402 S.n15478 S.n15477 6.105
R36403 S.n15481 S.n15480 6.105
R36404 S.n15471 S.t627 6.105
R36405 S.n15245 S.t1989 6.105
R36406 S.n15253 S.n15252 6.105
R36407 S.n15250 S.n15249 6.105
R36408 S.n15242 S.t2944 6.105
R36409 S.n14537 S.t3588 6.105
R36410 S.n14541 S.n14540 6.105
R36411 S.n14544 S.n14543 6.105
R36412 S.n14534 S.t4051 6.105
R36413 S.n14292 S.t4591 6.105
R36414 S.n14300 S.n14299 6.105
R36415 S.n14297 S.n14296 6.105
R36416 S.n14289 S.t994 6.105
R36417 S.n13578 S.t2393 6.105
R36418 S.n13582 S.n13581 6.105
R36419 S.n13585 S.n13584 6.105
R36420 S.n13575 S.t2640 6.105
R36421 S.n13313 S.t3530 6.105
R36422 S.n13321 S.n13320 6.105
R36423 S.n13318 S.n13317 6.105
R36424 S.n13310 S.t4491 6.105
R36425 S.n12606 S.t1123 6.105
R36426 S.n12610 S.n12609 6.105
R36427 S.n12613 S.n12612 6.105
R36428 S.n12603 S.t4325 6.105
R36429 S.n12325 S.t656 6.105
R36430 S.n12333 S.n12332 6.105
R36431 S.n12330 S.n12329 6.105
R36432 S.n12322 S.t1627 6.105
R36433 S.n11612 S.t1077 6.105
R36434 S.n11616 S.n11615 6.105
R36435 S.n11619 S.n11618 6.105
R36436 S.n11609 S.t4270 6.105
R36437 S.n11311 S.t595 6.105
R36438 S.n11319 S.n11318 6.105
R36439 S.n11316 S.n11315 6.105
R36440 S.n11308 S.t1581 6.105
R36441 S.n10605 S.t1037 6.105
R36442 S.n10609 S.n10608 6.105
R36443 S.n10612 S.n10611 6.105
R36444 S.n10602 S.t4217 6.105
R36445 S.n10288 S.t549 6.105
R36446 S.n10296 S.n10295 6.105
R36447 S.n10293 S.n10292 6.105
R36448 S.n10285 S.t1528 6.105
R36449 S.n9576 S.t997 6.105
R36450 S.n9580 S.n9579 6.105
R36451 S.n9583 S.n9582 6.105
R36452 S.n9573 S.t4166 6.105
R36453 S.n9239 S.t3483 6.105
R36454 S.n9247 S.n9246 6.105
R36455 S.n9244 S.n9243 6.105
R36456 S.n9236 S.t1472 6.105
R36457 S.n8534 S.t957 6.105
R36458 S.n8538 S.n8537 6.105
R36459 S.n8541 S.n8540 6.105
R36460 S.n8531 S.t4120 6.105
R36461 S.n8181 S.t3673 6.105
R36462 S.n8189 S.n8188 6.105
R36463 S.n8186 S.n8185 6.105
R36464 S.n8178 S.t85 6.105
R36465 S.n7470 S.t925 6.105
R36466 S.n7474 S.n7473 6.105
R36467 S.n7477 S.n7476 6.105
R36468 S.n7467 S.t4076 6.105
R36469 S.n7097 S.t3629 6.105
R36470 S.n7105 S.n7104 6.105
R36471 S.n7102 S.n7101 6.105
R36472 S.n7094 S.t4606 6.105
R36473 S.n6393 S.t883 6.105
R36474 S.n6397 S.n6396 6.105
R36475 S.n6400 S.n6399 6.105
R36476 S.n6390 S.t4038 6.105
R36477 S.n6004 S.t3573 6.105
R36478 S.n6012 S.n6011 6.105
R36479 S.n6009 S.n6008 6.105
R36480 S.n6001 S.t4556 6.105
R36481 S.n5293 S.t842 6.105
R36482 S.n5297 S.n5296 6.105
R36483 S.n5300 S.n5299 6.105
R36484 S.n5290 S.t3997 6.105
R36485 S.n4884 S.t4009 6.105
R36486 S.n4892 S.n4891 6.105
R36487 S.n4889 S.n4888 6.105
R36488 S.n4881 S.t488 6.105
R36489 S.n4180 S.t1274 6.105
R36490 S.n4184 S.n4183 6.105
R36491 S.n4187 S.n4186 6.105
R36492 S.n4177 S.t4488 6.105
R36493 S.n3724 S.t3626 6.105
R36494 S.n1444 S.t2239 6.105
R36495 S.n1890 S.n1889 6.105
R36496 S.n1893 S.n1892 6.105
R36497 S.n1896 S.t3063 6.105
R36498 S.n2625 S.t3442 6.105
R36499 S.n2633 S.n2632 6.105
R36500 S.n2630 S.n2629 6.105
R36501 S.n2622 S.t1179 6.105
R36502 S.n22830 S.t3849 6.105
R36503 S.n22364 S.t852 6.105
R36504 S.n22370 S.n22369 6.105
R36505 S.n22373 S.n22372 6.105
R36506 S.n22361 S.t2864 6.105
R36507 S.n22688 S.t3872 6.105
R36508 S.n22699 S.n22698 6.105
R36509 S.n22696 S.n22695 6.105
R36510 S.n22685 S.t308 6.105
R36511 S.n21652 S.t2034 6.105
R36512 S.n21649 S.n21648 6.105
R36513 S.n21646 S.n21645 6.105
R36514 S.n21279 S.t2325 6.105
R36515 S.n21274 S.t3193 6.105
R36516 S.n21658 S.n21657 6.105
R36517 S.n21661 S.n21660 6.105
R36518 S.n21271 S.t4086 6.105
R36519 S.n20505 S.t968 6.105
R36520 S.n20509 S.n20508 6.105
R36521 S.n20512 S.n20511 6.105
R36522 S.n20502 S.t1506 6.105
R36523 S.n20858 S.t2145 6.105
R36524 S.n20863 S.n20862 6.105
R36525 S.n20866 S.n20865 6.105
R36526 S.n20855 S.t3100 6.105
R36527 S.n19894 S.t2369 6.105
R36528 S.n19898 S.n19897 6.105
R36529 S.n19901 S.n19900 6.105
R36530 S.n19891 S.t2853 6.105
R36531 S.n19787 S.t3498 6.105
R36532 S.n19795 S.n19794 6.105
R36533 S.n19792 S.n19791 6.105
R36534 S.n19784 S.t4453 6.105
R36535 S.n19040 S.t1290 6.105
R36536 S.n19044 S.n19043 6.105
R36537 S.n19047 S.n19046 6.105
R36538 S.n19037 S.t1832 6.105
R36539 S.n18915 S.t2977 6.105
R36540 S.n18923 S.n18922 6.105
R36541 S.n18920 S.n18919 6.105
R36542 S.n18912 S.t3410 6.105
R36543 S.n18174 S.t278 6.105
R36544 S.n18178 S.n18177 6.105
R36545 S.n18181 S.n18180 6.105
R36546 S.n18171 S.t796 6.105
R36547 S.n18032 S.t1934 6.105
R36548 S.n18040 S.n18039 6.105
R36549 S.n18037 S.n18036 6.105
R36550 S.n18029 S.t2873 6.105
R36551 S.n17285 S.t3755 6.105
R36552 S.n17289 S.n17288 6.105
R36553 S.n17292 S.n17291 6.105
R36554 S.n17282 S.t4216 6.105
R36555 S.n17123 S.t1075 6.105
R36556 S.n17131 S.n17130 6.105
R36557 S.n17128 S.n17127 6.105
R36558 S.n17120 S.t2075 6.105
R36559 S.n16383 S.t2671 6.105
R36560 S.n16387 S.n16386 6.105
R36561 S.n16390 S.n16389 6.105
R36562 S.n16380 S.t3223 6.105
R36563 S.n16205 S.t4602 6.105
R36564 S.n16213 S.n16212 6.105
R36565 S.n16210 S.n16209 6.105
R36566 S.n16202 S.t1001 6.105
R36567 S.n15459 S.t1680 6.105
R36568 S.n15463 S.n15462 6.105
R36569 S.n15466 S.n15465 6.105
R36570 S.n15456 S.t2186 6.105
R36571 S.n15261 S.t3539 6.105
R36572 S.n15269 S.n15268 6.105
R36573 S.n15266 S.n15265 6.105
R36574 S.n15258 S.t4499 6.105
R36575 S.n14522 S.t632 6.105
R36576 S.n14526 S.n14525 6.105
R36577 S.n14529 S.n14528 6.105
R36578 S.n14519 S.t1087 6.105
R36579 S.n14308 S.t1634 6.105
R36580 S.n14316 S.n14315 6.105
R36581 S.n14313 S.n14312 6.105
R36582 S.n14305 S.t2541 6.105
R36583 S.n13563 S.t3727 6.105
R36584 S.n13567 S.n13566 6.105
R36585 S.n13570 S.n13569 6.105
R36586 S.n13560 S.t4186 6.105
R36587 S.n13329 S.t579 6.105
R36588 S.n13337 S.n13336 6.105
R36589 S.n13334 S.n13333 6.105
R36590 S.n13326 S.t1544 6.105
R36591 S.n12591 S.t2895 6.105
R36592 S.n12595 S.n12594 6.105
R36593 S.n12598 S.n12597 6.105
R36594 S.n12588 S.t3201 6.105
R36595 S.n12341 S.t4016 6.105
R36596 S.n12349 S.n12348 6.105
R36597 S.n12346 S.n12345 6.105
R36598 S.n12338 S.t481 6.105
R36599 S.n11597 S.t2633 6.105
R36600 S.n11601 S.n11600 6.105
R36601 S.n11604 S.n11603 6.105
R36602 S.n11594 S.t1322 6.105
R36603 S.n11327 S.t2163 6.105
R36604 S.n11335 S.n11334 6.105
R36605 S.n11332 S.n11331 6.105
R36606 S.n11324 S.t3138 6.105
R36607 S.n10590 S.t2588 6.105
R36608 S.n10594 S.n10593 6.105
R36609 S.n10597 S.n10596 6.105
R36610 S.n10587 S.t1266 6.105
R36611 S.n10304 S.t2109 6.105
R36612 S.n10312 S.n10311 6.105
R36613 S.n10309 S.n10308 6.105
R36614 S.n10301 S.t3082 6.105
R36615 S.n9561 S.t2544 6.105
R36616 S.n9565 S.n9564 6.105
R36617 S.n9568 S.n9567 6.105
R36618 S.n9558 S.t1216 6.105
R36619 S.n9255 S.t524 6.105
R36620 S.n9263 S.n9262 6.105
R36621 S.n9260 S.n9259 6.105
R36622 S.n9252 S.t3028 6.105
R36623 S.n8519 S.t2507 6.105
R36624 S.n8523 S.n8522 6.105
R36625 S.n8526 S.n8525 6.105
R36626 S.n8516 S.t1165 6.105
R36627 S.n8197 S.t474 6.105
R36628 S.n8205 S.n8204 6.105
R36629 S.n8202 S.n8201 6.105
R36630 S.n8194 S.t1449 6.105
R36631 S.n7455 S.t2467 6.105
R36632 S.n7459 S.n7458 6.105
R36633 S.n7462 S.n7461 6.105
R36634 S.n7452 S.t1118 6.105
R36635 S.n7113 S.t669 6.105
R36636 S.n7121 S.n7120 6.105
R36637 S.n7118 S.n7117 6.105
R36638 S.n7110 S.t1651 6.105
R36639 S.n6378 S.t2426 6.105
R36640 S.n6382 S.n6381 6.105
R36641 S.n6385 S.n6384 6.105
R36642 S.n6375 S.t1072 6.105
R36643 S.n6020 S.t622 6.105
R36644 S.n6028 S.n6027 6.105
R36645 S.n6025 S.n6024 6.105
R36646 S.n6017 S.t1600 6.105
R36647 S.n5278 S.t2395 6.105
R36648 S.n5282 S.n5281 6.105
R36649 S.n5285 S.n5284 6.105
R36650 S.n5275 S.t1032 6.105
R36651 S.n4900 S.t1041 6.105
R36652 S.n4908 S.n4907 6.105
R36653 S.n4905 S.n4904 6.105
R36654 S.n4897 S.t2052 6.105
R36655 S.n4165 S.t2843 6.105
R36656 S.n4169 S.n4168 6.105
R36657 S.n4172 S.n4171 6.105
R36658 S.n4162 S.t1538 6.105
R36659 S.n3772 S.t1006 6.105
R36660 S.n3780 S.n3779 6.105
R36661 S.n3777 S.n3776 6.105
R36662 S.n3769 S.t2002 6.105
R36663 S.n3039 S.t1250 6.105
R36664 S.n3043 S.n3042 6.105
R36665 S.n3046 S.n3045 6.105
R36666 S.n3036 S.t4463 6.105
R36667 S.n2593 S.t621 6.105
R36668 S.n22813 S.t4110 6.105
R36669 S.n21982 S.t605 6.105
R36670 S.n1421 S.t3548 6.105
R36671 S.n1185 S.t2390 6.105
R36672 S.n1175 S.t2884 6.105
R36673 S.n895 S.t3830 6.105
R36674 S.n919 S.n918 6.105
R36675 S.n916 S.n915 6.105
R36676 S.n898 S.t1611 6.105
R36677 S.n1977 S.t4015 6.105
R36678 S.n1987 S.n1986 6.105
R36679 S.n1990 S.n1989 6.105
R36680 S.n1974 S.t496 6.105
R36681 S.n22291 S.t3943 6.105
R36682 S.n22270 S.t1468 6.105
R36683 S.n22728 S.t2454 6.105
R36684 S.n22746 S.n22745 6.105
R36685 S.n22743 S.n22742 6.105
R36686 S.n22725 S.t3417 6.105
R36687 S.n21308 S.t395 6.105
R36688 S.n21319 S.n21318 6.105
R36689 S.n21316 S.n21315 6.105
R36690 S.n21305 S.t898 6.105
R36691 S.n21207 S.t1778 6.105
R36692 S.n21222 S.n21221 6.105
R36693 S.n21219 S.n21218 6.105
R36694 S.n21204 S.t2690 6.105
R36695 S.n20485 S.t3871 6.105
R36696 S.n20496 S.n20495 6.105
R36697 S.n20493 S.n20492 6.105
R36698 S.n20482 S.t4356 6.105
R36699 S.n20388 S.t736 6.105
R36700 S.n20403 S.n20402 6.105
R36701 S.n20400 S.n20399 6.105
R36702 S.n20385 S.t1695 6.105
R36703 S.n19874 S.t3064 6.105
R36704 S.n19885 S.n19884 6.105
R36705 S.n19882 S.n19881 6.105
R36706 S.n19871 S.t3334 6.105
R36707 S.n20261 S.t4156 6.105
R36708 S.n20273 S.n20272 6.105
R36709 S.n20276 S.n20275 6.105
R36710 S.n20258 S.t650 6.105
R36711 S.n19020 S.t2017 6.105
R36712 S.n19031 S.n19030 6.105
R36713 S.n19028 S.n19027 6.105
R36714 S.n19017 S.t2499 6.105
R36715 S.n19393 S.t3675 6.105
R36716 S.n19405 S.n19404 6.105
R36717 S.n19408 S.n19407 6.105
R36718 S.n19390 S.t4072 6.105
R36719 S.n18154 S.t3384 6.105
R36720 S.n18165 S.n18164 6.105
R36721 S.n18162 S.n18161 6.105
R36722 S.n18151 S.t3885 6.105
R36723 S.n18506 S.t519 6.105
R36724 S.n18518 S.n18517 6.105
R36725 S.n18521 S.n18520 6.105
R36726 S.n18503 S.t1477 6.105
R36727 S.n17265 S.t2356 6.105
R36728 S.n17276 S.n17275 6.105
R36729 S.n17273 S.n17272 6.105
R36730 S.n17262 S.t2832 6.105
R36731 S.n17606 S.t3975 6.105
R36732 S.n17618 S.n17617 6.105
R36733 S.n17621 S.n17620 6.105
R36734 S.n17603 S.t430 6.105
R36735 S.n16363 S.t1270 6.105
R36736 S.n16374 S.n16373 6.105
R36737 S.n16371 S.n16370 6.105
R36738 S.n16360 S.t1815 6.105
R36739 S.n16683 S.t2957 6.105
R36740 S.n16695 S.n16694 6.105
R36741 S.n16698 S.n16697 6.105
R36742 S.n16680 S.t3899 6.105
R36743 S.n15439 S.t254 6.105
R36744 S.n15450 S.n15449 6.105
R36745 S.n15447 S.n15446 6.105
R36746 S.n15436 S.t776 6.105
R36747 S.n15748 S.t2152 6.105
R36748 S.n15760 S.n15759 6.105
R36749 S.n15763 S.n15762 6.105
R36750 S.n15745 S.t3106 6.105
R36751 S.n14502 S.t3739 6.105
R36752 S.n14513 S.n14512 6.105
R36753 S.n14510 S.n14509 6.105
R36754 S.n14499 S.t4197 6.105
R36755 S.n14790 S.t206 6.105
R36756 S.n14802 S.n14801 6.105
R36757 S.n14805 S.n14804 6.105
R36758 S.n14787 S.t1125 6.105
R36759 S.n13543 S.t2327 6.105
R36760 S.n13554 S.n13553 6.105
R36761 S.n13551 S.n13550 6.105
R36762 S.n13540 S.t2795 6.105
R36763 S.n13820 S.t3689 6.105
R36764 S.n13832 S.n13831 6.105
R36765 S.n13835 S.n13834 6.105
R36766 S.n13817 S.t86 6.105
R36767 S.n12571 S.t1239 6.105
R36768 S.n12582 S.n12581 6.105
R36769 S.n12579 S.n12578 6.105
R36770 S.n12568 S.t1784 6.105
R36771 S.n12827 S.t2603 6.105
R36772 S.n12839 S.n12838 6.105
R36773 S.n12842 S.n12841 6.105
R36774 S.n12824 S.t3601 6.105
R36775 S.n11577 S.t224 6.105
R36776 S.n11588 S.n11587 6.105
R36777 S.n11585 S.n11584 6.105
R36778 S.n11574 S.t744 6.105
R36779 S.n11822 S.t1617 6.105
R36780 S.n11834 S.n11833 6.105
R36781 S.n11837 S.n11836 6.105
R36782 S.n11819 S.t2525 6.105
R36783 S.n10570 S.t3912 6.105
R36784 S.n10581 S.n10580 6.105
R36785 S.n10578 S.n10577 6.105
R36786 S.n10567 S.t4165 6.105
R36787 S.n10794 S.t560 6.105
R36788 S.n10806 S.n10805 6.105
R36789 S.n10809 S.n10808 6.105
R36790 S.n10791 S.t1523 6.105
R36791 S.n9541 S.t1130 6.105
R36792 S.n9552 S.n9551 6.105
R36793 S.n9549 S.n9548 6.105
R36794 S.n9538 S.t4331 6.105
R36795 S.n9754 S.t3641 6.105
R36796 S.n9766 S.n9765 6.105
R36797 S.n9769 S.n9768 6.105
R36798 S.n9751 S.t1637 6.105
R36799 S.n8499 S.t1084 6.105
R36800 S.n8510 S.n8509 6.105
R36801 S.n8507 S.n8506 6.105
R36802 S.n8496 S.t4282 6.105
R36803 S.n8691 S.t3592 6.105
R36804 S.n8703 S.n8702 6.105
R36805 S.n8706 S.n8705 6.105
R36806 S.n8688 S.t4569 6.105
R36807 S.n7435 S.t1040 6.105
R36808 S.n7446 S.n7445 6.105
R36809 S.n7443 S.n7442 6.105
R36810 S.n7432 S.t4226 6.105
R36811 S.n7616 S.t3536 6.105
R36812 S.n7628 S.n7627 6.105
R36813 S.n7631 S.n7630 6.105
R36814 S.n7613 S.t4519 6.105
R36815 S.n6358 S.t1005 6.105
R36816 S.n6369 S.n6368 6.105
R36817 S.n6366 S.n6365 6.105
R36818 S.n6355 S.t4176 6.105
R36819 S.n6518 S.t3487 6.105
R36820 S.n6530 S.n6529 6.105
R36821 S.n6533 S.n6532 6.105
R36822 S.n6515 S.t4461 6.105
R36823 S.n5258 S.t966 6.105
R36824 S.n5269 S.n5268 6.105
R36825 S.n5266 S.n5265 6.105
R36826 S.n5255 S.t4127 6.105
R36827 S.n5407 S.t4142 6.105
R36828 S.n5419 S.n5418 6.105
R36829 S.n5422 S.n5421 6.105
R36830 S.n5404 S.t652 6.105
R36831 S.n4145 S.t1446 6.105
R36832 S.n4156 S.n4155 6.105
R36833 S.n4153 S.n4152 6.105
R36834 S.n4142 S.t82 6.105
R36835 S.n4273 S.t4095 6.105
R36836 S.n4285 S.n4284 6.105
R36837 S.n4288 S.n4287 6.105
R36838 S.n4270 S.t598 6.105
R36839 S.n3019 S.t4366 6.105
R36840 S.n3030 S.n3029 6.105
R36841 S.n3027 S.n3026 6.105
R36842 S.n3016 S.t3069 6.105
R36843 S.n3137 S.t4057 6.105
R36844 S.n3148 S.n3147 6.105
R36845 S.n3151 S.n3150 6.105
R36846 S.n3134 S.t545 6.105
R36847 S.n1858 S.t4313 6.105
R36848 S.n1870 S.n1869 6.105
R36849 S.n1867 S.n1866 6.105
R36850 S.n1855 S.t3018 6.105
R36851 S.n873 S.t4262 6.105
R36852 S.n876 S.n875 6.105
R36853 S.n879 S.n878 6.105
R36854 S.n882 S.t2970 6.105
R36855 S.n797 S.t138 6.105
R36856 S.n808 S.n807 6.105
R36857 S.n811 S.n810 6.105
R36858 S.n800 S.t1017 6.105
R36859 S.n953 S.t2133 6.105
R36860 S.n22821 S.t888 6.105
R36861 S.n22345 S.t2404 6.105
R36862 S.n22353 S.n22352 6.105
R36863 S.n22356 S.n22355 6.105
R36864 S.n22348 S.t4418 6.105
R36865 S.n22707 S.t909 6.105
R36866 S.n22718 S.n22717 6.105
R36867 S.n22715 S.n22714 6.105
R36868 S.n22710 S.t1872 6.105
R36869 S.n21339 S.t3358 6.105
R36870 S.n21347 S.n21346 6.105
R36871 S.n21350 S.n21349 6.105
R36872 S.n21342 S.t3863 6.105
R36873 S.n21255 S.t212 6.105
R36874 S.n21263 S.n21262 6.105
R36875 S.n21266 S.n21265 6.105
R36876 S.n21258 S.t1129 6.105
R36877 S.n20433 S.t2518 6.105
R36878 S.n20826 S.n20825 6.105
R36879 S.n20829 S.n20828 6.105
R36880 S.n20832 S.t2801 6.105
R36881 S.n20839 S.t3693 6.105
R36882 S.n20847 S.n20846 6.105
R36883 S.n20850 S.n20849 6.105
R36884 S.n20842 S.t92 6.105
R36885 S.n19799 S.t1515 6.105
R36886 S.n20191 S.n20190 6.105
R36887 S.n20194 S.n20193 6.105
R36888 S.n20197 S.t2010 6.105
R36889 S.n20204 S.t2606 6.105
R36890 S.n20215 S.n20214 6.105
R36891 S.n20212 S.n20211 6.105
R36892 S.n20207 S.t3606 6.105
R36893 S.n18927 S.t2857 6.105
R36894 S.n19321 S.n19320 6.105
R36895 S.n19324 S.n19323 6.105
R36896 S.n19327 S.t3377 6.105
R36897 S.n19334 S.t4537 6.105
R36898 S.n19345 S.n19344 6.105
R36899 S.n19342 S.n19341 6.105
R36900 S.n19337 S.t454 6.105
R36901 S.n18044 S.t1842 6.105
R36902 S.n18439 S.n18438 6.105
R36903 S.n18442 S.n18441 6.105
R36904 S.n18445 S.t2350 6.105
R36905 S.n18452 S.t3481 6.105
R36906 S.n18463 S.n18462 6.105
R36907 S.n18460 S.n18459 6.105
R36908 S.n18455 S.t4428 6.105
R36909 S.n17135 S.t801 6.105
R36910 S.n17534 S.n17533 6.105
R36911 S.n17537 S.n17536 6.105
R36912 S.n17540 S.t1264 6.105
R36913 S.n17547 S.t2436 6.105
R36914 S.n17558 S.n17557 6.105
R36915 S.n17555 S.n17554 6.105
R36916 S.n17550 S.t3391 6.105
R36917 S.n16217 S.t4221 6.105
R36918 S.n16616 S.n16615 6.105
R36919 S.n16619 S.n16618 6.105
R36920 S.n16622 S.t247 6.105
R36921 S.n16629 S.t1648 6.105
R36922 S.n16640 S.n16639 6.105
R36923 S.n16637 S.n16636 6.105
R36924 S.n16632 S.t2548 6.105
R36925 S.n15273 S.t3231 6.105
R36926 S.n15676 S.n15675 6.105
R36927 S.n15679 S.n15678 6.105
R36928 S.n15682 S.t3733 6.105
R36929 S.n15689 S.t587 6.105
R36930 S.n15700 S.n15699 6.105
R36931 S.n15697 S.n15696 6.105
R36932 S.n15692 S.t1555 6.105
R36933 S.n14320 S.t2194 6.105
R36934 S.n14723 S.n14722 6.105
R36935 S.n14726 S.n14725 6.105
R36936 S.n14729 S.t2648 6.105
R36937 S.n14736 S.t3186 6.105
R36938 S.n14747 S.n14746 6.105
R36939 S.n14744 S.n14743 6.105
R36940 S.n14739 S.t4083 6.105
R36941 S.n13341 S.t772 6.105
R36942 S.n13748 S.n13747 6.105
R36943 S.n13751 S.n13750 6.105
R36944 S.n13754 S.t1233 6.105
R36945 S.n13761 S.t2143 6.105
R36946 S.n13772 S.n13771 6.105
R36947 S.n13769 S.n13768 6.105
R36948 S.n13764 S.t3097 6.105
R36949 S.n12353 S.t4192 6.105
R36950 S.n12760 S.n12759 6.105
R36951 S.n12763 S.n12762 6.105
R36952 S.n12766 S.t222 6.105
R36953 S.n12773 S.t1049 6.105
R36954 S.n12784 S.n12783 6.105
R36955 S.n12781 S.n12780 6.105
R36956 S.n12776 S.t2045 6.105
R36957 S.n11339 S.t3412 6.105
R36958 S.n11750 S.n11749 6.105
R36959 S.n11753 S.n11752 6.105
R36960 S.n11756 S.t3701 6.105
R36961 S.n11763 S.t4572 6.105
R36962 S.n11774 S.n11773 6.105
R36963 S.n11771 S.n11770 6.105
R36964 S.n11766 S.t980 6.105
R36965 S.n10316 S.t4134 6.105
R36966 S.n10727 S.n10726 6.105
R36967 S.n10730 S.n10729 6.105
R36968 S.n10733 S.t2830 6.105
R36969 S.n10740 S.t3664 6.105
R36970 S.n10751 S.n10750 6.105
R36971 S.n10748 S.n10747 6.105
R36972 S.n10743 S.t66 6.105
R36973 S.n9267 S.t4087 6.105
R36974 S.n9682 S.n9681 6.105
R36975 S.n9685 S.n9684 6.105
R36976 S.n9688 S.t2778 6.105
R36977 S.n9695 S.t2090 6.105
R36978 S.n9706 S.n9705 6.105
R36979 S.n9703 S.n9702 6.105
R36980 S.n9698 S.t4590 6.105
R36981 S.n8209 S.t4048 6.105
R36982 S.n8624 S.n8623 6.105
R36983 S.n8627 S.n8626 6.105
R36984 S.n8630 S.t2725 6.105
R36985 S.n8637 S.t2036 6.105
R36986 S.n8648 S.n8647 6.105
R36987 S.n8645 S.n8644 6.105
R36988 S.n8640 S.t3011 6.105
R36989 S.n7125 S.t4008 6.105
R36990 S.n7544 S.n7543 6.105
R36991 S.n7547 S.n7546 6.105
R36992 S.n7550 S.t2674 6.105
R36993 S.n7557 S.t1986 6.105
R36994 S.n7568 S.n7567 6.105
R36995 S.n7565 S.n7564 6.105
R36996 S.n7560 S.t2961 6.105
R36997 S.n6032 S.t3968 6.105
R36998 S.n6451 S.n6450 6.105
R36999 S.n6454 S.n6453 6.105
R37000 S.n6457 S.t2626 6.105
R37001 S.n6464 S.t2183 6.105
R37002 S.n6475 S.n6474 6.105
R37003 S.n6472 S.n6471 6.105
R37004 S.n6467 S.t3157 6.105
R37005 S.n4912 S.t3932 6.105
R37006 S.n5335 S.n5334 6.105
R37007 S.n5338 S.n5337 6.105
R37008 S.n5341 S.t2585 6.105
R37009 S.n5348 S.t2594 6.105
R37010 S.n5359 S.n5358 6.105
R37011 S.n5356 S.n5355 6.105
R37012 S.n5351 S.t3608 6.105
R37013 S.n3784 S.t4398 6.105
R37014 S.n4206 S.n4205 6.105
R37015 S.n4209 S.n4208 6.105
R37016 S.n4212 S.t3093 6.105
R37017 S.n4219 S.t2554 6.105
R37018 S.n4230 S.n4229 6.105
R37019 S.n4227 S.n4226 6.105
R37020 S.n4222 S.t3552 6.105
R37021 S.n2637 S.t2813 6.105
R37022 S.n3065 S.n3064 6.105
R37023 S.n3068 S.n3067 6.105
R37024 S.n3071 S.t1518 6.105
R37025 S.n3078 S.t2516 6.105
R37026 S.n3089 S.n3088 6.105
R37027 S.n3086 S.n3085 6.105
R37028 S.n3081 S.t3501 6.105
R37029 S.n1876 S.t2757 6.105
R37030 S.n1884 S.n1883 6.105
R37031 S.n1887 S.n1886 6.105
R37032 S.n1879 S.t1457 6.105
R37033 S.n1921 S.t1365 6.105
R37034 S.n1936 S.n1935 6.105
R37035 S.n1933 S.n1932 6.105
R37036 S.n1924 S.t3668 6.105
R37037 S.n1300 S.t1673 6.105
R37038 S.n1293 S.t2990 6.105
R37039 S.n400 S.t2493 6.105
R37040 S.n411 S.n410 6.105
R37041 S.n408 S.n407 6.105
R37042 S.n403 S.t3480 6.105
R37043 S.n2129 S.t2534 6.105
R37044 S.n2139 S.n2138 6.105
R37045 S.n2142 S.n2141 6.105
R37046 S.n2126 S.t3522 6.105
R37047 S.n18062 S.t3977 6.105
R37048 S.n18046 S.t4511 6.105
R37049 S.n18471 S.t1350 6.105
R37050 S.n18488 S.n18487 6.105
R37051 S.n18485 S.n18484 6.105
R37052 S.n18468 S.t2332 6.105
R37053 S.n17163 S.t2960 6.105
R37054 S.n17174 S.n17173 6.105
R37055 S.n17171 S.n17170 6.105
R37056 S.n17160 S.t3459 6.105
R37057 S.n17755 S.t320 6.105
R37058 S.n17767 S.n17766 6.105
R37059 S.n17770 S.n17769 6.105
R37060 S.n17752 S.t1245 6.105
R37061 S.n16263 S.t1918 6.105
R37062 S.n16274 S.n16273 6.105
R37063 S.n16271 S.n16270 6.105
R37064 S.n16260 S.t2415 6.105
R37065 S.n16828 S.t3802 6.105
R37066 S.n16840 S.n16839 6.105
R37067 S.n16843 S.n16842 6.105
R37068 S.n16825 S.t232 6.105
R37069 S.n15339 S.t1058 6.105
R37070 S.n15350 S.n15349 6.105
R37071 S.n15347 S.n15346 6.105
R37072 S.n15336 S.t1367 6.105
R37073 S.n15893 S.t2723 6.105
R37074 S.n15905 S.n15904 6.105
R37075 S.n15908 S.n15907 6.105
R37076 S.n15890 S.t3712 6.105
R37077 S.n14402 S.t4584 6.105
R37078 S.n14413 S.n14412 6.105
R37079 S.n14410 S.n14409 6.105
R37080 S.n14399 S.t566 6.105
R37081 S.n14935 S.t831 6.105
R37082 S.n14947 S.n14946 6.105
R37083 S.n14950 S.n14949 6.105
R37084 S.n14932 S.t1787 6.105
R37085 S.n13443 S.t1023 6.105
R37086 S.n13454 S.n13453 6.105
R37087 S.n13451 S.n13450 6.105
R37088 S.n13440 S.t1575 6.105
R37089 S.n13965 S.t2218 6.105
R37090 S.n13977 S.n13976 6.105
R37091 S.n13980 S.n13979 6.105
R37092 S.n13962 S.t3164 6.105
R37093 S.n12471 S.t4536 6.105
R37094 S.n12482 S.n12481 6.105
R37095 S.n12479 S.n12478 6.105
R37096 S.n12468 S.t516 6.105
R37097 S.n12972 S.t1120 6.105
R37098 S.n12984 S.n12983 6.105
R37099 S.n12987 S.n12986 6.105
R37100 S.n12969 S.t2120 6.105
R37101 S.n11477 S.t3478 6.105
R37102 S.n11488 S.n11487 6.105
R37103 S.n11485 S.n11484 6.105
R37104 S.n11474 S.t3966 6.105
R37105 S.n11967 S.t68 6.105
R37106 S.n11979 S.n11978 6.105
R37107 S.n11982 S.n11981 6.105
R37108 S.n11964 S.t1036 6.105
R37109 S.n10470 S.t2435 6.105
R37110 S.n10481 S.n10480 6.105
R37111 S.n10478 S.n10477 6.105
R37112 S.n10467 S.t2946 6.105
R37113 S.n10939 S.t3816 6.105
R37114 S.n10951 S.n10950 6.105
R37115 S.n10954 S.n10953 6.105
R37116 S.n10936 S.t246 6.105
R37117 S.n9441 S.t1389 6.105
R37118 S.n9452 S.n9451 6.105
R37119 S.n9449 S.n9448 6.105
R37120 S.n9438 S.t1910 6.105
R37121 S.n9899 S.t3283 6.105
R37122 S.n9911 S.n9910 6.105
R37123 S.n9914 S.n9913 6.105
R37124 S.n9896 S.t3728 6.105
R37125 S.n8399 S.t355 6.105
R37126 S.n8410 S.n8409 6.105
R37127 S.n8407 S.n8406 6.105
R37128 S.n8396 S.t866 6.105
R37129 S.n8836 S.t2253 6.105
R37130 S.n8848 S.n8847 6.105
R37131 S.n8851 S.n8850 6.105
R37132 S.n8833 S.t3205 6.105
R37133 S.n7335 S.t3833 6.105
R37134 S.n7346 S.n7345 6.105
R37135 S.n7343 S.n7342 6.105
R37136 S.n7332 S.t4308 6.105
R37137 S.n7761 S.t1159 6.105
R37138 S.n7773 S.n7772 6.105
R37139 S.n7776 S.n7775 6.105
R37140 S.n7758 S.t2164 6.105
R37141 S.n6258 S.t2759 6.105
R37142 S.n6269 S.n6268 6.105
R37143 S.n6266 S.n6265 6.105
R37144 S.n6255 S.t3298 6.105
R37145 S.n6663 S.t131 6.105
R37146 S.n6675 S.n6674 6.105
R37147 S.n6678 S.n6677 6.105
R37148 S.n6660 S.t1067 6.105
R37149 S.n5158 S.t1971 6.105
R37150 S.n5169 S.n5168 6.105
R37151 S.n5166 S.n5165 6.105
R37152 S.n5155 S.t2266 6.105
R37153 S.n5553 S.t1708 6.105
R37154 S.n5565 S.n5564 6.105
R37155 S.n5568 S.n5567 6.105
R37156 S.n5550 S.t2611 6.105
R37157 S.n4046 S.t177 6.105
R37158 S.n4057 S.n4056 6.105
R37159 S.n4054 S.n4053 6.105
R37160 S.n4043 S.t3375 6.105
R37161 S.n4418 S.t2614 6.105
R37162 S.n4430 S.n4429 6.105
R37163 S.n4433 S.n4432 6.105
R37164 S.n4415 S.t3630 6.105
R37165 S.n2919 S.t3142 6.105
R37166 S.n2930 S.n2929 6.105
R37167 S.n2927 S.n2926 6.105
R37168 S.n2916 S.t1805 6.105
R37169 S.n3281 S.t2575 6.105
R37170 S.n3292 S.n3291 6.105
R37171 S.n3295 S.n3294 6.105
R37172 S.n3278 S.t3575 6.105
R37173 S.n1750 S.t3091 6.105
R37174 S.n1762 S.n1761 6.105
R37175 S.n1759 S.n1758 6.105
R37176 S.n1747 S.t1760 6.105
R37177 S.n1418 S.t52 6.105
R37178 S.n1419 S.t1430 6.105
R37179 S.n12 S.t1149 6.105
R37180 S.n15 S.n14 6.105
R37181 S.n18 S.n17 6.105
R37182 S.n21 S.t2170 6.105
R37183 S.n18946 S.t3482 6.105
R37184 S.n18929 S.t3972 6.105
R37185 S.n19357 S.t858 6.105
R37186 S.n19375 S.n19374 6.105
R37187 S.n19372 S.n19371 6.105
R37188 S.n19360 S.t1268 6.105
R37189 S.n18071 S.t2437 6.105
R37190 S.n18082 S.n18081 6.105
R37191 S.n18079 S.n18078 6.105
R37192 S.n18074 S.t2954 6.105
R37193 S.n18618 S.t4297 6.105
R37194 S.n18635 S.n18634 6.105
R37195 S.n18638 S.n18637 6.105
R37196 S.n18621 S.t778 6.105
R37197 S.n17182 S.t1393 6.105
R37198 S.n17193 S.n17192 6.105
R37199 S.n17190 S.n17189 6.105
R37200 S.n17185 S.t1913 6.105
R37201 S.n17718 S.t3291 6.105
R37202 S.n17735 S.n17734 6.105
R37203 S.n17738 S.n17737 6.105
R37204 S.n17721 S.t4200 6.105
R37205 S.n16280 S.t590 6.105
R37206 S.n16291 S.n16290 6.105
R37207 S.n16288 S.n16287 6.105
R37208 S.n16283 S.t870 6.105
R37209 S.n16791 S.t2259 6.105
R37210 S.n16808 S.n16807 6.105
R37211 S.n16811 S.n16810 6.105
R37212 S.n16794 S.t3208 6.105
R37213 S.n15356 S.t4029 6.105
R37214 S.n15367 S.n15366 6.105
R37215 S.n15364 S.n15363 6.105
R37216 S.n15359 S.t4576 6.105
R37217 S.n15856 S.t1162 6.105
R37218 S.n15873 S.n15872 6.105
R37219 S.n15876 S.n15875 6.105
R37220 S.n15859 S.t2169 6.105
R37221 S.n14419 S.t911 6.105
R37222 S.n14430 S.n14429 6.105
R37223 S.n14427 S.n14426 6.105
R37224 S.n14422 S.t1416 6.105
R37225 S.n14898 S.t1700 6.105
R37226 S.n14915 S.n14914 6.105
R37227 S.n14918 S.n14917 6.105
R37228 S.n14901 S.t2599 6.105
R37229 S.n13460 S.t3991 6.105
R37230 S.n13471 S.n13470 6.105
R37231 S.n13468 S.n13467 6.105
R37232 S.n13463 S.t4528 6.105
R37233 S.n13928 S.t659 6.105
R37234 S.n13945 S.n13944 6.105
R37235 S.n13948 S.n13947 6.105
R37236 S.n13931 S.t1609 6.105
R37237 S.n12488 S.t2976 6.105
R37238 S.n12499 S.n12498 6.105
R37239 S.n12496 S.n12495 6.105
R37240 S.n12491 S.t3474 6.105
R37241 S.n12935 S.t4077 6.105
R37242 S.n12952 S.n12951 6.105
R37243 S.n12955 S.n12954 6.105
R37244 S.n12938 S.t554 6.105
R37245 S.n11494 S.t1932 6.105
R37246 S.n11505 S.n11504 6.105
R37247 S.n11502 S.n11501 6.105
R37248 S.n11497 S.t2425 6.105
R37249 S.n11930 S.t3307 6.105
R37250 S.n11947 S.n11946 6.105
R37251 S.n11950 S.n11949 6.105
R37252 S.n11933 S.t4215 6.105
R37253 S.n10487 S.t887 6.105
R37254 S.n10498 S.n10497 6.105
R37255 S.n10495 S.n10494 6.105
R37256 S.n10490 S.t1380 6.105
R37257 S.n10902 S.t2276 6.105
R37258 S.n10919 S.n10918 6.105
R37259 S.n10922 S.n10921 6.105
R37260 S.n10905 S.t3222 6.105
R37261 S.n9458 S.t4337 6.105
R37262 S.n9469 S.n9468 6.105
R37263 S.n9466 S.n9465 6.105
R37264 S.n9461 S.t350 6.105
R37265 S.n9862 S.t1735 6.105
R37266 S.n9879 S.n9878 6.105
R37267 S.n9882 S.n9881 6.105
R37268 S.n9865 S.t2184 6.105
R37269 S.n8416 S.t3324 6.105
R37270 S.n8427 S.n8426 6.105
R37271 S.n8424 S.n8423 6.105
R37272 S.n8419 S.t3825 6.105
R37273 S.n8799 S.t694 6.105
R37274 S.n8816 S.n8815 6.105
R37275 S.n8819 S.n8818 6.105
R37276 S.n8802 S.t1655 6.105
R37277 S.n7352 S.t2293 6.105
R37278 S.n7363 S.n7362 6.105
R37279 S.n7360 S.n7359 6.105
R37280 S.n7355 S.t2752 6.105
R37281 S.n7724 S.t4112 6.105
R37282 S.n7741 S.n7740 6.105
R37283 S.n7744 S.n7743 6.105
R37284 S.n7727 S.t599 6.105
R37285 S.n6275 S.t1460 6.105
R37286 S.n6286 S.n6285 6.105
R37287 S.n6283 S.n6282 6.105
R37288 S.n6278 S.t1746 6.105
R37289 S.n6626 S.t3132 6.105
R37290 S.n6643 S.n6642 6.105
R37291 S.n6646 S.n6645 6.105
R37292 S.n6629 S.t4036 6.105
R37293 S.n5175 S.t2655 6.105
R37294 S.n5186 S.n5185 6.105
R37295 S.n5183 S.n5182 6.105
R37296 S.n5178 S.t1340 6.105
R37297 S.n5516 S.t1103 6.105
R37298 S.n5533 S.n5532 6.105
R37299 S.n5536 S.n5535 6.105
R37300 S.n5519 S.t2130 6.105
R37301 S.n4063 S.t3161 6.105
R37302 S.n4074 S.n4073 6.105
R37303 S.n4071 S.n4070 6.105
R37304 S.n4066 S.t1828 6.105
R37305 S.n4381 S.t1060 6.105
R37306 S.n4398 S.n4397 6.105
R37307 S.n4401 S.n4400 6.105
R37308 S.n4384 S.t2076 6.105
R37309 S.n2936 S.t1586 6.105
R37310 S.n2947 S.n2946 6.105
R37311 S.n2944 S.n2943 6.105
R37312 S.n2939 S.t239 6.105
R37313 S.n3244 S.t1025 6.105
R37314 S.n3261 S.n3260 6.105
R37315 S.n3264 S.n3263 6.105
R37316 S.n3247 S.t2024 6.105
R37317 S.n1768 S.t1537 6.105
R37318 S.n1781 S.n1780 6.105
R37319 S.n1778 S.n1777 6.105
R37320 S.n1771 S.t190 6.105
R37321 S.n1790 S.t4483 6.105
R37322 S.n1804 S.n1803 6.105
R37323 S.n1801 S.n1800 6.105
R37324 S.n1793 S.t3173 6.105
R37325 S.n2060 S.t4151 6.105
R37326 S.n2081 S.n2080 6.105
R37327 S.n2084 S.n2083 6.105
R37328 S.n2063 S.t661 6.105
R37329 S.n415 S.t4435 6.105
R37330 S.n814 S.n813 6.105
R37331 S.n817 S.n816 6.105
R37332 S.n820 S.t3130 6.105
R37333 S.n828 S.t4102 6.105
R37334 S.n843 S.n842 6.105
R37335 S.n840 S.n839 6.105
R37336 S.n831 S.t612 6.105
R37337 S.n1315 S.t3076 6.105
R37338 S.n1307 S.t4376 6.105
R37339 S.n3221 S.t3989 6.105
R37340 S.n3232 S.n3231 6.105
R37341 S.n3235 S.n3234 6.105
R37342 S.n3218 S.t463 6.105
R37343 S.n4357 S.t4027 6.105
R37344 S.n4369 S.n4368 6.105
R37345 S.n4372 S.n4371 6.105
R37346 S.n4354 S.t511 6.105
R37347 S.n5492 S.t4065 6.105
R37348 S.n5504 S.n5503 6.105
R37349 S.n5507 S.n5506 6.105
R37350 S.n5489 S.t562 6.105
R37351 S.n6602 S.t3647 6.105
R37352 S.n6614 S.n6613 6.105
R37353 S.n6617 S.n6616 6.105
R37354 S.n6599 S.t36 6.105
R37355 S.n7700 S.t2568 6.105
R37356 S.n7712 S.n7711 6.105
R37357 S.n7715 S.n7714 6.105
R37358 S.n7697 S.t3554 6.105
R37359 S.n8775 S.t3652 6.105
R37360 S.n8787 S.n8786 6.105
R37361 S.n8790 S.n8789 6.105
R37362 S.n8772 S.t5 6.105
R37363 S.n9838 S.t161 6.105
R37364 S.n9850 S.n9849 6.105
R37365 S.n9853 S.n9852 6.105
R37366 S.n9835 S.t626 6.105
R37367 S.n10878 S.t710 6.105
R37368 S.n10890 S.n10889 6.105
R37369 S.n10893 S.n10892 6.105
R37370 S.n10875 S.t1672 6.105
R37371 S.n11906 S.t1756 6.105
R37372 S.n11918 S.n11917 6.105
R37373 S.n11921 S.n11920 6.105
R37374 S.n11903 S.t2664 6.105
R37375 S.n12911 S.t2760 6.105
R37376 S.n12923 S.n12922 6.105
R37377 S.n12926 S.n12925 6.105
R37378 S.n12908 S.t3745 6.105
R37379 S.n13904 S.t3614 6.105
R37380 S.n13916 S.n13915 6.105
R37381 S.n13919 S.n13918 6.105
R37382 S.n13901 S.t4571 6.105
R37383 S.n14874 S.t103 6.105
R37384 S.n14886 S.n14885 6.105
R37385 S.n14889 S.n14888 6.105
R37386 S.n14871 S.t1046 6.105
R37387 S.n15832 S.t2066 6.105
R37388 S.n15844 S.n15843 6.105
R37389 S.n15847 S.n15846 6.105
R37390 S.n15829 S.t3017 6.105
R37391 S.n16767 S.t700 6.105
R37392 S.n16779 S.n16778 6.105
R37393 S.n16782 S.n16781 6.105
R37394 S.n16764 S.t1658 6.105
R37395 S.n17690 S.t1741 6.105
R37396 S.n17702 S.n17701 6.105
R37397 S.n17705 S.n17704 6.105
R37398 S.n17687 S.t2650 6.105
R37399 S.n18590 S.t2742 6.105
R37400 S.n18602 S.n18601 6.105
R37401 S.n18605 S.n18604 6.105
R37402 S.n18587 S.t3734 6.105
R37403 S.n19480 S.t3818 6.105
R37404 S.n19492 S.n19491 6.105
R37405 S.n19495 S.n19494 6.105
R37406 S.n19477 S.t4219 6.105
R37407 S.n20226 S.t4322 6.105
R37408 S.n20243 S.n20242 6.105
R37409 S.n20240 S.n20239 6.105
R37410 S.n20223 S.t800 6.105
R37411 S.n19817 S.t2981 6.105
R37412 S.n19801 S.t3477 6.105
R37413 S.n18955 S.t1935 6.105
R37414 S.n18966 S.n18965 6.105
R37415 S.n18963 S.n18962 6.105
R37416 S.n18952 S.t2433 6.105
R37417 S.n18090 S.t889 6.105
R37418 S.n18101 S.n18100 6.105
R37419 S.n18098 S.n18097 6.105
R37420 S.n18087 S.t1388 6.105
R37421 S.n17201 S.t4605 6.105
R37422 S.n17212 S.n17211 6.105
R37423 S.n17209 S.n17208 6.105
R37424 S.n17198 S.t354 6.105
R37425 S.n16299 S.t3544 6.105
R37426 S.n16310 S.n16309 6.105
R37427 S.n16307 S.n16306 6.105
R37428 S.n16296 S.t4022 6.105
R37429 S.n15375 S.t403 6.105
R37430 S.n15386 S.n15385 6.105
R37431 S.n15383 S.n15382 6.105
R37432 S.n15372 S.t907 6.105
R37433 S.n14438 S.t3874 6.105
R37434 S.n14449 S.n14448 6.105
R37435 S.n14446 S.n14445 6.105
R37436 S.n14435 S.t4361 6.105
R37437 S.n13479 S.t2450 6.105
R37438 S.n13490 S.n13489 6.105
R37439 S.n13487 S.n13486 6.105
R37440 S.n13476 S.t2972 6.105
R37441 S.n12507 S.t1409 6.105
R37442 S.n12518 S.n12517 6.105
R37443 S.n12515 S.n12514 6.105
R37444 S.n12504 S.t1925 6.105
R37445 S.n11513 S.t373 6.105
R37446 S.n11524 S.n11523 6.105
R37447 S.n11521 S.n11520 6.105
R37448 S.n11510 S.t879 6.105
R37449 S.n10506 S.t3848 6.105
R37450 S.n10517 S.n10516 6.105
R37451 S.n10514 S.n10513 6.105
R37452 S.n10503 S.t4332 6.105
R37453 S.n9477 S.t2781 6.105
R37454 S.n9488 S.n9487 6.105
R37455 S.n9485 S.n9484 6.105
R37456 S.n9474 S.t3319 6.105
R37457 S.n8435 S.t1772 6.105
R37458 S.n8446 S.n8445 6.105
R37459 S.n8443 S.n8442 6.105
R37460 S.n8432 S.t2287 6.105
R37461 S.n7371 S.t933 6.105
R37462 S.n7382 S.n7381 6.105
R37463 S.n7379 S.n7378 6.105
R37464 S.n7368 S.t1192 6.105
R37465 S.n6294 S.t1140 6.105
R37466 S.n6305 S.n6304 6.105
R37467 S.n6302 S.n6301 6.105
R37468 S.n6291 S.t4343 6.105
R37469 S.n5194 S.t1093 6.105
R37470 S.n5205 S.n5204 6.105
R37471 S.n5202 S.n5201 6.105
R37472 S.n5191 S.t4289 6.105
R37473 S.n4082 S.t1606 6.105
R37474 S.n4093 S.n4092 6.105
R37475 S.n4090 S.n4089 6.105
R37476 S.n4079 S.t261 6.105
R37477 S.n2955 S.t4542 6.105
R37478 S.n2966 S.n2965 6.105
R37479 S.n2963 S.n2962 6.105
R37480 S.n2952 S.t3218 6.105
R37481 S.n2032 S.t2601 6.105
R37482 S.n2047 S.n2046 6.105
R37483 S.n2050 S.n2049 6.105
R37484 S.n2035 S.t3621 6.105
R37485 S.n753 S.t2879 6.105
R37486 S.n772 S.n771 6.105
R37487 S.n769 S.n768 6.105
R37488 S.n756 S.t1577 6.105
R37489 S.n1324 S.t2560 6.105
R37490 S.n1327 S.n1326 6.105
R37491 S.n1330 S.n1329 6.105
R37492 S.n1333 S.t3563 6.105
R37493 S.n1362 S.t1526 6.105
R37494 S.n1318 S.t2822 6.105
R37495 S.n20454 S.t2451 6.105
R37496 S.n20435 S.t2975 6.105
R37497 S.n20418 S.t3835 6.105
R37498 S.n20426 S.n20425 6.105
R37499 S.n20429 S.n20428 6.105
R37500 S.n20415 S.t275 6.105
R37501 S.n19835 S.t1417 6.105
R37502 S.n19844 S.n19843 6.105
R37503 S.n19841 S.n19840 6.105
R37504 S.n19832 S.t1929 6.105
R37505 S.n20314 S.t2767 6.105
R37506 S.n20332 S.n20331 6.105
R37507 S.n20335 S.n20334 6.105
R37508 S.n20311 S.t3754 6.105
R37509 S.n18983 S.t374 6.105
R37510 S.n18992 S.n18991 6.105
R37511 S.n18989 S.n18988 6.105
R37512 S.n18980 S.t885 6.105
R37513 S.n19442 S.t2279 6.105
R37514 S.n19460 S.n19459 6.105
R37515 S.n19463 S.n19462 6.105
R37516 S.n19439 S.t2668 6.105
R37517 S.n18118 S.t4046 6.105
R37518 S.n18126 S.n18125 6.105
R37519 S.n18123 S.n18122 6.105
R37520 S.n18115 S.t4335 6.105
R37521 S.n18555 S.t1183 6.105
R37522 S.n18570 S.n18569 6.105
R37523 S.n18573 S.n18572 6.105
R37524 S.n18552 S.t2187 6.105
R37525 S.n17229 S.t3047 6.105
R37526 S.n17237 S.n17236 6.105
R37527 S.n17234 S.n17233 6.105
R37528 S.n17226 S.t3538 6.105
R37529 S.n17655 S.t170 6.105
R37530 S.n17670 S.n17669 6.105
R37531 S.n17673 S.n17672 6.105
R37532 S.n17652 S.t1089 6.105
R37533 S.n16327 S.t4393 6.105
R37534 S.n16335 S.n16334 6.105
R37535 S.n16332 S.n16331 6.105
R37536 S.n16324 S.t397 6.105
R37537 S.n16732 S.t1564 6.105
R37538 S.n16747 S.n16746 6.105
R37539 S.n16750 S.n16749 6.105
R37540 S.n16729 S.t2481 6.105
R37541 S.n15403 S.t3366 6.105
R37542 S.n15411 S.n15410 6.105
R37543 S.n15408 S.n15407 6.105
R37544 S.n15400 S.t3870 6.105
R37545 S.n15797 S.t501 6.105
R37546 S.n15812 S.n15811 6.105
R37547 S.n15815 S.n15814 6.105
R37548 S.n15794 S.t1455 6.105
R37549 S.n14466 S.t2340 6.105
R37550 S.n14474 S.n14473 6.105
R37551 S.n14471 S.n14470 6.105
R37552 S.n14463 S.t2804 6.105
R37553 S.n14839 S.t3107 6.105
R37554 S.n14854 S.n14853 6.105
R37555 S.n14857 S.n14856 6.105
R37556 S.n14836 S.t4014 6.105
R37557 S.n13507 S.t903 6.105
R37558 S.n13515 S.n13514 6.105
R37559 S.n13512 S.n13511 6.105
R37560 S.n13504 S.t1404 6.105
R37561 S.n13869 S.t2294 6.105
R37562 S.n13884 S.n13883 6.105
R37563 S.n13887 S.n13886 6.105
R37564 S.n13866 S.t3243 6.105
R37565 S.n12535 S.t4358 6.105
R37566 S.n12543 S.n12542 6.105
R37567 S.n12540 S.n12539 6.105
R37568 S.n12532 S.t365 6.105
R37569 S.n12876 S.t1200 6.105
R37570 S.n12891 S.n12890 6.105
R37571 S.n12894 S.n12893 6.105
R37572 S.n12873 S.t2207 6.105
R37573 S.n11541 S.t3337 6.105
R37574 S.n11549 S.n11548 6.105
R37575 S.n11546 S.n11545 6.105
R37576 S.n11538 S.t3842 6.105
R37577 S.n11871 S.t186 6.105
R37578 S.n11886 S.n11885 6.105
R37579 S.n11889 S.n11888 6.105
R37580 S.n11868 S.t1104 6.105
R37581 S.n10534 S.t2310 6.105
R37582 S.n10542 S.n10541 6.105
R37583 S.n10539 S.n10538 6.105
R37584 S.n10531 S.t2775 6.105
R37585 S.n10843 S.t3669 6.105
R37586 S.n10858 S.n10857 6.105
R37587 S.n10861 S.n10860 6.105
R37588 S.n10840 S.t46 6.105
R37589 S.n9505 S.t1219 6.105
R37590 S.n9513 S.n9512 6.105
R37591 S.n9510 S.n9509 6.105
R37592 S.n9502 S.t1768 6.105
R37593 S.n9803 S.t3151 6.105
R37594 S.n9818 S.n9817 6.105
R37595 S.n9821 S.n9820 6.105
R37596 S.n9800 S.t3577 6.105
R37597 S.n8463 S.t431 6.105
R37598 S.n8471 S.n8470 6.105
R37599 S.n8468 S.n8467 6.105
R37600 S.n8460 S.t727 6.105
R37601 S.n8740 S.t2099 6.105
R37602 S.n8755 S.n8754 6.105
R37603 S.n8758 S.n8757 6.105
R37604 S.n8737 S.t3053 6.105
R37605 S.n7399 S.t4143 6.105
R37606 S.n7407 S.n7406 6.105
R37607 S.n7404 S.n7403 6.105
R37608 S.n7396 S.t2844 6.105
R37609 S.n7665 S.t2150 6.105
R37610 S.n7680 S.n7679 6.105
R37611 S.n7683 S.n7682 6.105
R37612 S.n7662 S.t3119 6.105
R37613 S.n6322 S.t4096 6.105
R37614 S.n6330 S.n6329 6.105
R37615 S.n6327 S.n6326 6.105
R37616 S.n6319 S.t2785 6.105
R37617 S.n6567 S.t2095 6.105
R37618 S.n6582 S.n6581 6.105
R37619 S.n6585 S.n6584 6.105
R37620 S.n6564 S.t3068 6.105
R37621 S.n5222 S.t4056 6.105
R37622 S.n5230 S.n5229 6.105
R37623 S.n5227 S.n5226 6.105
R37624 S.n5219 S.t2733 6.105
R37625 S.n5457 S.t2524 6.105
R37626 S.n5472 S.n5471 6.105
R37627 S.n5475 S.n5474 6.105
R37628 S.n5454 S.t3514 6.105
R37629 S.n4110 S.t4567 6.105
R37630 S.n4118 S.n4117 6.105
R37631 S.n4115 S.n4114 6.105
R37632 S.n4107 S.t3241 6.105
R37633 S.n4322 S.t2486 6.105
R37634 S.n4337 S.n4336 6.105
R37635 S.n4340 S.n4339 6.105
R37636 S.n4319 S.t3471 6.105
R37637 S.n2983 S.t2983 6.105
R37638 S.n2991 S.n2990 6.105
R37639 S.n2988 S.n2987 6.105
R37640 S.n2980 S.t1668 6.105
R37641 S.n3185 S.t2654 6.105
R37642 S.n3200 S.n3199 6.105
R37643 S.n3203 S.n3202 6.105
R37644 S.n3182 S.t3660 6.105
R37645 S.n1820 S.t2929 6.105
R37646 S.n1828 S.n1827 6.105
R37647 S.n1825 S.n1824 6.105
R37648 S.n1817 S.t1620 6.105
R37649 S.n1999 S.t1047 6.105
R37650 S.n2014 S.n2013 6.105
R37651 S.n2017 S.n2016 6.105
R37652 S.n2002 S.t2062 6.105
R37653 S.n777 S.t1312 6.105
R37654 S.n791 S.n790 6.105
R37655 S.n788 S.n787 6.105
R37656 S.n780 S.t4531 6.105
R37657 S.n1841 S.t1364 6.105
R37658 S.n1850 S.n1849 6.105
R37659 S.n1847 S.n1846 6.105
R37660 S.n1838 S.t4577 6.105
R37661 S.n3160 S.t1092 6.105
R37662 S.n3168 S.n3167 6.105
R37663 S.n3171 S.n3170 6.105
R37664 S.n3163 S.t2112 6.105
R37665 S.n2997 S.t1420 6.105
R37666 S.n3011 S.n3010 6.105
R37667 S.n3008 S.n3007 6.105
R37668 S.n3000 S.t34 6.105
R37669 S.n4297 S.t1139 6.105
R37670 S.n4305 S.n4304 6.105
R37671 S.n4308 S.n4307 6.105
R37672 S.n4300 S.t2159 6.105
R37673 S.n4124 S.t3009 6.105
R37674 S.n4137 S.n4136 6.105
R37675 S.n4134 S.n4133 6.105
R37676 S.n4127 S.t1690 6.105
R37677 S.n5431 S.t976 6.105
R37678 S.n5440 S.n5439 6.105
R37679 S.n5443 S.n5442 6.105
R37680 S.n5434 S.t1966 6.105
R37681 S.n5236 S.t2514 6.105
R37682 S.n5250 S.n5249 6.105
R37683 S.n5247 S.n5246 6.105
R37684 S.n5239 S.t1173 6.105
R37685 S.n6542 S.t529 6.105
R37686 S.n6550 S.n6549 6.105
R37687 S.n6553 S.n6552 6.105
R37688 S.n6545 S.t1517 6.105
R37689 S.n6336 S.t2553 6.105
R37690 S.n6350 S.n6349 6.105
R37691 S.n6347 S.n6346 6.105
R37692 S.n6339 S.t1225 6.105
R37693 S.n7640 S.t584 6.105
R37694 S.n7648 S.n7647 6.105
R37695 S.n7651 S.n7650 6.105
R37696 S.n7643 S.t1568 6.105
R37697 S.n7413 S.t2595 6.105
R37698 S.n7427 S.n7426 6.105
R37699 S.n7424 S.n7423 6.105
R37700 S.n7416 S.t1275 6.105
R37701 S.n8715 S.t640 6.105
R37702 S.n8723 S.n8722 6.105
R37703 S.n8726 S.n8725 6.105
R37704 S.n8718 S.t1612 6.105
R37705 S.n8477 S.t2644 6.105
R37706 S.n8491 S.n8490 6.105
R37707 S.n8488 S.n8487 6.105
R37708 S.n8480 S.t1329 6.105
R37709 S.n9778 S.t1596 6.105
R37710 S.n9786 S.n9785 6.105
R37711 S.n9789 S.n9788 6.105
R37712 S.n9781 S.t2026 6.105
R37713 S.n9519 S.t4431 6.105
R37714 S.n9533 S.n9532 6.105
R37715 S.n9530 S.n9529 6.105
R37716 S.n9522 S.t199 6.105
R37717 S.n10818 S.t2123 6.105
R37718 S.n10826 S.n10825 6.105
R37719 S.n10829 S.n10828 6.105
R37720 S.n10821 S.t3074 6.105
R37721 S.n10548 S.t748 6.105
R37722 S.n10562 S.n10561 6.105
R37723 S.n10559 S.n10558 6.105
R37724 S.n10551 S.t1214 6.105
R37725 S.n11846 S.t3170 6.105
R37726 S.n11854 S.n11853 6.105
R37727 S.n11857 S.n11856 6.105
R37728 S.n11849 S.t4066 6.105
R37729 S.n11555 S.t1790 6.105
R37730 S.n11569 S.n11568 6.105
R37731 S.n11566 S.n11565 6.105
R37732 S.n11558 S.t2306 6.105
R37733 S.n12851 S.t4154 6.105
R37734 S.n12859 S.n12858 6.105
R37735 S.n12862 S.n12861 6.105
R37736 S.n12854 S.t646 6.105
R37737 S.n12549 S.t2800 6.105
R37738 S.n12563 S.n12562 6.105
R37739 S.n12560 S.n12559 6.105
R37740 S.n12552 S.t3332 6.105
R37741 S.n13844 S.t732 6.105
R37742 S.n13852 S.n13851 6.105
R37743 S.n13855 S.n13854 6.105
R37744 S.n13847 S.t1691 6.105
R37745 S.n13521 S.t3866 6.105
R37746 S.n13535 S.n13534 6.105
R37747 S.n13532 S.n13531 6.105
R37748 S.n13524 S.t4352 6.105
R37749 S.n14814 S.t1773 6.105
R37750 S.n14822 S.n14821 6.105
R37751 S.n14825 S.n14824 6.105
R37752 S.n14817 S.t2683 6.105
R37753 S.n14480 S.t785 6.105
R37754 S.n14494 S.n14493 6.105
R37755 S.n14491 S.n14490 6.105
R37756 S.n14483 S.t1244 6.105
R37757 S.n15772 S.t3461 6.105
R37758 S.n15780 S.n15779 6.105
R37759 S.n15783 S.n15782 6.105
R37760 S.n15775 S.t4404 6.105
R37761 S.n15417 S.t1821 6.105
R37762 S.n15431 S.n15430 6.105
R37763 S.n15428 S.n15427 6.105
R37764 S.n15420 S.t2331 6.105
R37765 S.n16707 S.t4514 6.105
R37766 S.n16715 S.n16714 6.105
R37767 S.n16718 S.n16717 6.105
R37768 S.n16710 S.t931 6.105
R37769 S.n16341 S.t2837 6.105
R37770 S.n16355 S.n16354 6.105
R37771 S.n16352 S.n16351 6.105
R37772 S.n16344 S.t3361 6.105
R37773 S.n17630 S.t1011 6.105
R37774 S.n17638 S.n17637 6.105
R37775 S.n17641 S.n17640 6.105
R37776 S.n17633 S.t1988 6.105
R37777 S.n17243 S.t3893 6.105
R37778 S.n17257 S.n17256 6.105
R37779 S.n17254 S.n17253 6.105
R37780 S.n17246 S.t4385 6.105
R37781 S.n18530 S.t4138 6.105
R37782 S.n18538 S.n18537 6.105
R37783 S.n18541 S.n18540 6.105
R37784 S.n18533 S.t628 6.105
R37785 S.n18132 S.t2504 6.105
R37786 S.n18146 S.n18145 6.105
R37787 S.n18143 S.n18142 6.105
R37788 S.n18135 S.t3040 6.105
R37789 S.n19417 S.t716 6.105
R37790 S.n19425 S.n19424 6.105
R37791 S.n19428 S.n19427 6.105
R37792 S.n19420 S.t1112 6.105
R37793 S.n18998 S.t3568 6.105
R37794 S.n19012 S.n19011 6.105
R37795 S.n19009 S.n19008 6.105
R37796 S.n19001 S.t3846 6.105
R37797 S.n20289 S.t1203 6.105
R37798 S.n20297 S.n20296 6.105
R37799 S.n20300 S.n20299 6.105
R37800 S.n20292 S.t2212 6.105
R37801 S.n19852 S.t4362 6.105
R37802 S.n19866 S.n19865 6.105
R37803 S.n19863 S.n19862 6.105
R37804 S.n19855 S.t372 6.105
R37805 S.n20360 S.t2301 6.105
R37806 S.n20371 S.n20370 6.105
R37807 S.n20368 S.n20367 6.105
R37808 S.n20363 S.t3250 6.105
R37809 S.n20463 S.t905 6.105
R37810 S.n20477 S.n20476 6.105
R37811 S.n20474 S.n20473 6.105
R37812 S.n20466 S.t1407 6.105
R37813 S.n21236 S.t3327 6.105
R37814 S.n21244 S.n21243 6.105
R37815 S.n21247 S.n21246 6.105
R37816 S.n21239 S.t4239 6.105
R37817 S.n21299 S.t1952 6.105
R37818 S.n21281 S.t2445 6.105
R37819 S.n1379 S.t4471 6.105
R37820 S.n1366 S.t1257 6.105
R37821 S.n852 S.t1013 6.105
R37822 S.n869 S.n868 6.105
R37823 S.n866 S.n865 6.105
R37824 S.n855 S.t2013 6.105
R37825 S.n2093 S.t984 6.105
R37826 S.n2109 S.n2108 6.105
R37827 S.n2112 S.n2111 6.105
R37828 S.n2096 S.t1976 6.105
R37829 S.n737 S.t1487 6.105
R37830 S.n748 S.n747 6.105
R37831 S.n745 S.n744 6.105
R37832 S.n740 S.t123 6.105
R37833 S.n720 S.t3044 6.105
R37834 S.n731 S.n730 6.105
R37835 S.n728 S.n727 6.105
R37836 S.n723 S.t1716 6.105
R37837 S.n1288 S.t248 6.105
R37838 S.n1281 S.t1594 6.105
R37839 S.n368 S.t1069 6.105
R37840 S.n379 S.n378 6.105
R37841 S.n376 S.n375 6.105
R37842 S.n371 S.t2085 6.105
R37843 S.n2188 S.t1117 6.105
R37844 S.n2198 S.n2197 6.105
R37845 S.n2201 S.n2200 6.105
R37846 S.n2185 S.t2135 6.105
R37847 S.n16235 S.t505 6.105
R37848 S.n16219 S.t991 6.105
R37849 S.n16648 S.t2392 6.105
R37850 S.n16665 S.n16664 6.105
R37851 S.n16662 S.n16661 6.105
R37852 S.n16645 S.t3343 6.105
R37853 S.n15301 S.t3959 6.105
R37854 S.n15312 S.n15311 6.105
R37855 S.n15309 S.n15308 6.105
R37856 S.n15298 S.t4485 6.105
R37857 S.n15958 S.t1326 6.105
R37858 S.n15970 S.n15969 6.105
R37859 S.n15973 S.n15972 6.105
R37860 S.n15955 S.t2317 6.105
R37861 S.n14366 S.t2938 6.105
R37862 S.n14377 S.n14376 6.105
R37863 S.n14374 S.n14373 6.105
R37864 S.n14363 S.t3439 6.105
R37865 S.n14996 S.t3924 6.105
R37866 S.n15008 S.n15007 6.105
R37867 S.n15011 S.n15010 6.105
R37868 S.n14993 S.t369 6.105
R37869 S.n13407 S.t1758 6.105
R37870 S.n13418 S.n13417 6.105
R37871 S.n13415 S.n13414 6.105
R37872 S.n13404 S.t2032 6.105
R37873 S.n14026 S.t2887 6.105
R37874 S.n14038 S.n14037 6.105
R37875 S.n14041 S.n14040 6.105
R37876 S.n14023 S.t3845 6.105
R37877 S.n12435 S.t715 6.105
R37878 S.n12446 S.n12445 6.105
R37879 S.n12443 S.n12442 6.105
R37880 S.n12432 S.t1177 6.105
R37881 S.n13033 S.t1857 6.105
R37882 S.n13045 S.n13044 6.105
R37883 S.n13048 S.n13047 6.105
R37884 S.n13030 S.t2780 6.105
R37885 S.n11441 S.t2087 6.105
R37886 S.n11452 S.n11451 6.105
R37887 S.n11449 S.n11448 6.105
R37888 S.n11438 S.t2552 6.105
R37889 S.n12028 S.t3236 6.105
R37890 S.n12040 S.n12039 6.105
R37891 S.n12043 S.n12042 6.105
R37892 S.n12025 S.t4132 6.105
R37893 S.n10434 S.t1008 6.105
R37894 S.n10445 S.n10444 6.105
R37895 S.n10442 S.n10441 6.105
R37896 S.n10431 S.t1557 6.105
R37897 S.n11000 S.t2198 6.105
R37898 S.n11012 S.n11011 6.105
R37899 S.n11015 S.n11014 6.105
R37900 S.n10997 S.t3147 6.105
R37901 S.n9405 S.t4513 6.105
R37902 S.n9416 S.n9415 6.105
R37903 S.n9413 S.n9412 6.105
R37904 S.n9402 S.t493 6.105
R37905 S.n9960 S.t1666 6.105
R37906 S.n9972 S.n9971 6.105
R37907 S.n9975 S.n9974 6.105
R37908 S.n9957 S.t2100 6.105
R37909 S.n8363 S.t3460 6.105
R37910 S.n8374 S.n8373 6.105
R37911 S.n8371 S.n8370 6.105
R37912 S.n8360 S.t3950 6.105
R37913 S.n8897 S.t834 6.105
R37914 S.n8909 S.n8908 6.105
R37915 S.n8912 S.n8911 6.105
R37916 S.n8894 S.t1791 6.105
R37917 S.n7299 S.t2417 6.105
R37918 S.n7310 S.n7309 6.105
R37919 S.n7307 S.n7306 6.105
R37920 S.n7296 S.t2926 6.105
R37921 S.n7822 S.t4273 6.105
R37922 S.n7834 S.n7833 6.105
R37923 S.n7837 S.n7836 6.105
R37924 S.n7819 S.t752 6.105
R37925 S.n6222 S.t1369 6.105
R37926 S.n6233 S.n6232 6.105
R37927 S.n6230 S.n6229 6.105
R37928 S.n6219 S.t1892 6.105
R37929 S.n6724 S.t3272 6.105
R37930 S.n6736 S.n6735 6.105
R37931 S.n6739 S.n6738 6.105
R37932 S.n6721 S.t4173 6.105
R37933 S.n5122 S.t337 6.105
R37934 S.n5133 S.n5132 6.105
R37935 S.n5130 S.n5129 6.105
R37936 S.n5119 S.t848 6.105
R37937 S.n5614 S.t289 6.105
R37938 S.n5626 S.n5625 6.105
R37939 S.n5629 S.n5628 6.105
R37940 S.n5611 S.t1205 6.105
R37941 S.n4010 S.t1884 6.105
R37942 S.n4021 S.n4020 6.105
R37943 S.n4018 S.n4017 6.105
R37944 S.n4007 S.t2389 6.105
R37945 S.n4479 S.t3772 6.105
R37946 S.n4491 S.n4490 6.105
R37947 S.n4494 S.n4493 6.105
R37948 S.n4476 S.t195 6.105
R37949 S.n2883 S.t1589 6.105
R37950 S.n2894 S.n2893 6.105
R37951 S.n2891 S.n2890 6.105
R37952 S.n2880 S.t1863 6.105
R37953 S.n3341 S.t2687 6.105
R37954 S.n3352 S.n3351 6.105
R37955 S.n3355 S.n3354 6.105
R37956 S.n3338 S.t3678 6.105
R37957 S.n1713 S.t1687 6.105
R37958 S.n1725 S.n1724 6.105
R37959 S.n1722 S.n1721 6.105
R37960 S.n1710 S.t343 6.105
R37961 S.n1414 S.t3226 6.105
R37962 S.n1415 S.t4551 6.105
R37963 S.n59 S.t4035 6.105
R37964 S.n62 S.n61 6.105
R37965 S.n65 S.n64 6.105
R37966 S.n68 S.t521 6.105
R37967 S.n17154 S.t4518 6.105
R37968 S.n17137 S.t499 6.105
R37969 S.n17570 S.t1880 6.105
R37970 S.n17588 S.n17587 6.105
R37971 S.n17585 S.n17584 6.105
R37972 S.n17573 S.t2807 6.105
R37973 S.n16244 S.t3465 6.105
R37974 S.n16255 S.n16254 6.105
R37975 S.n16252 S.n16251 6.105
R37976 S.n16247 S.t3953 6.105
R37977 S.n16856 S.t839 6.105
R37978 S.n16873 S.n16872 6.105
R37979 S.n16876 S.n16875 6.105
R37980 S.n16859 S.t1796 6.105
R37981 S.n15320 S.t2420 6.105
R37982 S.n15331 S.n15330 6.105
R37983 S.n15328 S.n15327 6.105
R37984 S.n15323 S.t2931 6.105
R37985 S.n15921 S.t4277 6.105
R37986 S.n15938 S.n15937 6.105
R37987 S.n15941 S.n15940 6.105
R37988 S.n15924 S.t757 6.105
R37989 S.n14383 S.t1630 6.105
R37990 S.n14394 S.n14393 6.105
R37991 S.n14391 S.n14390 6.105
R37992 S.n14386 S.t1893 6.105
R37993 S.n14959 S.t2384 6.105
R37994 S.n14976 S.n14975 6.105
R37995 S.n14979 S.n14978 6.105
R37996 S.n14962 S.t3333 6.105
R37997 S.n13424 S.t189 6.105
R37998 S.n13435 S.n13434 6.105
R37999 S.n13432 S.n13431 6.105
R38000 S.n13427 S.t708 6.105
R38001 S.n13989 S.t1318 6.105
R38002 S.n14006 S.n14005 6.105
R38003 S.n14009 S.n14008 6.105
R38004 S.n13992 S.t2308 6.105
R38005 S.n12452 S.t1582 6.105
R38006 S.n12463 S.n12462 6.105
R38007 S.n12460 S.n12459 6.105
R38008 S.n12455 S.t2078 6.105
R38009 S.n12996 S.t2673 6.105
R38010 S.n13013 S.n13012 6.105
R38011 S.n13016 S.n13015 6.105
R38012 S.n12999 S.t3666 6.105
R38013 S.n11458 S.t518 6.105
R38014 S.n11469 S.n11468 6.105
R38015 S.n11466 S.n11465 6.105
R38016 S.n11461 S.t1003 6.105
R38017 S.n11991 S.t1683 6.105
R38018 S.n12008 S.n12007 6.105
R38019 S.n12011 S.n12010 6.105
R38020 S.n11994 S.t2587 6.105
R38021 S.n10451 S.t3973 6.105
R38022 S.n10462 S.n10461 6.105
R38023 S.n10459 S.n10458 6.105
R38024 S.n10454 S.t4502 6.105
R38025 S.n10963 S.t636 6.105
R38026 S.n10980 S.n10979 6.105
R38027 S.n10983 S.n10982 6.105
R38028 S.n10966 S.t1592 6.105
R38029 S.n9422 S.t2956 6.105
R38030 S.n9433 S.n9432 6.105
R38031 S.n9430 S.n9429 6.105
R38032 S.n9425 S.t3454 6.105
R38033 S.n9923 S.t313 6.105
R38034 S.n9940 S.n9939 6.105
R38035 S.n9943 S.n9942 6.105
R38036 S.n9926 S.t775 6.105
R38037 S.n8380 S.t1914 6.105
R38038 S.n8391 S.n8390 6.105
R38039 S.n8388 S.n8387 6.105
R38040 S.n8383 S.t2412 6.105
R38041 S.n8860 S.t3796 6.105
R38042 S.n8877 S.n8876 6.105
R38043 S.n8880 S.n8879 6.105
R38044 S.n8863 S.t225 6.105
R38045 S.n7316 S.t871 6.105
R38046 S.n7327 S.n7326 6.105
R38047 S.n7324 S.n7323 6.105
R38048 S.n7319 S.t1359 6.105
R38049 S.n7785 S.t2718 6.105
R38050 S.n7802 S.n7801 6.105
R38051 S.n7805 S.n7804 6.105
R38052 S.n7788 S.t3709 6.105
R38053 S.n6239 S.t4317 6.105
R38054 S.n6250 S.n6249 6.105
R38055 S.n6247 S.n6246 6.105
R38056 S.n6242 S.t333 6.105
R38057 S.n6687 S.t1719 6.105
R38058 S.n6704 S.n6703 6.105
R38059 S.n6707 S.n6706 6.105
R38060 S.n6690 S.t2621 6.105
R38061 S.n5139 S.t3303 6.105
R38062 S.n5150 S.n5149 6.105
R38063 S.n5147 S.n5146 6.105
R38064 S.n5142 S.t3809 6.105
R38065 S.n5577 S.t3262 6.105
R38066 S.n5594 S.n5593 6.105
R38067 S.n5597 S.n5596 6.105
R38068 S.n5580 S.t4161 6.105
R38069 S.n4027 S.t551 6.105
R38070 S.n4038 S.n4037 6.105
R38071 S.n4035 S.n4034 6.105
R38072 S.n4030 S.t837 6.105
R38073 S.n4442 S.t2228 6.105
R38074 S.n4459 S.n4458 6.105
R38075 S.n4462 S.n4461 6.105
R38076 S.n4445 S.t3176 6.105
R38077 S.n2900 S.t145 6.105
R38078 S.n2911 S.n2910 6.105
R38079 S.n2908 S.n2907 6.105
R38080 S.n2903 S.t3350 6.105
R38081 S.n3304 S.t4119 6.105
R38082 S.n3321 S.n3320 6.105
R38083 S.n3324 S.n3323 6.105
R38084 S.n3307 S.t623 6.105
R38085 S.n1731 S.t76 6.105
R38086 S.n1742 S.n1741 6.105
R38087 S.n1739 S.n1738 6.105
R38088 S.n1734 S.t3311 6.105
R38089 S.n2151 S.t4074 6.105
R38090 S.n2168 S.n2167 6.105
R38091 S.n2171 S.n2170 6.105
R38092 S.n2154 S.t572 6.105
R38093 S.n702 S.t4600 6.105
R38094 S.n713 S.n712 6.105
R38095 S.n710 S.n709 6.105
R38096 S.n705 S.t3268 6.105
R38097 S.n685 S.t1646 6.105
R38098 S.n696 S.n695 6.105
R38099 S.n693 S.n692 6.105
R38100 S.n688 S.t299 6.105
R38101 S.n1276 S.t3364 6.105
R38102 S.n1268 S.t159 6.105
R38103 S.n336 S.t3751 6.105
R38104 S.n347 S.n346 6.105
R38105 S.n344 S.n343 6.105
R38106 S.n339 S.t171 6.105
R38107 S.n2247 S.t271 6.105
R38108 S.n2257 S.n2256 6.105
R38109 S.n2260 S.n2259 6.105
R38110 S.n2244 S.t1184 6.105
R38111 S.n14338 S.t1547 6.105
R38112 S.n14322 S.t2042 6.105
R38113 S.n14755 S.t2506 6.105
R38114 S.n14772 S.n14771 6.105
R38115 S.n14769 S.n14768 6.105
R38116 S.n14752 S.t3476 6.105
R38117 S.n13369 S.t74 6.105
R38118 S.n13380 S.n13379 6.105
R38119 S.n13377 S.n13376 6.105
R38120 S.n13366 S.t635 6.105
R38121 S.n14091 S.t1494 6.105
R38122 S.n14103 S.n14102 6.105
R38123 S.n14106 S.n14105 6.105
R38124 S.n14088 S.t2429 6.105
R38125 S.n12399 S.t3591 6.105
R38126 S.n12410 S.n12409 6.105
R38127 S.n12407 S.n12406 6.105
R38128 S.n12396 S.t4059 6.105
R38129 S.n13094 S.t444 6.105
R38130 S.n13106 S.n13105 6.105
R38131 S.n13109 S.n13108 6.105
R38132 S.n13091 S.t1387 6.105
R38133 S.n11405 S.t2739 6.105
R38134 S.n11416 S.n11415 6.105
R38135 S.n11413 S.n11412 6.105
R38136 S.n11402 S.t3065 6.105
R38137 S.n12089 S.t3905 6.105
R38138 S.n12101 S.n12100 6.105
R38139 S.n12104 S.n12103 6.105
R38140 S.n12086 S.t353 6.105
R38141 S.n10398 S.t1740 6.105
R38142 S.n10409 S.n10408 6.105
R38143 S.n10406 S.n10405 6.105
R38144 S.n10395 S.t2250 6.105
R38145 S.n11061 S.t2863 6.105
R38146 S.n11073 S.n11072 6.105
R38147 S.n11076 S.n11075 6.105
R38148 S.n11058 S.t3828 6.105
R38149 S.n9369 S.t3113 6.105
R38150 S.n9380 S.n9379 6.105
R38151 S.n9377 S.n9376 6.105
R38152 S.n9366 S.t3615 6.105
R38153 S.n10021 S.t236 6.105
R38154 S.n10033 S.n10032 6.105
R38155 S.n10036 S.n10035 6.105
R38156 S.n10018 S.t692 6.105
R38157 S.n8327 S.t2065 6.105
R38158 S.n8338 S.n8337 6.105
R38159 S.n8335 S.n8334 6.105
R38160 S.n8324 S.t2537 6.105
R38161 S.n8958 S.t3720 6.105
R38162 S.n8970 S.n8969 6.105
R38163 S.n8973 S.n8972 6.105
R38164 S.n8955 S.t124 6.105
R38165 S.n7263 S.t992 6.105
R38166 S.n7274 S.n7273 6.105
R38167 S.n7271 S.n7270 6.105
R38168 S.n7260 S.t1533 6.105
R38169 S.n7883 S.t2636 6.105
R38170 S.n7895 S.n7894 6.105
R38171 S.n7898 S.n7897 6.105
R38172 S.n7880 S.t3632 6.105
R38173 S.n6186 S.t4484 6.105
R38174 S.n6197 S.n6196 6.105
R38175 S.n6194 S.n6193 6.105
R38176 S.n6183 S.t476 6.105
R38177 S.n6785 S.t1864 6.105
R38178 S.n6797 S.n6796 6.105
R38179 S.n6800 S.n6799 6.105
R38180 S.n6782 S.t2783 6.105
R38181 S.n5086 S.t3443 6.105
R38182 S.n5097 S.n5096 6.105
R38183 S.n5094 S.n5093 6.105
R38184 S.n5083 S.t3940 6.105
R38185 S.n5675 S.t3392 6.105
R38186 S.n5687 S.n5686 6.105
R38187 S.n5690 S.n5689 6.105
R38188 S.n5672 S.t4326 6.105
R38189 S.n3974 S.t469 6.105
R38190 S.n3985 S.n3984 6.105
R38191 S.n3982 S.n3981 6.105
R38192 S.n3971 S.t962 6.105
R38193 S.n4540 S.t2366 6.105
R38194 S.n4552 S.n4551 6.105
R38195 S.n4555 S.n4554 6.105
R38196 S.n4537 S.t3314 6.105
R38197 S.n2847 S.t4452 6.105
R38198 S.n2858 S.n2857 6.105
R38199 S.n2855 S.n2854 6.105
R38200 S.n2844 S.t449 6.105
R38201 S.n3401 S.t1288 6.105
R38202 S.n3412 S.n3411 6.105
R38203 S.n3415 S.n3414 6.105
R38204 S.n3398 S.t2284 6.105
R38205 S.n1676 S.t3408 6.105
R38206 S.n1688 S.n1687 6.105
R38207 S.n1685 S.n1684 6.105
R38208 S.n1673 S.t3907 6.105
R38209 S.n1410 S.t1817 6.105
R38210 S.n1411 S.t3149 6.105
R38211 S.n91 S.t2624 6.105
R38212 S.n94 S.n93 6.105
R38213 S.n97 S.n96 6.105
R38214 S.n100 S.t3637 6.105
R38215 S.n15292 S.t996 6.105
R38216 S.n15275 S.t1535 6.105
R38217 S.n15712 S.t2892 6.105
R38218 S.n15730 S.n15729 6.105
R38219 S.n15727 S.n15726 6.105
R38220 S.n15715 S.t3854 6.105
R38221 S.n14347 S.t4494 6.105
R38222 S.n14358 S.n14357 6.105
R38223 S.n14355 S.n14354 6.105
R38224 S.n14350 S.t479 6.105
R38225 S.n15024 S.t955 6.105
R38226 S.n15041 S.n15040 6.105
R38227 S.n15044 S.n15043 6.105
R38228 S.n15027 S.t1928 6.105
R38229 S.n13388 S.t3088 6.105
R38230 S.n13399 S.n13398 6.105
R38231 S.n13396 S.n13395 6.105
R38232 S.n13391 S.t3586 6.105
R38233 S.n14054 S.t4442 6.105
R38234 S.n14071 S.n14070 6.105
R38235 S.n14074 S.n14073 6.105
R38236 S.n14057 S.t882 6.105
R38237 S.n12416 S.t2278 6.105
R38238 S.n12427 S.n12426 6.105
R38239 S.n12424 S.n12423 6.105
R38240 S.n12419 S.t2517 6.105
R38241 S.n13057 S.t3400 6.105
R38242 S.n13074 S.n13073 6.105
R38243 S.n13077 S.n13076 6.105
R38244 S.n13060 S.t4334 6.105
R38245 S.n11422 S.t1182 6.105
R38246 S.n11433 S.n11432 6.105
R38247 S.n11430 S.n11429 6.105
R38248 S.n11425 S.t1732 6.105
R38249 S.n12052 S.t2373 6.105
R38250 S.n12069 S.n12068 6.105
R38251 S.n12072 S.n12071 6.105
R38252 S.n12055 S.t3321 6.105
R38253 S.n10415 S.t2556 6.105
R38254 S.n10426 S.n10425 6.105
R38255 S.n10423 S.n10422 6.105
R38256 S.n10418 S.t3109 6.105
R38257 S.n11024 S.t3741 6.105
R38258 S.n11041 S.n11040 6.105
R38259 S.n11044 S.n11043 6.105
R38260 S.n11027 S.t155 6.105
R38261 S.n9386 S.t1562 6.105
R38262 S.n9397 S.n9396 6.105
R38263 S.n9394 S.n9393 6.105
R38264 S.n9389 S.t2059 6.105
R38265 S.n9984 S.t3215 6.105
R38266 S.n10001 S.n10000 6.105
R38267 S.n10004 S.n10003 6.105
R38268 S.n9987 S.t3649 6.105
R38269 S.n8344 S.t500 6.105
R38270 S.n8355 S.n8354 6.105
R38271 S.n8352 S.n8351 6.105
R38272 S.n8347 S.t988 6.105
R38273 S.n8921 S.t2178 6.105
R38274 S.n8938 S.n8937 6.105
R38275 S.n8941 S.n8940 6.105
R38276 S.n8924 S.t3128 6.105
R38277 S.n7280 S.t3955 6.105
R38278 S.n7291 S.n7290 6.105
R38279 S.n7288 S.n7287 6.105
R38280 S.n7283 S.t4480 6.105
R38281 S.n7846 S.t1323 6.105
R38282 S.n7863 S.n7862 6.105
R38283 S.n7866 S.n7865 6.105
R38284 S.n7849 S.t2311 6.105
R38285 S.n6203 S.t2935 6.105
R38286 S.n6214 S.n6213 6.105
R38287 S.n6211 S.n6210 6.105
R38288 S.n6206 S.t3435 6.105
R38289 S.n6748 S.t302 6.105
R38290 S.n6765 S.n6764 6.105
R38291 S.n6768 S.n6767 6.105
R38292 S.n6751 S.t1223 6.105
R38293 S.n5103 S.t1897 6.105
R38294 S.n5114 S.n5113 6.105
R38295 S.n5111 S.n5110 6.105
R38296 S.n5106 S.t2401 6.105
R38297 S.n5638 S.t1849 6.105
R38298 S.n5655 S.n5654 6.105
R38299 S.n5658 S.n5657 6.105
R38300 S.n5641 S.t2770 6.105
R38301 S.n3991 S.t3429 6.105
R38302 S.n4002 S.n4001 6.105
R38303 S.n3999 S.n3998 6.105
R38304 S.n3994 S.t3929 6.105
R38305 S.n4503 S.t812 6.105
R38306 S.n4520 S.n4519 6.105
R38307 S.n4523 S.n4522 6.105
R38308 S.n4506 S.t1764 6.105
R38309 S.n2864 S.t2896 6.105
R38310 S.n2875 S.n2874 6.105
R38311 S.n2872 S.n2871 6.105
R38312 S.n2867 S.t3405 6.105
R38313 S.n3364 S.t4238 6.105
R38314 S.n3381 S.n3380 6.105
R38315 S.n3384 S.n3383 6.105
R38316 S.n3367 S.t721 6.105
R38317 S.n1694 S.t2094 6.105
R38318 S.n1705 S.n1704 6.105
R38319 S.n1702 S.n1701 6.105
R38320 S.n1697 S.t2374 6.105
R38321 S.n2210 S.t3245 6.105
R38322 S.n2227 S.n2226 6.105
R38323 S.n2230 S.n2229 6.105
R38324 S.n2213 S.t4139 6.105
R38325 S.n667 S.t3197 6.105
R38326 S.n678 S.n677 6.105
R38327 S.n675 S.n674 6.105
R38328 S.n670 S.t1859 6.105
R38329 S.n650 S.t2564 6.105
R38330 S.n661 S.n660 6.105
R38331 S.n658 S.n657 6.105
R38332 S.n653 S.t2866 6.105
R38333 S.n1263 S.t425 6.105
R38334 S.n1255 S.t4426 6.105
R38335 S.n304 S.t2352 6.105
R38336 S.n315 S.n314 6.105
R38337 S.n312 S.n311 6.105
R38338 S.n307 S.t3293 6.105
R38339 S.n2306 S.t3380 6.105
R38340 S.n2316 S.n2315 6.105
R38341 S.n2319 S.n2318 6.105
R38342 S.n2303 S.t4301 6.105
R38343 S.n12371 S.t2199 6.105
R38344 S.n12355 S.t2657 6.105
R38345 S.n12792 S.t3549 6.105
R38346 S.n12809 S.n12808 6.105
R38347 S.n12806 S.n12805 6.105
R38348 S.n12789 S.t4505 6.105
R38349 S.n11367 S.t1098 6.105
R38350 S.n11378 S.n11377 6.105
R38351 S.n11375 S.n11374 6.105
R38352 S.n11364 S.t1664 6.105
R38353 S.n12154 S.t2490 6.105
R38354 S.n12166 S.n12165 6.105
R38355 S.n12169 S.n12168 6.105
R38356 S.n12151 S.t3458 6.105
R38357 S.n10362 S.t32 6.105
R38358 S.n10373 S.n10372 6.105
R38359 S.n10370 S.n10369 6.105
R38360 S.n10359 S.t615 6.105
R38361 S.n11122 S.t1469 6.105
R38362 S.n11134 S.n11133 6.105
R38363 S.n11137 S.n11136 6.105
R38364 S.n11119 S.t2414 6.105
R38365 S.n9333 S.t3801 6.105
R38366 S.n9344 S.n9343 6.105
R38367 S.n9341 S.n9340 6.105
R38368 S.n9330 S.t4045 6.105
R38369 S.n10082 S.t928 6.105
R38370 S.n10094 S.n10093 6.105
R38371 S.n10097 S.n10096 6.105
R38372 S.n10079 S.t1361 6.105
R38373 S.n8291 S.t2722 6.105
R38374 S.n8302 S.n8301 6.105
R38375 S.n8299 S.n8298 6.105
R38376 S.n8288 S.t3269 6.105
R38377 S.n9019 S.t4395 6.105
R38378 S.n9031 S.n9030 6.105
R38379 S.n9034 S.n9033 6.105
R38380 S.n9016 S.t850 6.105
R38381 S.n7227 S.t4084 6.105
R38382 S.n7238 S.n7237 6.105
R38383 S.n7235 S.n7234 6.105
R38384 S.n7224 S.t69 6.105
R38385 S.n7944 S.t1231 6.105
R38386 S.n7956 S.n7955 6.105
R38387 S.n7959 S.n7958 6.105
R38388 S.n7941 S.t2234 6.105
R38389 S.n6150 S.t3094 6.105
R38390 S.n6161 S.n6160 6.105
R38391 S.n6158 S.n6157 6.105
R38392 S.n6147 S.t3594 6.105
R38393 S.n6846 S.t220 6.105
R38394 S.n6858 S.n6857 6.105
R38395 S.n6861 S.n6860 6.105
R38396 S.n6843 S.t1133 6.105
R38397 S.n5050 S.t2041 6.105
R38398 S.n5061 S.n5060 6.105
R38399 S.n5058 S.n5057 6.105
R38400 S.n5047 S.t2519 6.105
R38401 S.n5736 S.t1770 6.105
R38402 S.n5748 S.n5747 6.105
R38403 S.n5751 S.n5750 6.105
R38404 S.n5733 S.t2681 6.105
R38405 S.n3938 S.t3584 6.105
R38406 S.n3949 S.n3948 6.105
R38407 S.n3946 S.n3945 6.105
R38408 S.n3935 S.t4053 6.105
R38409 S.n4601 S.t934 6.105
R38410 S.n4613 S.n4612 6.105
R38411 S.n4616 S.n4615 6.105
R38412 S.n4598 S.t1905 6.105
R38413 S.n2811 S.t3058 6.105
R38414 S.n2822 S.n2821 6.105
R38415 S.n2819 S.n2818 6.105
R38416 S.n2808 S.t3555 6.105
R38417 S.n3461 S.t4406 6.105
R38418 S.n3472 S.n3471 6.105
R38419 S.n3475 S.n3474 6.105
R38420 S.n3458 S.t863 6.105
R38421 S.n1639 S.t2011 6.105
R38422 S.n1651 S.n1650 6.105
R38423 S.n1648 S.n1647 6.105
R38424 S.n1636 S.t2492 6.105
R38425 S.n1406 S.t3388 6.105
R38426 S.n1407 S.t3126 6.105
R38427 S.n123 S.t795 6.105
R38428 S.n981 S.n980 6.105
R38429 S.n984 S.n983 6.105
R38430 S.n987 S.t1743 6.105
R38431 S.n13360 S.t1686 6.105
R38432 S.n13343 S.t2196 6.105
R38433 S.n13784 S.t3049 6.105
R38434 S.n13802 S.n13801 6.105
R38435 S.n13799 S.n13798 6.105
R38436 S.n13787 S.t3971 6.105
R38437 S.n12380 S.t637 6.105
R38438 S.n12391 S.n12390 6.105
R38439 S.n12388 S.n12387 6.105
R38440 S.n12383 S.t1095 6.105
R38441 S.n13122 S.t1999 6.105
R38442 S.n13139 S.n13138 6.105
R38443 S.n13142 S.n13141 6.105
R38444 S.n13125 S.t2953 6.105
R38445 S.n11386 S.t4062 6.105
R38446 S.n11397 S.n11396 6.105
R38447 S.n11394 S.n11393 6.105
R38448 S.n11389 S.t26 6.105
R38449 S.n12117 S.t941 6.105
R38450 S.n12134 S.n12133 6.105
R38451 S.n12137 S.n12136 6.105
R38452 S.n12120 S.t1912 6.105
R38453 S.n10379 S.t3287 6.105
R38454 S.n10390 S.n10389 6.105
R38455 S.n10387 S.n10386 6.105
R38456 S.n10382 S.t3565 6.105
R38457 S.n11085 S.t4416 6.105
R38458 S.n11102 S.n11101 6.105
R38459 S.n11105 S.n11104 6.105
R38460 S.n11088 S.t867 6.105
R38461 S.n9350 S.t2258 6.105
R38462 S.n9361 S.n9360 6.105
R38463 S.n9358 S.n9357 6.105
R38464 S.n9353 S.t2713 6.105
R38465 S.n10045 S.t3895 6.105
R38466 S.n10062 S.n10061 6.105
R38467 S.n10065 S.n10064 6.105
R38468 S.n10048 S.t4315 6.105
R38469 S.n8308 S.t3623 6.105
R38470 S.n8319 S.n8318 6.105
R38471 S.n8316 S.n8315 6.105
R38472 S.n8311 S.t4078 6.105
R38473 S.n8982 S.t764 6.105
R38474 S.n8999 S.n8998 6.105
R38475 S.n9002 S.n9001 6.105
R38476 S.n8985 S.t1715 6.105
R38477 S.n7244 S.t2539 6.105
R38478 S.n7255 S.n7254 6.105
R38479 S.n7252 S.n7251 6.105
R38480 S.n7247 S.t3089 6.105
R38481 S.n7907 S.t4187 6.105
R38482 S.n7924 S.n7923 6.105
R38483 S.n7927 S.n7926 6.105
R38484 S.n7910 S.t671 6.105
R38485 S.n6167 S.t1539 6.105
R38486 S.n6178 S.n6177 6.105
R38487 S.n6175 S.n6174 6.105
R38488 S.n6170 S.t2038 6.105
R38489 S.n6809 S.t3200 6.105
R38490 S.n6826 S.n6825 6.105
R38491 S.n6829 S.n6828 6.105
R38492 S.n6812 S.t4090 6.105
R38493 S.n5067 S.t482 6.105
R38494 S.n5078 S.n5077 6.105
R38495 S.n5075 S.n5074 6.105
R38496 S.n5070 S.t971 6.105
R38497 S.n5699 S.t432 6.105
R38498 S.n5716 S.n5715 6.105
R38499 S.n5719 S.n5718 6.105
R38500 S.n5702 S.t1378 6.105
R38501 S.n3955 S.t2031 6.105
R38502 S.n3966 S.n3965 6.105
R38503 S.n3963 S.n3962 6.105
R38504 S.n3958 S.t2510 6.105
R38505 S.n4564 S.t3900 6.105
R38506 S.n4581 S.n4580 6.105
R38507 S.n4584 S.n4583 6.105
R38508 S.n4567 S.t344 6.105
R38509 S.n2828 S.t1504 6.105
R38510 S.n2839 S.n2838 6.105
R38511 S.n2836 S.n2835 6.105
R38512 S.n2831 S.t2005 6.105
R38513 S.n3424 S.t2855 6.105
R38514 S.n3441 S.n3440 6.105
R38515 S.n3444 S.n3443 6.105
R38516 S.n3427 S.t3823 6.105
R38517 S.n1657 S.t453 6.105
R38518 S.n1668 S.n1667 6.105
R38519 S.n1665 S.n1664 6.105
R38520 S.n1660 S.t943 6.105
R38521 S.n2269 S.t1835 6.105
R38522 S.n2286 S.n2285 6.105
R38523 S.n2289 S.n2288 6.105
R38524 S.n2272 S.t2744 6.105
R38525 S.n632 S.t3909 6.105
R38526 S.n643 S.n642 6.105
R38527 S.n640 S.n639 6.105
R38528 S.n635 S.t4421 6.105
R38529 S.n615 S.t947 6.105
R38530 S.n626 S.n625 6.105
R38531 S.n623 S.n622 6.105
R38532 S.n618 S.t1471 6.105
R38533 S.n1250 S.t3532 6.105
R38534 S.n1242 S.t3038 6.105
R38535 S.n272 S.t923 6.105
R38536 S.n283 S.n282 6.105
R38537 S.n280 S.n279 6.105
R38538 S.n275 S.t1885 6.105
R38539 S.n2365 S.t1968 6.105
R38540 S.n2375 S.n2374 6.105
R38541 S.n2378 S.n2377 6.105
R38542 S.n2362 S.t2921 6.105
R38543 S.n10334 S.t3217 6.105
R38544 S.n10318 S.t3718 6.105
R38545 S.n10759 S.t4586 6.105
R38546 S.n10776 S.n10775 6.105
R38547 S.n10773 S.n10772 6.105
R38548 S.n10756 S.t990 6.105
R38549 S.n9295 S.t2182 6.105
R38550 S.n9306 S.n9305 6.105
R38551 S.n9303 S.n9302 6.105
R38552 S.n9292 S.t2635 6.105
R38553 S.n10147 S.t4012 6.105
R38554 S.n10159 S.n10158 6.105
R38555 S.n10162 S.n10161 6.105
R38556 S.n10144 S.t4481 6.105
R38557 S.n8255 S.t1082 6.105
R38558 S.n8266 S.n8265 6.105
R38559 S.n8263 S.n8262 6.105
R38560 S.n8252 S.t1649 6.105
R38561 S.n9080 S.t3007 6.105
R38562 S.n9092 S.n9091 6.105
R38563 S.n9095 S.n9094 6.105
R38564 S.n9077 S.t3941 6.105
R38565 S.n7191 S.t303 6.105
R38566 S.n7202 S.n7201 6.105
R38567 S.n7199 S.n7198 6.105
R38568 S.n7188 S.t588 6.105
R38569 S.n8005 S.t1960 6.105
R38570 S.n8017 S.n8016 6.105
R38571 S.n8020 S.n8019 6.105
R38572 S.n8002 S.t2908 6.105
R38573 S.n6114 S.t3782 6.105
R38574 S.n6125 S.n6124 6.105
R38575 S.n6122 S.n6121 6.105
R38576 S.n6111 S.t4245 6.105
R38577 S.n6907 S.t913 6.105
R38578 S.n6919 S.n6918 6.105
R38579 S.n6922 S.n6921 6.105
R38580 S.n6904 S.t1875 6.105
R38581 S.n5014 S.t643 6.105
R38582 S.n5025 S.n5024 6.105
R38583 S.n5022 S.n5021 6.105
R38584 S.n5011 S.t1101 6.105
R38585 S.n5797 S.t356 6.105
R38586 S.n5809 S.n5808 6.105
R38587 S.n5812 S.n5811 6.105
R38588 S.n5794 S.t1282 6.105
R38589 S.n3902 S.t2190 6.105
R38590 S.n3913 S.n3912 6.105
R38591 S.n3910 S.n3909 6.105
R38592 S.n3899 S.t2646 6.105
R38593 S.n4662 S.t3832 6.105
R38594 S.n4674 S.n4673 6.105
R38595 S.n4677 S.n4676 6.105
R38596 S.n4659 S.t265 6.105
R38597 S.n2775 S.t1661 6.105
R38598 S.n2786 S.n2785 6.105
R38599 S.n2783 S.n2782 6.105
R38600 S.n2772 S.t2165 6.105
R38601 S.n3521 S.t2761 6.105
R38602 S.n3532 S.n3531 6.105
R38603 S.n3535 S.n3534 6.105
R38604 S.n3518 S.t3746 6.105
R38605 S.n1602 S.t606 6.105
R38606 S.n1614 S.n1613 6.105
R38607 S.n1611 S.n1610 6.105
R38608 S.n1599 S.t1068 6.105
R38609 S.n1402 S.t1981 6.105
R38610 S.n1403 S.t1480 6.105
R38611 S.n1010 S.t3888 6.105
R38612 S.n1013 S.n1012 6.105
R38613 S.n1016 S.n1015 6.105
R38614 S.n1019 S.t324 6.105
R38615 S.n11358 S.t2660 6.105
R38616 S.n11341 S.t3213 6.105
R38617 S.n11786 S.t4030 6.105
R38618 S.n11804 S.n11803 6.105
R38619 S.n11801 S.n11800 6.105
R38620 S.n11789 S.t498 6.105
R38621 S.n10343 S.t1667 6.105
R38622 S.n10354 S.n10353 6.105
R38623 S.n10351 S.n10350 6.105
R38624 S.n10346 S.t2173 6.105
R38625 S.n11150 S.t3026 6.105
R38626 S.n11167 S.n11166 6.105
R38627 S.n11170 S.n11169 6.105
R38628 S.n11153 S.t3952 6.105
R38629 S.n9314 S.t620 6.105
R38630 S.n9325 S.n9324 6.105
R38631 S.n9322 S.n9321 6.105
R38632 S.n9317 S.t1080 6.105
R38633 S.n10110 S.t2475 6.105
R38634 S.n10127 S.n10126 6.105
R38635 S.n10130 S.n10129 6.105
R38636 S.n10113 S.t2927 6.105
R38637 S.n8272 S.t4276 6.105
R38638 S.n8283 S.n8282 6.105
R38639 S.n8280 S.n8279 6.105
R38640 S.n8275 S.t4603 6.105
R38641 S.n9043 S.t1448 6.105
R38642 S.n9060 S.n9059 6.105
R38643 S.n9063 S.n9062 6.105
R38644 S.n9046 S.t2402 6.105
R38645 S.n7208 S.t3274 6.105
R38646 S.n7219 S.n7218 6.105
R38647 S.n7216 S.n7215 6.105
R38648 S.n7211 S.t3779 6.105
R38649 S.n7968 S.t407 6.105
R38650 S.n7985 S.n7984 6.105
R38651 S.n7988 S.n7987 6.105
R38652 S.n7971 S.t1342 6.105
R38653 S.n6131 S.t84 6.105
R38654 S.n6142 S.n6141 6.105
R38655 S.n6139 S.n6138 6.105
R38656 S.n6134 S.t641 6.105
R38657 S.n6870 S.t1785 6.105
R38658 S.n6887 S.n6886 6.105
R38659 S.n6890 S.n6889 6.105
R38660 S.n6873 S.t2693 6.105
R38661 S.n5031 S.t3596 6.105
R38662 S.n5042 S.n5041 6.105
R38663 S.n5039 S.n5038 6.105
R38664 S.n5034 S.t4061 6.105
R38665 S.n5760 S.t3323 6.105
R38666 S.n5777 S.n5776 6.105
R38667 S.n5780 S.n5779 6.105
R38668 S.n5763 S.t4233 6.105
R38669 S.n3919 S.t633 6.105
R38670 S.n3930 S.n3929 6.105
R38671 S.n3927 S.n3926 6.105
R38672 S.n3922 S.t1085 6.105
R38673 S.n4625 S.t2295 6.105
R38674 S.n4642 S.n4641 6.105
R38675 S.n4645 S.n4644 6.105
R38676 S.n4628 S.t3244 6.105
R38677 S.n2792 S.t15 6.105
R38678 S.n2803 S.n2802 6.105
R38679 S.n2800 S.n2799 6.105
R38680 S.n2795 S.t600 6.105
R38681 S.n3484 S.t1458 6.105
R38682 S.n3501 S.n3500 6.105
R38683 S.n3504 S.n3503 6.105
R38684 S.n3487 S.t2410 6.105
R38685 S.n1620 S.t3559 6.105
R38686 S.n1631 S.n1630 6.105
R38687 S.n1628 S.n1627 6.105
R38688 S.n1623 S.t4034 6.105
R38689 S.n2328 S.t416 6.105
R38690 S.n2345 S.n2344 6.105
R38691 S.n2348 S.n2347 6.105
R38692 S.n2331 S.t1356 6.105
R38693 S.n597 S.t2498 6.105
R38694 S.n608 S.n607 6.105
R38695 S.n605 S.n604 6.105
R38696 S.n600 S.t3031 6.105
R38697 S.n580 S.t4041 6.105
R38698 S.n591 S.n590 6.105
R38699 S.n588 S.n587 6.105
R38700 S.n583 S.t4587 6.105
R38701 S.n1237 S.t2141 6.105
R38702 S.n1229 S.t1644 6.105
R38703 S.n243 S.t3812 6.105
R38704 S.n251 S.n250 6.105
R38705 S.n222 S.n221 6.105
R38706 S.n246 S.t244 6.105
R38707 S.n2424 S.t338 6.105
R38708 S.n2434 S.n2433 6.105
R38709 S.n2437 S.n2436 6.105
R38710 S.n2421 S.t1261 6.105
R38711 S.n8227 S.t4190 6.105
R38712 S.n8211 S.t217 6.105
R38713 S.n8656 S.t1605 6.105
R38714 S.n8673 S.n8672 6.105
R38715 S.n8670 S.n8669 6.105
R38716 S.n8653 S.t2521 6.105
R38717 S.n7153 S.t3202 6.105
R38718 S.n7164 S.n7163 6.105
R38719 S.n7161 S.n7160 6.105
R38720 S.n7150 S.t3699 6.105
R38721 S.n8070 S.t550 6.105
R38722 S.n8082 S.n8081 6.105
R38723 S.n8085 S.n8084 6.105
R38724 S.n8067 S.t1519 6.105
R38725 S.n6078 S.t2157 6.105
R38726 S.n6089 S.n6088 6.105
R38727 S.n6086 S.n6085 6.105
R38728 S.n6075 S.t2612 6.105
R38729 S.n6968 S.t4000 6.105
R38730 S.n6980 S.n6979 6.105
R38731 S.n6983 S.n6982 6.105
R38732 S.n6965 S.t461 6.105
R38733 S.n4978 S.t1302 6.105
R38734 S.n4989 S.n4988 6.105
R38735 S.n4986 S.n4985 6.105
R38736 S.n4975 S.t1626 6.105
R38737 S.n5858 S.t1024 6.105
R38738 S.n5870 S.n5869 6.105
R38739 S.n5873 S.n5872 6.105
R38740 S.n5855 S.t2007 6.105
R38741 S.n3866 S.t2858 6.105
R38742 S.n3877 S.n3876 6.105
R38743 S.n3874 S.n3873 6.105
R38744 S.n3863 S.t3378 6.105
R38745 S.n4723 S.t4538 6.105
R38746 S.n4735 S.n4734 6.105
R38747 S.n4738 S.n4737 6.105
R38748 S.n4720 S.t945 6.105
R38749 S.n2739 S.t234 6.105
R38750 S.n2750 S.n2749 6.105
R38751 S.n2747 S.n2746 6.105
R38752 S.n2736 S.t749 6.105
R38753 S.n3581 S.t1366 6.105
R38754 S.n3592 S.n3591 6.105
R38755 S.n3595 S.n3594 6.105
R38756 S.n3578 S.t2348 6.105
R38757 S.n1565 S.t3715 6.105
R38758 S.n1577 S.n1576 6.105
R38759 S.n1574 S.n1573 6.105
R38760 S.n1562 S.t4174 6.105
R38761 S.n1398 S.t581 6.105
R38762 S.n1399 S.t4598 6.105
R38763 S.n1042 S.t2469 6.105
R38764 S.n1045 S.n1044 6.105
R38765 S.n1048 S.n1047 6.105
R38766 S.n1051 S.t3432 6.105
R38767 S.n9286 S.t3725 6.105
R38768 S.n9269 S.t4183 6.105
R38769 S.n9718 S.t1045 6.105
R38770 S.n9736 S.n9735 6.105
R38771 S.n9733 S.n9732 6.105
R38772 S.n9721 S.t1534 6.105
R38773 S.n8236 S.t2641 6.105
R38774 S.n8247 S.n8246 6.105
R38775 S.n8244 S.n8243 6.105
R38776 S.n8239 S.t3198 6.105
R38777 S.n9108 S.t4565 6.105
R38778 S.n9125 S.n9124 6.105
R38779 S.n9128 S.n9127 6.105
R38780 S.n9111 S.t973 6.105
R38781 S.n7172 S.t1652 6.105
R38782 S.n7183 S.n7182 6.105
R38783 S.n7180 S.n7179 6.105
R38784 S.n7175 S.t2153 6.105
R38785 S.n8033 S.t3509 6.105
R38786 S.n8050 S.n8049 6.105
R38787 S.n8053 S.n8052 6.105
R38788 S.n8036 S.t4464 6.105
R38789 S.n6095 S.t819 6.105
R38790 S.n6106 S.n6105 6.105
R38791 S.n6103 S.n6102 6.105
R38792 S.n6098 S.t1059 6.105
R38793 S.n6931 S.t2457 6.105
R38794 S.n6948 S.n6947 6.105
R38795 S.n6951 S.n6950 6.105
R38796 S.n6934 S.t3420 6.105
R38797 S.n4995 S.t4255 6.105
R38798 S.n5006 S.n5005 6.105
R38799 S.n5003 S.n5002 6.105
R38800 S.n4998 S.t283 6.105
R38801 S.n5821 S.t3988 6.105
R38802 S.n5838 S.n5837 6.105
R38803 S.n5841 S.n5840 6.105
R38804 S.n5824 S.t451 6.105
R38805 S.n3883 S.t3737 6.105
R38806 S.n3894 S.n3893 6.105
R38807 S.n3891 S.n3890 6.105
R38808 S.n3886 S.t4194 6.105
R38809 S.n4686 S.t869 6.105
R38810 S.n4703 S.n4702 6.105
R38811 S.n4706 S.n4705 6.105
R38812 S.n4689 S.t1830 6.105
R38813 S.n2756 S.t3210 6.105
R38814 S.n2767 S.n2766 6.105
R38815 S.n2764 S.n2763 6.105
R38816 S.n2759 S.t3705 6.105
R38817 S.n3544 S.t4318 6.105
R38818 S.n3561 S.n3560 6.105
R38819 S.n3564 S.n3563 6.105
R38820 S.n3547 S.t793 6.105
R38821 S.n1583 S.t2168 6.105
R38822 S.n1594 S.n1593 6.105
R38823 S.n1591 S.n1590 6.105
R38824 S.n1586 S.t2622 6.105
R38825 S.n2387 S.t3304 6.105
R38826 S.n2404 S.n2403 6.105
R38827 S.n2407 S.n2406 6.105
R38828 S.n2390 S.t4213 6.105
R38829 S.n562 S.t1073 6.105
R38830 S.n573 S.n572 6.105
R38831 S.n570 S.n569 6.105
R38832 S.n565 S.t1635 6.105
R38833 S.n545 S.t2629 6.105
R38834 S.n556 S.n555 6.105
R38835 S.n553 S.n552 6.105
R38836 S.n548 S.t3187 6.105
R38837 S.n1224 S.t733 6.105
R38838 S.n1216 S.t211 6.105
R38839 S.n208 S.t2405 6.105
R38840 S.n219 S.n218 6.105
R38841 S.n216 S.n215 6.105
R38842 S.n211 S.t3357 6.105
R38843 S.n2483 S.t1009 6.105
R38844 S.n2493 S.n2492 6.105
R38845 S.n2496 S.n2495 6.105
R38846 S.n2480 S.t1985 6.105
R38847 S.n6050 S.t745 6.105
R38848 S.n6034 S.t1209 6.105
R38849 S.n6483 S.t2584 6.105
R38850 S.n6500 S.n6499 6.105
R38851 S.n6497 S.n6496 6.105
R38852 S.n6480 S.t3571 6.105
R38853 S.n4940 S.t4169 6.105
R38854 S.n4951 S.n4950 6.105
R38855 S.n4948 S.n4947 6.105
R38856 S.n4937 S.t196 6.105
R38857 S.n5923 S.t4117 6.105
R38858 S.n5935 S.n5934 6.105
R38859 S.n5938 S.n5937 6.105
R38860 S.n5920 S.t603 6.105
R38861 S.n3830 S.t1202 6.105
R38862 S.n3841 S.n3840 6.105
R38863 S.n3838 S.n3837 6.105
R38864 S.n3827 S.t1751 6.105
R38865 S.n4784 S.t3136 6.105
R38866 S.n4796 S.n4795 6.105
R38867 S.n4799 S.n4798 6.105
R38868 S.n4781 S.t4037 6.105
R38869 S.n2703 S.t924 6.105
R38870 S.n2714 S.n2713 6.105
R38871 S.n2711 S.n2710 6.105
R38872 S.n2700 S.t1172 6.105
R38873 S.n3641 S.t2088 6.105
R38874 S.n3652 S.n3651 6.105
R38875 S.n3655 S.n3654 6.105
R38876 S.n3638 S.t3035 6.105
R38877 S.n1528 S.t4389 6.105
R38878 S.n1540 S.n1539 6.105
R38879 S.n1537 S.n1536 6.105
R38880 S.n1525 S.t393 6.105
R38881 S.n1394 S.t3690 6.105
R38882 S.n1395 S.t3192 6.105
R38883 S.n1074 S.t854 6.105
R38884 S.n1077 S.n1076 6.105
R38885 S.n1080 S.n1079 6.105
R38886 S.n1083 S.t1812 6.105
R38887 S.n7144 S.t223 6.105
R38888 S.n7127 S.t742 6.105
R38889 S.n7580 S.t2114 6.105
R38890 S.n7598 S.n7597 6.105
R38891 S.n7595 S.n7594 6.105
R38892 S.n7583 S.t3067 6.105
R38893 S.n6059 S.t3702 6.105
R38894 S.n6070 S.n6069 6.105
R38895 S.n6067 S.n6066 6.105
R38896 S.n6062 S.t4162 6.105
R38897 S.n6996 S.t1034 6.105
R38898 S.n7013 S.n7012 6.105
R38899 S.n7016 S.n7015 6.105
R38900 S.n6999 S.t2021 6.105
R38901 S.n4959 S.t2618 6.105
R38902 S.n4970 S.n4969 6.105
R38903 S.n4967 S.n4966 6.105
R38904 S.n4962 S.t3178 6.105
R38905 S.n5886 S.t2574 6.105
R38906 S.n5903 S.n5902 6.105
R38907 S.n5906 S.n5905 6.105
R38908 S.n5889 S.t3557 6.105
R38909 S.n3847 S.t4410 6.105
R38910 S.n3858 S.n3857 6.105
R38911 S.n3855 S.n3854 6.105
R38912 S.n3850 S.t180 6.105
R38913 S.n4747 S.t1580 6.105
R38914 S.n4764 S.n4763 6.105
R38915 S.n4767 S.n4766 6.105
R38916 S.n4750 S.t2496 6.105
R38917 S.n2720 S.t3889 6.105
R38918 S.n2731 S.n2730 6.105
R38919 S.n2728 S.n2727 6.105
R38920 S.n2723 S.t4381 6.105
R38921 S.n3604 S.t520 6.105
R38922 S.n3621 S.n3620 6.105
R38923 S.n3624 S.n3623 6.105
R38924 S.n3607 S.t1478 6.105
R38925 S.n1546 S.t760 6.105
R38926 S.n1557 S.n1556 6.105
R38927 S.n1554 S.n1553 6.105
R38928 S.n1549 S.t1220 6.105
R38929 S.n2446 S.t1898 6.105
R38930 S.n2463 S.n2462 6.105
R38931 S.n2466 S.n2465 6.105
R38932 S.n2449 S.t2829 6.105
R38933 S.n527 S.t4179 6.105
R38934 S.n538 S.n537 6.105
R38935 S.n535 S.n534 6.105
R38936 S.n530 S.t208 6.105
R38937 S.n510 S.t1229 6.105
R38938 S.n521 S.n520 6.105
R38939 S.n518 S.n517 6.105
R38940 S.n513 S.t1775 6.105
R38941 S.n1211 S.t1411 6.105
R38942 S.n1203 S.t908 6.105
R38943 S.n176 S.t3114 6.105
R38944 S.n187 S.n186 6.105
R38945 S.n184 S.n183 6.105
R38946 S.n179 S.t4020 6.105
R38947 S.n2542 S.t4098 6.105
R38948 S.n2552 S.n2551 6.105
R38949 S.n2555 S.n2554 6.105
R38950 S.n2539 S.t583 6.105
R38951 S.n3802 S.t4321 6.105
R38952 S.n3786 S.t334 6.105
R38953 S.n4238 S.t1722 6.105
R38954 S.n4255 S.n4254 6.105
R38955 S.n4252 S.n4251 6.105
R38956 S.n4235 S.t2625 6.105
R38957 S.n2665 S.t3814 6.105
R38958 S.n2676 S.n2675 6.105
R38959 S.n2673 S.n2672 6.105
R38960 S.n2662 S.t4291 6.105
R38961 S.n3705 S.t677 6.105
R38962 S.n3716 S.n3715 6.105
R38963 S.n3719 S.n3718 6.105
R38964 S.n3702 S.t1639 6.105
R38965 S.n1491 S.t2740 6.105
R38966 S.n1503 S.n1502 6.105
R38967 S.n1500 S.n1499 6.105
R38968 S.n1488 S.t3281 6.105
R38969 S.n1390 S.t2297 6.105
R38970 S.n1391 S.t1779 6.105
R38971 S.n1106 S.t1563 6.105
R38972 S.n1109 S.n1108 6.105
R38973 S.n1112 S.n1111 6.105
R38974 S.n1115 S.t2479 6.105
R38975 S.n4931 S.t1215 6.105
R38976 S.n4914 S.t1765 6.105
R38977 S.n5371 S.t1163 6.105
R38978 S.n5389 S.n5388 6.105
R38979 S.n5386 S.n5385 6.105
R38980 S.n5374 S.t2167 6.105
R38981 S.n3811 S.t2765 6.105
R38982 S.n3822 S.n3821 6.105
R38983 S.n3819 S.n3818 6.105
R38984 S.n3814 S.t3300 6.105
R38985 S.n4812 S.t135 6.105
R38986 S.n4829 S.n4828 6.105
R38987 S.n4832 S.n4831 6.105
R38988 S.n4815 S.t1071 6.105
R38989 S.n2684 S.t2273 6.105
R38990 S.n2695 S.n2694 6.105
R38991 S.n2692 S.n2691 6.105
R38992 S.n2687 S.t2732 6.105
R38993 S.n3668 S.t3638 6.105
R38994 S.n3685 S.n3684 6.105
R38995 S.n3688 S.n3687 6.105
R38996 S.n3671 S.t4595 6.105
R38997 S.n1509 S.t1440 6.105
R38998 S.n1520 S.n1519 6.105
R38999 S.n1517 S.n1516 6.105
R39000 S.n1512 S.t1729 6.105
R39001 S.n2505 S.t2557 6.105
R39002 S.n2522 S.n2521 6.105
R39003 S.n2525 S.n2524 6.105
R39004 S.n2508 S.t3535 6.105
R39005 S.n492 S.t398 6.105
R39006 S.n503 S.n502 6.105
R39007 S.n500 S.n499 6.105
R39008 S.n495 S.t904 6.105
R39009 S.n475 S.t1954 6.105
R39010 S.n486 S.n485 6.105
R39011 S.n483 S.n482 6.105
R39012 S.n478 S.t2251 6.105
R39013 S.n1198 S.t4267 6.105
R39014 S.n1190 S.t3798 6.105
R39015 S.n144 S.t1704 6.105
R39016 S.n155 S.n154 6.105
R39017 S.n152 S.n151 6.105
R39018 S.n147 S.t2607 6.105
R39019 S.n1944 S.t2701 6.105
R39020 S.n1959 S.n1958 6.105
R39021 S.n1956 S.n1955 6.105
R39022 S.n1941 S.t3692 6.105
R39023 S.n1463 S.t1348 6.105
R39024 S.n1446 S.t1876 6.105
R39025 S.n1386 S.t2714 6.105
R39026 S.n1387 S.t2453 6.105
R39027 S.n1144 S.t110 6.105
R39028 S.n1147 S.n1146 6.105
R39029 S.n1150 S.n1149 6.105
R39030 S.n1153 S.t1053 6.105
R39031 S.n2656 S.t856 6.105
R39032 S.n2639 S.t1343 6.105
R39033 S.n3101 S.t2238 6.105
R39034 S.n3119 S.n3118 6.105
R39035 S.n3116 S.n3115 6.105
R39036 S.n3104 S.t3190 6.105
R39037 S.n1472 S.t4295 6.105
R39038 S.n1483 S.n1482 6.105
R39039 S.n1480 S.n1479 6.105
R39040 S.n1475 S.t312 6.105
R39041 S.n2568 S.t1146 6.105
R39042 S.n2585 S.n2584 6.105
R39043 S.n2588 S.n2587 6.105
R39044 S.n2571 S.t2147 6.105
R39045 S.n457 S.t3288 6.105
R39046 S.n468 S.n467 6.105
R39047 S.n465 S.n464 6.105
R39048 S.n460 S.t3793 6.105
R39049 S.n441 S.t318 6.105
R39050 S.n452 S.n451 6.105
R39051 S.n449 S.n448 6.105
R39052 S.n444 S.t829 6.105
R39053 S.n1382 S.t1319 6.105
R39054 S.n1383 S.t836 6.105
R39055 S.n931 S.t3259 6.105
R39056 S.n944 S.n943 6.105
R39057 S.n947 S.n946 6.105
R39058 S.n934 S.t4157 6.105
R39059 S.n435 S.t1878 6.105
R39060 S.n417 S.t2385 6.105
R39061 S.n1428 S.t2571 6.105
R39062 S.n22309 S.t4257 6.105
R39063 S.n22312 S.n22311 6.105
R39064 S.n21974 S.t3768 6.105
R39065 S.n22996 S.t860 6.105
R39066 S.n22759 S.t297 6.105
R39067 S.n22767 S.n22766 6.105
R39068 S.n22770 S.n22769 6.105
R39069 S.n22762 S.t2549 6.105
R39070 S.n21322 S.t2080 6.105
R39071 S.n21333 S.n21332 6.105
R39072 S.n21330 S.n21329 6.105
R39073 S.n21325 S.t4147 6.105
R39074 S.n22302 S.t1308 6.105
R39075 S.n22305 S.n22304 6.105
R39076 S.n22335 S.t3996 6.105
R39077 S.n22338 S.n22337 6.105
R39078 S.n22330 S.t1301 6.105
R39079 S.n22315 S.n22314 6.105
R39080 S.n22280 S.n22278 4.263
R39081 S.n965 S.n964 3.857
R39082 S.n1906 S.n1905 3.857
R39083 S.n2606 S.n2605 3.857
R39084 S.n3737 S.n3736 3.857
R39085 S.n4850 S.n4849 3.857
R39086 S.n5955 S.n5954 3.857
R39087 S.n7033 S.n7032 3.857
R39088 S.n8102 S.n8101 3.857
R39089 S.n9145 S.n9144 3.857
R39090 S.n10179 S.n10178 3.857
R39091 S.n11187 S.n11186 3.857
R39092 S.n12186 S.n12185 3.857
R39093 S.n13159 S.n13158 3.857
R39094 S.n14123 S.n14122 3.857
R39095 S.n15061 S.n15060 3.857
R39096 S.n15990 S.n15989 3.857
R39097 S.n16893 S.n16892 3.857
R39098 S.n17787 S.n17786 3.857
R39099 S.n18655 S.n18654 3.857
R39100 S.n19512 S.n19511 3.857
R39101 S.n21162 S.n21161 3.857
R39102 S.n21180 S.n21179 3.857
R39103 S.n22778 S.n22777 3.857
R39104 S.n22802 S.n22799 0.178
R39105 S.n1180 S.n1177 0.164
R39106 S.n23011 S.n23010 0.144
R39107 S.n962 S.n961 0.136
R39108 S.n5437 S.n5436 0.133
R39109 S.n1441 S.n1433 0.123
R39110 S.n105 S.n83 0.123
R39111 S.n992 S.n115 0.123
R39112 S.n1024 S.n1002 0.123
R39113 S.n1056 S.n1034 0.123
R39114 S.n1088 S.n1066 0.123
R39115 S.n1120 S.n1098 0.123
R39116 S.n1158 S.n1130 0.123
R39117 S.n1271 S.n1270 0.123
R39118 S.n1258 S.n1257 0.123
R39119 S.n1245 S.n1244 0.123
R39120 S.n1232 S.n1231 0.123
R39121 S.n1219 S.n1218 0.123
R39122 S.n1206 S.n1205 0.123
R39123 S.n1193 S.n1192 0.123
R39124 S.n1170 S.n1168 0.123
R39125 S.n967 S.n966 0.117
R39126 S.n2608 S.n2607 0.117
R39127 S.n3739 S.n3738 0.117
R39128 S.n4852 S.n4851 0.117
R39129 S.n5957 S.n5956 0.117
R39130 S.n7035 S.n7034 0.117
R39131 S.n8104 S.n8103 0.117
R39132 S.n9147 S.n9146 0.117
R39133 S.n10181 S.n10180 0.117
R39134 S.n11189 S.n11188 0.117
R39135 S.n12188 S.n12187 0.117
R39136 S.n13161 S.n13160 0.117
R39137 S.n14125 S.n14124 0.117
R39138 S.n15063 S.n15062 0.117
R39139 S.n15992 S.n15991 0.117
R39140 S.n16895 S.n16894 0.117
R39141 S.n17789 S.n17788 0.117
R39142 S.n18657 S.n18656 0.117
R39143 S.n19514 S.n19513 0.117
R39144 S.n21164 S.n21163 0.117
R39145 S.n21182 S.n21181 0.117
R39146 S.n22780 S.n22779 0.117
R39147 S.n23031 S.n3729 0.116
R39148 S.n23030 S.n4842 0.114
R39149 S.n23032 S.n2598 0.113
R39150 S.n23011 S.n22791 0.11
R39151 S.n23013 S.n21172 0.11
R39152 S.n23014 S.n20344 0.11
R39153 S.n23015 S.n19504 0.11
R39154 S.n23016 S.n18647 0.11
R39155 S.n23017 S.n17779 0.11
R39156 S.n23018 S.n16885 0.11
R39157 S.n23019 S.n15982 0.11
R39158 S.n23020 S.n15053 0.11
R39159 S.n23021 S.n14115 0.11
R39160 S.n23022 S.n13151 0.11
R39161 S.n23023 S.n12178 0.11
R39162 S.n23024 S.n11179 0.11
R39163 S.n23025 S.n10171 0.11
R39164 S.n23026 S.n9137 0.11
R39165 S.n23027 S.n8094 0.11
R39166 S.n23028 S.n7025 0.11
R39167 S.n23029 S.n5947 0.11
R39168 S.n23012 S.n21980 0.11
R39169 S.n22812 S.n22811 0.109
R39170 S.n20471 S.n20469 0.109
R39171 S.n19860 S.n19858 0.109
R39172 S.n19006 S.n19004 0.109
R39173 S.n18140 S.n18138 0.109
R39174 S.n17251 S.n17249 0.109
R39175 S.n16349 S.n16347 0.109
R39176 S.n15425 S.n15423 0.109
R39177 S.n14488 S.n14486 0.109
R39178 S.n13529 S.n13527 0.109
R39179 S.n12557 S.n12555 0.109
R39180 S.n11563 S.n11561 0.109
R39181 S.n10556 S.n10554 0.109
R39182 S.n9527 S.n9525 0.109
R39183 S.n8485 S.n8483 0.109
R39184 S.n7421 S.n7419 0.109
R39185 S.n6344 S.n6342 0.109
R39186 S.n5244 S.n5242 0.109
R39187 S.n3005 S.n3003 0.109
R39188 S.n1834 S.n1831 0.109
R39189 S.n388 S.n383 0.104
R39190 S.n356 S.n351 0.104
R39191 S.n324 S.n319 0.104
R39192 S.n292 S.n287 0.104
R39193 S.n260 S.n255 0.104
R39194 S.n231 S.n226 0.104
R39195 S.n196 S.n191 0.104
R39196 S.n164 S.n159 0.104
R39197 S.n132 S.n127 0.104
R39198 S.n2603 S.n2602 0.103
R39199 S.n3734 S.n3733 0.103
R39200 S.n4847 S.n4846 0.103
R39201 S.n5952 S.n5951 0.103
R39202 S.n7030 S.n7029 0.103
R39203 S.n8099 S.n8098 0.103
R39204 S.n9142 S.n9141 0.103
R39205 S.n10176 S.n10175 0.103
R39206 S.n11184 S.n11183 0.103
R39207 S.n12183 S.n12182 0.103
R39208 S.n13156 S.n13155 0.103
R39209 S.n14120 S.n14119 0.103
R39210 S.n15058 S.n15057 0.103
R39211 S.n15987 S.n15986 0.103
R39212 S.n16890 S.n16889 0.103
R39213 S.n17784 S.n17783 0.103
R39214 S.n18652 S.n18651 0.103
R39215 S.n19509 S.n19508 0.103
R39216 S.n21159 S.n21158 0.103
R39217 S.n21177 S.n21176 0.103
R39218 S.n22787 S.n22786 0.103
R39219 S.n1929 S.n1928 0.097
R39220 S.n2008 S.n2007 0.097
R39221 S.n387 S.n384 0.097
R39222 S.n355 S.n352 0.097
R39223 S.n323 S.n320 0.097
R39224 S.n291 S.n288 0.097
R39225 S.n259 S.n256 0.097
R39226 S.n230 S.n227 0.097
R39227 S.n195 S.n192 0.097
R39228 S.n163 S.n160 0.097
R39229 S.n131 S.n128 0.097
R39230 S.n22274 S.n22273 0.093
R39231 S.n21284 S.n21283 0.093
R39232 S.n20459 S.n20458 0.093
R39233 S.n19848 S.n19847 0.093
R39234 S.n18067 S.n18065 0.093
R39235 S.n17178 S.n17176 0.093
R39236 S.n16240 S.n16238 0.093
R39237 S.n15316 S.n15314 0.093
R39238 S.n14343 S.n14341 0.093
R39239 S.n13384 S.n13382 0.093
R39240 S.n12376 S.n12374 0.093
R39241 S.n11382 S.n11380 0.093
R39242 S.n10339 S.n10337 0.093
R39243 S.n9310 S.n9308 0.093
R39244 S.n8232 S.n8230 0.093
R39245 S.n7168 S.n7166 0.093
R39246 S.n6055 S.n6053 0.093
R39247 S.n4955 S.n4953 0.093
R39248 S.n3807 S.n3805 0.093
R39249 S.n2680 S.n2678 0.093
R39250 S.n1468 S.n1466 0.093
R39251 S.n910 S.n906 0.092
R39252 S.n22297 S.n22296 0.092
R39253 S.n22319 S.n22318 0.092
R39254 S.n19838 S.n19837 0.091
R39255 S.n18986 S.n18985 0.091
R39256 S S.n23033 0.09
R39257 S.n2076 S.n2075 0.087
R39258 S.n972 S.n971 0.082
R39259 S.n1912 S.n1911 0.082
R39260 S.n2613 S.n2612 0.082
R39261 S.n3744 S.n3743 0.082
R39262 S.n4857 S.n4856 0.082
R39263 S.n5962 S.n5961 0.082
R39264 S.n7040 S.n7039 0.082
R39265 S.n8109 S.n8108 0.082
R39266 S.n9152 S.n9151 0.082
R39267 S.n10186 S.n10185 0.082
R39268 S.n11194 S.n11193 0.082
R39269 S.n12193 S.n12192 0.082
R39270 S.n13166 S.n13165 0.082
R39271 S.n14130 S.n14129 0.082
R39272 S.n15068 S.n15067 0.082
R39273 S.n15997 S.n15996 0.082
R39274 S.n16900 S.n16899 0.082
R39275 S.n17794 S.n17793 0.082
R39276 S.n18662 S.n18661 0.082
R39277 S.n19519 S.n19518 0.082
R39278 S.n21169 S.n21168 0.082
R39279 S.n21187 S.n21186 0.082
R39280 S.n22789 S.n22784 0.082
R39281 S.n2010 S.n2009 0.08
R39282 S.n22804 S.n22803 0.079
R39283 S.n805 S.n804 0.077
R39284 S.n1810 S.n1809 0.077
R39285 S.n2972 S.n2971 0.077
R39286 S.n4099 S.n4098 0.077
R39287 S.n5211 S.n5210 0.077
R39288 S.n6311 S.n6310 0.077
R39289 S.n7388 S.n7387 0.077
R39290 S.n8452 S.n8451 0.077
R39291 S.n9494 S.n9493 0.077
R39292 S.n10523 S.n10522 0.077
R39293 S.n11530 S.n11529 0.077
R39294 S.n12524 S.n12523 0.077
R39295 S.n13496 S.n13495 0.077
R39296 S.n14455 S.n14454 0.077
R39297 S.n15392 S.n15391 0.077
R39298 S.n16316 S.n16315 0.077
R39299 S.n17218 S.n17217 0.077
R39300 S.n18107 S.n18106 0.077
R39301 S.n18972 S.n18971 0.077
R39302 S.n19824 S.n19823 0.077
R39303 S.n766 S.n765 0.077
R39304 S.n785 S.n784 0.077
R39305 S.n20450 S.n20449 0.076
R39306 S.n22287 S.n22286 0.074
R39307 S.n19812 S.n19811 0.074
R39308 S.n21294 S.n21293 0.074
R39309 S.n18942 S.n18941 0.074
R39310 S.n18057 S.n18056 0.074
R39311 S.n17150 S.n17149 0.074
R39312 S.n16230 S.n16229 0.074
R39313 S.n15288 S.n15287 0.074
R39314 S.n14333 S.n14332 0.074
R39315 S.n13356 S.n13355 0.074
R39316 S.n12366 S.n12365 0.074
R39317 S.n11354 S.n11353 0.074
R39318 S.n10329 S.n10328 0.074
R39319 S.n9282 S.n9281 0.074
R39320 S.n8222 S.n8221 0.074
R39321 S.n7140 S.n7139 0.074
R39322 S.n6045 S.n6044 0.074
R39323 S.n4927 S.n4926 0.074
R39324 S.n3797 S.n3796 0.074
R39325 S.n1458 S.n1457 0.074
R39326 S.n2652 S.n2651 0.074
R39327 S.n430 S.n429 0.074
R39328 S.n22953 S.n22952 0.073
R39329 S.n22961 S.n22960 0.073
R39330 S.n22946 S.n22945 0.073
R39331 S.n22939 S.n22938 0.073
R39332 S.n22932 S.n22931 0.073
R39333 S.n22925 S.n22924 0.073
R39334 S.n22918 S.n22917 0.073
R39335 S.n22911 S.n22910 0.073
R39336 S.n22904 S.n22903 0.073
R39337 S.n22897 S.n22896 0.073
R39338 S.n22890 S.n22889 0.073
R39339 S.n22883 S.n22882 0.073
R39340 S.n22876 S.n22875 0.073
R39341 S.n22869 S.n22868 0.073
R39342 S.n22862 S.n22861 0.073
R39343 S.n22855 S.n22854 0.073
R39344 S.n22848 S.n22847 0.073
R39345 S.n22841 S.n22840 0.073
R39346 S.n22832 S.n22831 0.073
R39347 S.n22823 S.n22822 0.073
R39348 S.n1450 S.n1449 0.072
R39349 S.n22967 S.n22966 0.071
R39350 S.n22969 S.n22968 0.071
R39351 S.t41 S.n22835 0.068
R39352 S.t41 S.n22826 0.068
R39353 S.t41 S.n22808 0.068
R39354 S.n21169 S.n21156 0.067
R39355 S.n21169 S.n21155 0.067
R39356 S.n19519 S.n19506 0.067
R39357 S.n19519 S.n19505 0.067
R39358 S.n18662 S.n18649 0.067
R39359 S.n18662 S.n18648 0.067
R39360 S.n17794 S.n17781 0.067
R39361 S.n17794 S.n17780 0.067
R39362 S.n16900 S.n16887 0.067
R39363 S.n16900 S.n16886 0.067
R39364 S.n15997 S.n15984 0.067
R39365 S.n15997 S.n15983 0.067
R39366 S.n15068 S.n15055 0.067
R39367 S.n15068 S.n15054 0.067
R39368 S.n14130 S.n14117 0.067
R39369 S.n14130 S.n14116 0.067
R39370 S.n13166 S.n13153 0.067
R39371 S.n13166 S.n13152 0.067
R39372 S.n12193 S.n12180 0.067
R39373 S.n12193 S.n12179 0.067
R39374 S.n11194 S.n11181 0.067
R39375 S.n11194 S.n11180 0.067
R39376 S.n10186 S.n10173 0.067
R39377 S.n10186 S.n10172 0.067
R39378 S.n9152 S.n9139 0.067
R39379 S.n9152 S.n9138 0.067
R39380 S.n8109 S.n8096 0.067
R39381 S.n8109 S.n8095 0.067
R39382 S.n7040 S.n7027 0.067
R39383 S.n7040 S.n7026 0.067
R39384 S.n5962 S.n5949 0.067
R39385 S.n5962 S.n5948 0.067
R39386 S.n4857 S.n4844 0.067
R39387 S.n4857 S.n4843 0.067
R39388 S.n3744 S.n3731 0.067
R39389 S.n3744 S.n3730 0.067
R39390 S.n2613 S.n2600 0.067
R39391 S.n2613 S.n2599 0.067
R39392 S.n972 S.n959 0.067
R39393 S.n972 S.n957 0.067
R39394 S.n1425 S.n1424 0.067
R39395 S.n1304 S.n1302 0.067
R39396 S.n1304 S.n1303 0.067
R39397 S.n1342 S.n1341 0.067
R39398 S.n1342 S.n1340 0.067
R39399 S.n1376 S.n1374 0.067
R39400 S.n1376 S.n1375 0.067
R39401 S.n45 S.n28 0.067
R39402 S.n45 S.n27 0.067
R39403 S.n1291 S.n1289 0.067
R39404 S.n1291 S.n1290 0.067
R39405 S.n76 S.n75 0.067
R39406 S.n76 S.n74 0.067
R39407 S.n1279 S.n1277 0.067
R39408 S.n1279 S.n1278 0.067
R39409 S.n108 S.n107 0.067
R39410 S.n108 S.n106 0.067
R39411 S.n1266 S.n1264 0.067
R39412 S.n1266 S.n1265 0.067
R39413 S.n995 S.n994 0.067
R39414 S.n995 S.n993 0.067
R39415 S.n1253 S.n1251 0.067
R39416 S.n1253 S.n1252 0.067
R39417 S.n1027 S.n1026 0.067
R39418 S.n1027 S.n1025 0.067
R39419 S.n1240 S.n1238 0.067
R39420 S.n1240 S.n1239 0.067
R39421 S.n1059 S.n1058 0.067
R39422 S.n1059 S.n1057 0.067
R39423 S.n1227 S.n1225 0.067
R39424 S.n1227 S.n1226 0.067
R39425 S.n1091 S.n1090 0.067
R39426 S.n1091 S.n1089 0.067
R39427 S.n1214 S.n1212 0.067
R39428 S.n1214 S.n1213 0.067
R39429 S.n1123 S.n1122 0.067
R39430 S.n1123 S.n1121 0.067
R39431 S.n1201 S.n1199 0.067
R39432 S.n1201 S.n1200 0.067
R39433 S.n1188 S.n1186 0.067
R39434 S.n1161 S.n1160 0.067
R39435 S.n1161 S.n1159 0.067
R39436 S.n1188 S.n1187 0.067
R39437 S.n1173 S.n1172 0.067
R39438 S.n1173 S.n1171 0.067
R39439 S.n1425 S.n1423 0.067
R39440 S.n21187 S.n21174 0.067
R39441 S.n21187 S.n21173 0.067
R39442 S.n22789 S.n22788 0.067
R39443 S.n22789 S.n22775 0.067
R39444 S.n973 S.n955 0.064
R39445 S.n20816 S.n20815 0.064
R39446 S.n21190 S.n21187 0.063
R39447 S.n1985 S.n1984 0.063
R39448 S.n1865 S.n1864 0.063
R39449 S.n3146 S.n3145 0.063
R39450 S.n3025 S.n3024 0.063
R39451 S.n4283 S.n4282 0.063
R39452 S.n4151 S.n4150 0.063
R39453 S.n5417 S.n5416 0.063
R39454 S.n5264 S.n5263 0.063
R39455 S.n6528 S.n6527 0.063
R39456 S.n6364 S.n6363 0.063
R39457 S.n7626 S.n7625 0.063
R39458 S.n7441 S.n7440 0.063
R39459 S.n8701 S.n8700 0.063
R39460 S.n8505 S.n8504 0.063
R39461 S.n9764 S.n9763 0.063
R39462 S.n9547 S.n9546 0.063
R39463 S.n10804 S.n10803 0.063
R39464 S.n10576 S.n10575 0.063
R39465 S.n11832 S.n11831 0.063
R39466 S.n11583 S.n11582 0.063
R39467 S.n12837 S.n12836 0.063
R39468 S.n12577 S.n12576 0.063
R39469 S.n13830 S.n13829 0.063
R39470 S.n13549 S.n13548 0.063
R39471 S.n14800 S.n14799 0.063
R39472 S.n14508 S.n14507 0.063
R39473 S.n15758 S.n15757 0.063
R39474 S.n15445 S.n15444 0.063
R39475 S.n16693 S.n16692 0.063
R39476 S.n16369 S.n16368 0.063
R39477 S.n17616 S.n17615 0.063
R39478 S.n17271 S.n17270 0.063
R39479 S.n18516 S.n18515 0.063
R39480 S.n18160 S.n18159 0.063
R39481 S.n19403 S.n19402 0.063
R39482 S.n19026 S.n19025 0.063
R39483 S.n20271 S.n20270 0.063
R39484 S.n19880 S.n19879 0.063
R39485 S.n20491 S.n20490 0.063
R39486 S.n21314 S.n21313 0.063
R39487 S.n2079 S.n2053 0.063
R39488 S.n1799 S.n1784 0.063
R39489 S.n3230 S.n3229 0.063
R39490 S.n2961 S.n2960 0.063
R39491 S.n4367 S.n4366 0.063
R39492 S.n4088 S.n4087 0.063
R39493 S.n5502 S.n5501 0.063
R39494 S.n5200 S.n5199 0.063
R39495 S.n6612 S.n6611 0.063
R39496 S.n6300 S.n6299 0.063
R39497 S.n7710 S.n7709 0.063
R39498 S.n7377 S.n7376 0.063
R39499 S.n8785 S.n8784 0.063
R39500 S.n8441 S.n8440 0.063
R39501 S.n9848 S.n9847 0.063
R39502 S.n9483 S.n9482 0.063
R39503 S.n10888 S.n10887 0.063
R39504 S.n10512 S.n10511 0.063
R39505 S.n11916 S.n11915 0.063
R39506 S.n11519 S.n11518 0.063
R39507 S.n12921 S.n12920 0.063
R39508 S.n12513 S.n12512 0.063
R39509 S.n13914 S.n13913 0.063
R39510 S.n13485 S.n13484 0.063
R39511 S.n14884 S.n14883 0.063
R39512 S.n14444 S.n14443 0.063
R39513 S.n15842 S.n15841 0.063
R39514 S.n15381 S.n15380 0.063
R39515 S.n16777 S.n16776 0.063
R39516 S.n16305 S.n16304 0.063
R39517 S.n17700 S.n17699 0.063
R39518 S.n17207 S.n17206 0.063
R39519 S.n18096 S.n18095 0.063
R39520 S.n18961 S.n18960 0.063
R39521 S.n1337 S.n1336 0.063
R39522 S.n2012 S.n1993 0.063
R39523 S.n3166 S.n3154 0.063
R39524 S.n4303 S.n4291 0.063
R39525 S.n5438 S.n5425 0.063
R39526 S.n6548 S.n6536 0.063
R39527 S.n7646 S.n7634 0.063
R39528 S.n8721 S.n8709 0.063
R39529 S.n9784 S.n9772 0.063
R39530 S.n10824 S.n10812 0.063
R39531 S.n11852 S.n11840 0.063
R39532 S.n12857 S.n12845 0.063
R39533 S.n13850 S.n13838 0.063
R39534 S.n14820 S.n14808 0.063
R39535 S.n15778 S.n15766 0.063
R39536 S.n16713 S.n16701 0.063
R39537 S.n17636 S.n17624 0.063
R39538 S.n18536 S.n18524 0.063
R39539 S.n19423 S.n19411 0.063
R39540 S.n864 S.n848 0.063
R39541 S.n16806 S.n16785 0.063
R39542 S.n15871 S.n15850 0.063
R39543 S.n14913 S.n14892 0.063
R39544 S.n13943 S.n13922 0.063
R39545 S.n12950 S.n12929 0.063
R39546 S.n11945 S.n11924 0.063
R39547 S.n10917 S.n10896 0.063
R39548 S.n9877 S.n9856 0.063
R39549 S.n8814 S.n8793 0.063
R39550 S.n7739 S.n7718 0.063
R39551 S.n6641 S.n6620 0.063
R39552 S.n5531 S.n5510 0.063
R39553 S.n4396 S.n4375 0.063
R39554 S.n3259 S.n3238 0.063
R39555 S.n2107 S.n2088 0.063
R39556 S.n24 S.n8 0.063
R39557 S.n2137 S.n2136 0.063
R39558 S.n1757 S.n1756 0.063
R39559 S.n3290 S.n3289 0.063
R39560 S.n2925 S.n2924 0.063
R39561 S.n4428 S.n4427 0.063
R39562 S.n4052 S.n4051 0.063
R39563 S.n5563 S.n5562 0.063
R39564 S.n5164 S.n5163 0.063
R39565 S.n6673 S.n6672 0.063
R39566 S.n6264 S.n6263 0.063
R39567 S.n7771 S.n7770 0.063
R39568 S.n7341 S.n7340 0.063
R39569 S.n8846 S.n8845 0.063
R39570 S.n8405 S.n8404 0.063
R39571 S.n9909 S.n9908 0.063
R39572 S.n9447 S.n9446 0.063
R39573 S.n10949 S.n10948 0.063
R39574 S.n10476 S.n10475 0.063
R39575 S.n11977 S.n11976 0.063
R39576 S.n11483 S.n11482 0.063
R39577 S.n12982 S.n12981 0.063
R39578 S.n12477 S.n12476 0.063
R39579 S.n13975 S.n13974 0.063
R39580 S.n13449 S.n13448 0.063
R39581 S.n14945 S.n14944 0.063
R39582 S.n14408 S.n14407 0.063
R39583 S.n15903 S.n15902 0.063
R39584 S.n15345 S.n15344 0.063
R39585 S.n16269 S.n16268 0.063
R39586 S.n17169 S.n17168 0.063
R39587 S.n14974 S.n14953 0.063
R39588 S.n14004 S.n13983 0.063
R39589 S.n13011 S.n12990 0.063
R39590 S.n12006 S.n11985 0.063
R39591 S.n10978 S.n10957 0.063
R39592 S.n9938 S.n9917 0.063
R39593 S.n8875 S.n8854 0.063
R39594 S.n7800 S.n7779 0.063
R39595 S.n6702 S.n6681 0.063
R39596 S.n5592 S.n5571 0.063
R39597 S.n4457 S.n4436 0.063
R39598 S.n3319 S.n3298 0.063
R39599 S.n2166 S.n2146 0.063
R39600 S.n71 S.n55 0.063
R39601 S.n2196 S.n2195 0.063
R39602 S.n1720 S.n1719 0.063
R39603 S.n3350 S.n3349 0.063
R39604 S.n2889 S.n2888 0.063
R39605 S.n4489 S.n4488 0.063
R39606 S.n4016 S.n4015 0.063
R39607 S.n5624 S.n5623 0.063
R39608 S.n5128 S.n5127 0.063
R39609 S.n6734 S.n6733 0.063
R39610 S.n6228 S.n6227 0.063
R39611 S.n7832 S.n7831 0.063
R39612 S.n7305 S.n7304 0.063
R39613 S.n8907 S.n8906 0.063
R39614 S.n8369 S.n8368 0.063
R39615 S.n9970 S.n9969 0.063
R39616 S.n9411 S.n9410 0.063
R39617 S.n11010 S.n11009 0.063
R39618 S.n10440 S.n10439 0.063
R39619 S.n12038 S.n12037 0.063
R39620 S.n11447 S.n11446 0.063
R39621 S.n13043 S.n13042 0.063
R39622 S.n12441 S.n12440 0.063
R39623 S.n14036 S.n14035 0.063
R39624 S.n13413 S.n13412 0.063
R39625 S.n14372 S.n14371 0.063
R39626 S.n15307 S.n15306 0.063
R39627 S.n13072 S.n13051 0.063
R39628 S.n12067 S.n12046 0.063
R39629 S.n11039 S.n11018 0.063
R39630 S.n9999 S.n9978 0.063
R39631 S.n8936 S.n8915 0.063
R39632 S.n7861 S.n7840 0.063
R39633 S.n6763 S.n6742 0.063
R39634 S.n5653 S.n5632 0.063
R39635 S.n4518 S.n4497 0.063
R39636 S.n3379 S.n3358 0.063
R39637 S.n2225 S.n2205 0.063
R39638 S.n103 S.n85 0.063
R39639 S.n2255 S.n2254 0.063
R39640 S.n1683 S.n1682 0.063
R39641 S.n3410 S.n3409 0.063
R39642 S.n2853 S.n2852 0.063
R39643 S.n4550 S.n4549 0.063
R39644 S.n3980 S.n3979 0.063
R39645 S.n5685 S.n5684 0.063
R39646 S.n5092 S.n5091 0.063
R39647 S.n6795 S.n6794 0.063
R39648 S.n6192 S.n6191 0.063
R39649 S.n7893 S.n7892 0.063
R39650 S.n7269 S.n7268 0.063
R39651 S.n8968 S.n8967 0.063
R39652 S.n8333 S.n8332 0.063
R39653 S.n10031 S.n10030 0.063
R39654 S.n9375 S.n9374 0.063
R39655 S.n11071 S.n11070 0.063
R39656 S.n10404 S.n10403 0.063
R39657 S.n12099 S.n12098 0.063
R39658 S.n11411 S.n11410 0.063
R39659 S.n12405 S.n12404 0.063
R39660 S.n13375 S.n13374 0.063
R39661 S.n11100 S.n11079 0.063
R39662 S.n10060 S.n10039 0.063
R39663 S.n8997 S.n8976 0.063
R39664 S.n7922 S.n7901 0.063
R39665 S.n6824 S.n6803 0.063
R39666 S.n5714 S.n5693 0.063
R39667 S.n4579 S.n4558 0.063
R39668 S.n3439 S.n3418 0.063
R39669 S.n2284 S.n2264 0.063
R39670 S.n990 S.n119 0.063
R39671 S.n2314 S.n2313 0.063
R39672 S.n1646 S.n1645 0.063
R39673 S.n3470 S.n3469 0.063
R39674 S.n2817 S.n2816 0.063
R39675 S.n4611 S.n4610 0.063
R39676 S.n3944 S.n3943 0.063
R39677 S.n5746 S.n5745 0.063
R39678 S.n5056 S.n5055 0.063
R39679 S.n6856 S.n6855 0.063
R39680 S.n6156 S.n6155 0.063
R39681 S.n7954 S.n7953 0.063
R39682 S.n7233 S.n7232 0.063
R39683 S.n9029 S.n9028 0.063
R39684 S.n8297 S.n8296 0.063
R39685 S.n10092 S.n10091 0.063
R39686 S.n9339 S.n9338 0.063
R39687 S.n10368 S.n10367 0.063
R39688 S.n11373 S.n11372 0.063
R39689 S.n9058 S.n9037 0.063
R39690 S.n7983 S.n7962 0.063
R39691 S.n6885 S.n6864 0.063
R39692 S.n5775 S.n5754 0.063
R39693 S.n4640 S.n4619 0.063
R39694 S.n3499 S.n3478 0.063
R39695 S.n2343 S.n2323 0.063
R39696 S.n1022 S.n1006 0.063
R39697 S.n2373 S.n2372 0.063
R39698 S.n1609 S.n1608 0.063
R39699 S.n3530 S.n3529 0.063
R39700 S.n2781 S.n2780 0.063
R39701 S.n4672 S.n4671 0.063
R39702 S.n3908 S.n3907 0.063
R39703 S.n5807 S.n5806 0.063
R39704 S.n5020 S.n5019 0.063
R39705 S.n6917 S.n6916 0.063
R39706 S.n6120 S.n6119 0.063
R39707 S.n8015 S.n8014 0.063
R39708 S.n7197 S.n7196 0.063
R39709 S.n8261 S.n8260 0.063
R39710 S.n9301 S.n9300 0.063
R39711 S.n6946 S.n6925 0.063
R39712 S.n5836 S.n5815 0.063
R39713 S.n4701 S.n4680 0.063
R39714 S.n3559 S.n3538 0.063
R39715 S.n2402 S.n2382 0.063
R39716 S.n1054 S.n1036 0.063
R39717 S.n2432 S.n2431 0.063
R39718 S.n1572 S.n1571 0.063
R39719 S.n3590 S.n3589 0.063
R39720 S.n2745 S.n2744 0.063
R39721 S.n4733 S.n4732 0.063
R39722 S.n3872 S.n3871 0.063
R39723 S.n5868 S.n5867 0.063
R39724 S.n4984 S.n4983 0.063
R39725 S.n6084 S.n6083 0.063
R39726 S.n7159 S.n7158 0.063
R39727 S.n4762 S.n4741 0.063
R39728 S.n3619 S.n3598 0.063
R39729 S.n2461 S.n2441 0.063
R39730 S.n1086 S.n1070 0.063
R39731 S.n2491 S.n2490 0.063
R39732 S.n1535 S.n1534 0.063
R39733 S.n3650 S.n3649 0.063
R39734 S.n2709 S.n2708 0.063
R39735 S.n3836 S.n3835 0.063
R39736 S.n4946 S.n4945 0.063
R39737 S.n2520 S.n2500 0.063
R39738 S.n1118 S.n1102 0.063
R39739 S.n1498 S.n1497 0.063
R39740 S.n2671 S.n2670 0.063
R39741 S.n1156 S.n1132 0.063
R39742 S.n942 S.n941 0.063
R39743 S.n22691 S.n22690 0.062
R39744 S.n22693 S.n22692 0.062
R39745 S.n22704 S.n22701 0.062
R39746 S.n22703 S.n22702 0.062
R39747 S.n21252 S.n21249 0.062
R39748 S.n21251 S.n21250 0.062
R39749 S.n1426 S.n1425 0.062
R39750 S.n1292 S.n1291 0.062
R39751 S.n1280 S.n1279 0.062
R39752 S.n1267 S.n1266 0.062
R39753 S.n1254 S.n1253 0.062
R39754 S.n1241 S.n1240 0.062
R39755 S.n1228 S.n1227 0.062
R39756 S.n1215 S.n1214 0.062
R39757 S.n1202 S.n1201 0.062
R39758 S.n1189 S.n1188 0.062
R39759 S.n1353 S.n1342 0.061
R39760 S.n46 S.n45 0.06
R39761 S.n77 S.n76 0.06
R39762 S.n109 S.n108 0.06
R39763 S.n996 S.n995 0.06
R39764 S.n1028 S.n1027 0.06
R39765 S.n1060 S.n1059 0.06
R39766 S.n1092 S.n1091 0.06
R39767 S.n1124 S.n1123 0.06
R39768 S.n1162 S.n1161 0.06
R39769 S.n1174 S.n1173 0.06
R39770 S.n22737 S.n22736 0.059
R39771 S.n21226 S.n21225 0.059
R39772 S.n20350 S.n20349 0.059
R39773 S.n20279 S.n20278 0.059
R39774 S.n18610 S.n18609 0.059
R39775 S.n17710 S.n17709 0.059
R39776 S.n16848 S.n16847 0.059
R39777 S.n15913 S.n15912 0.059
R39778 S.n15016 S.n15015 0.059
R39779 S.n14046 S.n14045 0.059
R39780 S.n13114 S.n13113 0.059
R39781 S.n12109 S.n12108 0.059
R39782 S.n11142 S.n11141 0.059
R39783 S.n10102 S.n10101 0.059
R39784 S.n9100 S.n9099 0.059
R39785 S.n8025 S.n8024 0.059
R39786 S.n6988 S.n6987 0.059
R39787 S.n5878 S.n5877 0.059
R39788 S.n4804 S.n4803 0.059
R39789 S.n3660 S.n3659 0.059
R39790 S.n2560 S.n2559 0.059
R39791 S.n3216 S.n3206 0.059
R39792 S.n1305 S.n1304 0.059
R39793 S.n3745 S.n3744 0.058
R39794 S.n2614 S.n2613 0.058
R39795 S.n973 S.n972 0.058
R39796 S.n22790 S.n22789 0.058
R39797 S.n19520 S.n19519 0.058
R39798 S.n18663 S.n18662 0.058
R39799 S.n17795 S.n17794 0.058
R39800 S.n16901 S.n16900 0.058
R39801 S.n15998 S.n15997 0.058
R39802 S.n15069 S.n15068 0.058
R39803 S.n14131 S.n14130 0.058
R39804 S.n13167 S.n13166 0.058
R39805 S.n12194 S.n12193 0.058
R39806 S.n11195 S.n11194 0.058
R39807 S.n10187 S.n10186 0.058
R39808 S.n9153 S.n9152 0.058
R39809 S.n8110 S.n8109 0.058
R39810 S.n7041 S.n7040 0.058
R39811 S.n5963 S.n5962 0.058
R39812 S.n4858 S.n4857 0.058
R39813 S.n2 S.n1 0.056
R39814 S.n1371 S.n1370 0.056
R39815 S.n49 S.n48 0.056
R39816 S.n80 S.n79 0.056
R39817 S.n112 S.n111 0.056
R39818 S.n999 S.n998 0.056
R39819 S.n1031 S.n1030 0.056
R39820 S.n1063 S.n1062 0.056
R39821 S.n1095 S.n1094 0.056
R39822 S.n1127 S.n1126 0.056
R39823 S.n1165 S.n1164 0.056
R39824 S.n1184 S.n1175 0.055
R39825 S.n21144 S.n21143 0.055
R39826 S.n20343 S.n20342 0.055
R39827 S.n19503 S.n19502 0.055
R39828 S.n18646 S.n18645 0.055
R39829 S.n17778 S.n17777 0.055
R39830 S.n16884 S.n16883 0.055
R39831 S.n15981 S.n15980 0.055
R39832 S.n15052 S.n15051 0.055
R39833 S.n14114 S.n14113 0.055
R39834 S.n13150 S.n13149 0.055
R39835 S.n12177 S.n12176 0.055
R39836 S.n11178 S.n11177 0.055
R39837 S.n10170 S.n10169 0.055
R39838 S.n9136 S.n9135 0.055
R39839 S.n8093 S.n8092 0.055
R39840 S.n7024 S.n7023 0.055
R39841 S.n5946 S.n5945 0.055
R39842 S.n4840 S.n4839 0.055
R39843 S.n3727 S.n3726 0.055
R39844 S.n2596 S.n2595 0.055
R39845 S.n979 S.n978 0.055
R39846 S.n21973 S.n21972 0.055
R39847 S.n22774 S.n21982 0.054
R39848 S.n22289 S.n22270 0.054
R39849 S.n18060 S.n18046 0.054
R39850 S.n18944 S.n18929 0.054
R39851 S.n19815 S.n19801 0.054
R39852 S.n20452 S.n20435 0.054
R39853 S.n21297 S.n21281 0.054
R39854 S.n16233 S.n16219 0.054
R39855 S.n17152 S.n17137 0.054
R39856 S.n14336 S.n14322 0.054
R39857 S.n15290 S.n15275 0.054
R39858 S.n12369 S.n12355 0.054
R39859 S.n13358 S.n13343 0.054
R39860 S.n10332 S.n10318 0.054
R39861 S.n11356 S.n11341 0.054
R39862 S.n8225 S.n8211 0.054
R39863 S.n9284 S.n9269 0.054
R39864 S.n6048 S.n6034 0.054
R39865 S.n7142 S.n7127 0.054
R39866 S.n3800 S.n3786 0.054
R39867 S.n4929 S.n4914 0.054
R39868 S.n1461 S.n1446 0.054
R39869 S.n2654 S.n2639 0.054
R39870 S.n433 S.n417 0.054
R39871 S.n1814 S.n1813 0.054
R39872 S.n2977 S.n2976 0.054
R39873 S.n4104 S.n4103 0.054
R39874 S.n5216 S.n5215 0.054
R39875 S.n6316 S.n6315 0.054
R39876 S.n7393 S.n7392 0.054
R39877 S.n8457 S.n8456 0.054
R39878 S.n9499 S.n9498 0.054
R39879 S.n10528 S.n10527 0.054
R39880 S.n11535 S.n11534 0.054
R39881 S.n12529 S.n12528 0.054
R39882 S.n13501 S.n13500 0.054
R39883 S.n14460 S.n14459 0.054
R39884 S.n15397 S.n15396 0.054
R39885 S.n16321 S.n16320 0.054
R39886 S.n17223 S.n17222 0.054
R39887 S.n18112 S.n18111 0.054
R39888 S.n18977 S.n18976 0.054
R39889 S.n19829 S.n19828 0.054
R39890 S.n762 S.n761 0.054
R39891 S.n22804 S.n22802 0.054
R39892 S.n45 S.n44 0.054
R39893 S.n20189 S.n20188 0.054
R39894 S.n21139 S.n21138 0.054
R39895 S.n22646 S.n22645 0.054
R39896 S.n22013 S.n22012 0.054
R39897 S.n21623 S.n21622 0.054
R39898 S.n21948 S.n21947 0.054
R39899 S.n20800 S.n20799 0.054
R39900 S.n22662 S.n22661 0.054
R39901 S.n21998 S.n21997 0.054
R39902 S.n21644 S.n21643 0.054
R39903 S.n21968 S.n21967 0.054
R39904 S.n20824 S.n20823 0.054
R39905 S.n19319 S.n19318 0.054
R39906 S.n19536 S.n19535 0.054
R39907 S.n22630 S.n22629 0.054
R39908 S.n22028 S.n22027 0.054
R39909 S.n21607 S.n21606 0.054
R39910 S.n21933 S.n21932 0.054
R39911 S.n20784 S.n20783 0.054
R39912 S.n21123 S.n21122 0.054
R39913 S.n20173 S.n20172 0.054
R39914 S.n18437 S.n18436 0.054
R39915 S.n18679 S.n18678 0.054
R39916 S.n22614 S.n22613 0.054
R39917 S.n22043 S.n22042 0.054
R39918 S.n21591 S.n21590 0.054
R39919 S.n21918 S.n21917 0.054
R39920 S.n20768 S.n20767 0.054
R39921 S.n21108 S.n21107 0.054
R39922 S.n20157 S.n20156 0.054
R39923 S.n19551 S.n19550 0.054
R39924 S.n19303 S.n19302 0.054
R39925 S.n17532 S.n17531 0.054
R39926 S.n17811 S.n17810 0.054
R39927 S.n22598 S.n22597 0.054
R39928 S.n22058 S.n22057 0.054
R39929 S.n21575 S.n21574 0.054
R39930 S.n21903 S.n21902 0.054
R39931 S.n20752 S.n20751 0.054
R39932 S.n21093 S.n21092 0.054
R39933 S.n20141 S.n20140 0.054
R39934 S.n19566 S.n19565 0.054
R39935 S.n19287 S.n19286 0.054
R39936 S.n18694 S.n18693 0.054
R39937 S.n18421 S.n18420 0.054
R39938 S.n16614 S.n16613 0.054
R39939 S.n16917 S.n16916 0.054
R39940 S.n22582 S.n22581 0.054
R39941 S.n22073 S.n22072 0.054
R39942 S.n21559 S.n21558 0.054
R39943 S.n21888 S.n21887 0.054
R39944 S.n20736 S.n20735 0.054
R39945 S.n21078 S.n21077 0.054
R39946 S.n20125 S.n20124 0.054
R39947 S.n19581 S.n19580 0.054
R39948 S.n19271 S.n19270 0.054
R39949 S.n18709 S.n18708 0.054
R39950 S.n18405 S.n18404 0.054
R39951 S.n17826 S.n17825 0.054
R39952 S.n17516 S.n17515 0.054
R39953 S.n15674 S.n15673 0.054
R39954 S.n16014 S.n16013 0.054
R39955 S.n22566 S.n22565 0.054
R39956 S.n22088 S.n22087 0.054
R39957 S.n21543 S.n21542 0.054
R39958 S.n21873 S.n21872 0.054
R39959 S.n20720 S.n20719 0.054
R39960 S.n21063 S.n21062 0.054
R39961 S.n20109 S.n20108 0.054
R39962 S.n19596 S.n19595 0.054
R39963 S.n19255 S.n19254 0.054
R39964 S.n18724 S.n18723 0.054
R39965 S.n18389 S.n18388 0.054
R39966 S.n17841 S.n17840 0.054
R39967 S.n17500 S.n17499 0.054
R39968 S.n16932 S.n16931 0.054
R39969 S.n16598 S.n16597 0.054
R39970 S.n14721 S.n14720 0.054
R39971 S.n15085 S.n15084 0.054
R39972 S.n22550 S.n22549 0.054
R39973 S.n22103 S.n22102 0.054
R39974 S.n21527 S.n21526 0.054
R39975 S.n21858 S.n21857 0.054
R39976 S.n20704 S.n20703 0.054
R39977 S.n21048 S.n21047 0.054
R39978 S.n20093 S.n20092 0.054
R39979 S.n19611 S.n19610 0.054
R39980 S.n19239 S.n19238 0.054
R39981 S.n18739 S.n18738 0.054
R39982 S.n18373 S.n18372 0.054
R39983 S.n17856 S.n17855 0.054
R39984 S.n17484 S.n17483 0.054
R39985 S.n16947 S.n16946 0.054
R39986 S.n16582 S.n16581 0.054
R39987 S.n16029 S.n16028 0.054
R39988 S.n15658 S.n15657 0.054
R39989 S.n13746 S.n13745 0.054
R39990 S.n14147 S.n14146 0.054
R39991 S.n22534 S.n22533 0.054
R39992 S.n22118 S.n22117 0.054
R39993 S.n21511 S.n21510 0.054
R39994 S.n21843 S.n21842 0.054
R39995 S.n20688 S.n20687 0.054
R39996 S.n21033 S.n21032 0.054
R39997 S.n20077 S.n20076 0.054
R39998 S.n19626 S.n19625 0.054
R39999 S.n19223 S.n19222 0.054
R40000 S.n18754 S.n18753 0.054
R40001 S.n18357 S.n18356 0.054
R40002 S.n17871 S.n17870 0.054
R40003 S.n17468 S.n17467 0.054
R40004 S.n16962 S.n16961 0.054
R40005 S.n16566 S.n16565 0.054
R40006 S.n16044 S.n16043 0.054
R40007 S.n15642 S.n15641 0.054
R40008 S.n15100 S.n15099 0.054
R40009 S.n14705 S.n14704 0.054
R40010 S.n12758 S.n12757 0.054
R40011 S.n13183 S.n13182 0.054
R40012 S.n22518 S.n22517 0.054
R40013 S.n22133 S.n22132 0.054
R40014 S.n21495 S.n21494 0.054
R40015 S.n21828 S.n21827 0.054
R40016 S.n20672 S.n20671 0.054
R40017 S.n21018 S.n21017 0.054
R40018 S.n20061 S.n20060 0.054
R40019 S.n19641 S.n19640 0.054
R40020 S.n19207 S.n19206 0.054
R40021 S.n18769 S.n18768 0.054
R40022 S.n18341 S.n18340 0.054
R40023 S.n17886 S.n17885 0.054
R40024 S.n17452 S.n17451 0.054
R40025 S.n16977 S.n16976 0.054
R40026 S.n16550 S.n16549 0.054
R40027 S.n16059 S.n16058 0.054
R40028 S.n15626 S.n15625 0.054
R40029 S.n15115 S.n15114 0.054
R40030 S.n14689 S.n14688 0.054
R40031 S.n14162 S.n14161 0.054
R40032 S.n13730 S.n13729 0.054
R40033 S.n11748 S.n11747 0.054
R40034 S.n12210 S.n12209 0.054
R40035 S.n22502 S.n22501 0.054
R40036 S.n22148 S.n22147 0.054
R40037 S.n21479 S.n21478 0.054
R40038 S.n21813 S.n21812 0.054
R40039 S.n20656 S.n20655 0.054
R40040 S.n21003 S.n21002 0.054
R40041 S.n20045 S.n20044 0.054
R40042 S.n19656 S.n19655 0.054
R40043 S.n19191 S.n19190 0.054
R40044 S.n18784 S.n18783 0.054
R40045 S.n18325 S.n18324 0.054
R40046 S.n17901 S.n17900 0.054
R40047 S.n17436 S.n17435 0.054
R40048 S.n16992 S.n16991 0.054
R40049 S.n16534 S.n16533 0.054
R40050 S.n16074 S.n16073 0.054
R40051 S.n15610 S.n15609 0.054
R40052 S.n15130 S.n15129 0.054
R40053 S.n14673 S.n14672 0.054
R40054 S.n14177 S.n14176 0.054
R40055 S.n13714 S.n13713 0.054
R40056 S.n13198 S.n13197 0.054
R40057 S.n12742 S.n12741 0.054
R40058 S.n10725 S.n10724 0.054
R40059 S.n11211 S.n11210 0.054
R40060 S.n22486 S.n22485 0.054
R40061 S.n22163 S.n22162 0.054
R40062 S.n21463 S.n21462 0.054
R40063 S.n21798 S.n21797 0.054
R40064 S.n20640 S.n20639 0.054
R40065 S.n20988 S.n20987 0.054
R40066 S.n20029 S.n20028 0.054
R40067 S.n19671 S.n19670 0.054
R40068 S.n19175 S.n19174 0.054
R40069 S.n18799 S.n18798 0.054
R40070 S.n18309 S.n18308 0.054
R40071 S.n17916 S.n17915 0.054
R40072 S.n17420 S.n17419 0.054
R40073 S.n17007 S.n17006 0.054
R40074 S.n16518 S.n16517 0.054
R40075 S.n16089 S.n16088 0.054
R40076 S.n15594 S.n15593 0.054
R40077 S.n15145 S.n15144 0.054
R40078 S.n14657 S.n14656 0.054
R40079 S.n14192 S.n14191 0.054
R40080 S.n13698 S.n13697 0.054
R40081 S.n13213 S.n13212 0.054
R40082 S.n12726 S.n12725 0.054
R40083 S.n12225 S.n12224 0.054
R40084 S.n11732 S.n11731 0.054
R40085 S.n9680 S.n9679 0.054
R40086 S.n10203 S.n10202 0.054
R40087 S.n22470 S.n22469 0.054
R40088 S.n22178 S.n22177 0.054
R40089 S.n21447 S.n21446 0.054
R40090 S.n21783 S.n21782 0.054
R40091 S.n20624 S.n20623 0.054
R40092 S.n20973 S.n20972 0.054
R40093 S.n20013 S.n20012 0.054
R40094 S.n19686 S.n19685 0.054
R40095 S.n19159 S.n19158 0.054
R40096 S.n18814 S.n18813 0.054
R40097 S.n18293 S.n18292 0.054
R40098 S.n17931 S.n17930 0.054
R40099 S.n17404 S.n17403 0.054
R40100 S.n17022 S.n17021 0.054
R40101 S.n16502 S.n16501 0.054
R40102 S.n16104 S.n16103 0.054
R40103 S.n15578 S.n15577 0.054
R40104 S.n15160 S.n15159 0.054
R40105 S.n14641 S.n14640 0.054
R40106 S.n14207 S.n14206 0.054
R40107 S.n13682 S.n13681 0.054
R40108 S.n13228 S.n13227 0.054
R40109 S.n12710 S.n12709 0.054
R40110 S.n12240 S.n12239 0.054
R40111 S.n11716 S.n11715 0.054
R40112 S.n11226 S.n11225 0.054
R40113 S.n10709 S.n10708 0.054
R40114 S.n8622 S.n8621 0.054
R40115 S.n9169 S.n9168 0.054
R40116 S.n22454 S.n22453 0.054
R40117 S.n22193 S.n22192 0.054
R40118 S.n21431 S.n21430 0.054
R40119 S.n21768 S.n21767 0.054
R40120 S.n20608 S.n20607 0.054
R40121 S.n20958 S.n20957 0.054
R40122 S.n19997 S.n19996 0.054
R40123 S.n19701 S.n19700 0.054
R40124 S.n19143 S.n19142 0.054
R40125 S.n18829 S.n18828 0.054
R40126 S.n18277 S.n18276 0.054
R40127 S.n17946 S.n17945 0.054
R40128 S.n17388 S.n17387 0.054
R40129 S.n17037 S.n17036 0.054
R40130 S.n16486 S.n16485 0.054
R40131 S.n16119 S.n16118 0.054
R40132 S.n15562 S.n15561 0.054
R40133 S.n15175 S.n15174 0.054
R40134 S.n14625 S.n14624 0.054
R40135 S.n14222 S.n14221 0.054
R40136 S.n13666 S.n13665 0.054
R40137 S.n13243 S.n13242 0.054
R40138 S.n12694 S.n12693 0.054
R40139 S.n12255 S.n12254 0.054
R40140 S.n11700 S.n11699 0.054
R40141 S.n11241 S.n11240 0.054
R40142 S.n10693 S.n10692 0.054
R40143 S.n10218 S.n10217 0.054
R40144 S.n9664 S.n9663 0.054
R40145 S.n7542 S.n7541 0.054
R40146 S.n8126 S.n8125 0.054
R40147 S.n22438 S.n22437 0.054
R40148 S.n22208 S.n22207 0.054
R40149 S.n21415 S.n21414 0.054
R40150 S.n21753 S.n21752 0.054
R40151 S.n20592 S.n20591 0.054
R40152 S.n20943 S.n20942 0.054
R40153 S.n19981 S.n19980 0.054
R40154 S.n19716 S.n19715 0.054
R40155 S.n19127 S.n19126 0.054
R40156 S.n18844 S.n18843 0.054
R40157 S.n18261 S.n18260 0.054
R40158 S.n17961 S.n17960 0.054
R40159 S.n17372 S.n17371 0.054
R40160 S.n17052 S.n17051 0.054
R40161 S.n16470 S.n16469 0.054
R40162 S.n16134 S.n16133 0.054
R40163 S.n15546 S.n15545 0.054
R40164 S.n15190 S.n15189 0.054
R40165 S.n14609 S.n14608 0.054
R40166 S.n14237 S.n14236 0.054
R40167 S.n13650 S.n13649 0.054
R40168 S.n13258 S.n13257 0.054
R40169 S.n12678 S.n12677 0.054
R40170 S.n12270 S.n12269 0.054
R40171 S.n11684 S.n11683 0.054
R40172 S.n11256 S.n11255 0.054
R40173 S.n10677 S.n10676 0.054
R40174 S.n10233 S.n10232 0.054
R40175 S.n9648 S.n9647 0.054
R40176 S.n9184 S.n9183 0.054
R40177 S.n8606 S.n8605 0.054
R40178 S.n6449 S.n6448 0.054
R40179 S.n7057 S.n7056 0.054
R40180 S.n22422 S.n22421 0.054
R40181 S.n22223 S.n22222 0.054
R40182 S.n21399 S.n21398 0.054
R40183 S.n21738 S.n21737 0.054
R40184 S.n20576 S.n20575 0.054
R40185 S.n20928 S.n20927 0.054
R40186 S.n19965 S.n19964 0.054
R40187 S.n19731 S.n19730 0.054
R40188 S.n19111 S.n19110 0.054
R40189 S.n18859 S.n18858 0.054
R40190 S.n18245 S.n18244 0.054
R40191 S.n17976 S.n17975 0.054
R40192 S.n17356 S.n17355 0.054
R40193 S.n17067 S.n17066 0.054
R40194 S.n16454 S.n16453 0.054
R40195 S.n16149 S.n16148 0.054
R40196 S.n15530 S.n15529 0.054
R40197 S.n15205 S.n15204 0.054
R40198 S.n14593 S.n14592 0.054
R40199 S.n14252 S.n14251 0.054
R40200 S.n13634 S.n13633 0.054
R40201 S.n13273 S.n13272 0.054
R40202 S.n12662 S.n12661 0.054
R40203 S.n12285 S.n12284 0.054
R40204 S.n11668 S.n11667 0.054
R40205 S.n11271 S.n11270 0.054
R40206 S.n10661 S.n10660 0.054
R40207 S.n10248 S.n10247 0.054
R40208 S.n9632 S.n9631 0.054
R40209 S.n9199 S.n9198 0.054
R40210 S.n8590 S.n8589 0.054
R40211 S.n8141 S.n8140 0.054
R40212 S.n7526 S.n7525 0.054
R40213 S.n5333 S.n5332 0.054
R40214 S.n5979 S.n5978 0.054
R40215 S.n22406 S.n22405 0.054
R40216 S.n22238 S.n22237 0.054
R40217 S.n21383 S.n21382 0.054
R40218 S.n21723 S.n21722 0.054
R40219 S.n20560 S.n20559 0.054
R40220 S.n20913 S.n20912 0.054
R40221 S.n19949 S.n19948 0.054
R40222 S.n19746 S.n19745 0.054
R40223 S.n19095 S.n19094 0.054
R40224 S.n18874 S.n18873 0.054
R40225 S.n18229 S.n18228 0.054
R40226 S.n17991 S.n17990 0.054
R40227 S.n17340 S.n17339 0.054
R40228 S.n17082 S.n17081 0.054
R40229 S.n16438 S.n16437 0.054
R40230 S.n16164 S.n16163 0.054
R40231 S.n15514 S.n15513 0.054
R40232 S.n15220 S.n15219 0.054
R40233 S.n14577 S.n14576 0.054
R40234 S.n14267 S.n14266 0.054
R40235 S.n13618 S.n13617 0.054
R40236 S.n13288 S.n13287 0.054
R40237 S.n12646 S.n12645 0.054
R40238 S.n12300 S.n12299 0.054
R40239 S.n11652 S.n11651 0.054
R40240 S.n11286 S.n11285 0.054
R40241 S.n10645 S.n10644 0.054
R40242 S.n10263 S.n10262 0.054
R40243 S.n9616 S.n9615 0.054
R40244 S.n9214 S.n9213 0.054
R40245 S.n8574 S.n8573 0.054
R40246 S.n8156 S.n8155 0.054
R40247 S.n7510 S.n7509 0.054
R40248 S.n7072 S.n7071 0.054
R40249 S.n6433 S.n6432 0.054
R40250 S.n4204 S.n4203 0.054
R40251 S.n4874 S.n4873 0.054
R40252 S.n22390 S.n22389 0.054
R40253 S.n22253 S.n22252 0.054
R40254 S.n21367 S.n21366 0.054
R40255 S.n21708 S.n21707 0.054
R40256 S.n20544 S.n20543 0.054
R40257 S.n20898 S.n20897 0.054
R40258 S.n19933 S.n19932 0.054
R40259 S.n19761 S.n19760 0.054
R40260 S.n19079 S.n19078 0.054
R40261 S.n18889 S.n18888 0.054
R40262 S.n18213 S.n18212 0.054
R40263 S.n18006 S.n18005 0.054
R40264 S.n17324 S.n17323 0.054
R40265 S.n17097 S.n17096 0.054
R40266 S.n16422 S.n16421 0.054
R40267 S.n16179 S.n16178 0.054
R40268 S.n15498 S.n15497 0.054
R40269 S.n15235 S.n15234 0.054
R40270 S.n14561 S.n14560 0.054
R40271 S.n14282 S.n14281 0.054
R40272 S.n13602 S.n13601 0.054
R40273 S.n13303 S.n13302 0.054
R40274 S.n12630 S.n12629 0.054
R40275 S.n12315 S.n12314 0.054
R40276 S.n11636 S.n11635 0.054
R40277 S.n11301 S.n11300 0.054
R40278 S.n10629 S.n10628 0.054
R40279 S.n10278 S.n10277 0.054
R40280 S.n9600 S.n9599 0.054
R40281 S.n9220 S.n9219 0.054
R40282 S.n8558 S.n8557 0.054
R40283 S.n8171 S.n8170 0.054
R40284 S.n7494 S.n7493 0.054
R40285 S.n7087 S.n7086 0.054
R40286 S.n6417 S.n6416 0.054
R40287 S.n5994 S.n5993 0.054
R40288 S.n5317 S.n5316 0.054
R40289 S.n3063 S.n3062 0.054
R40290 S.n3762 S.n3761 0.054
R40291 S.n22665 S.n22664 0.054
R40292 S.n22678 S.n22677 0.054
R40293 S.n21678 S.n21677 0.054
R40294 S.n21693 S.n21692 0.054
R40295 S.n20528 S.n20527 0.054
R40296 S.n20883 S.n20882 0.054
R40297 S.n19917 S.n19916 0.054
R40298 S.n19777 S.n19776 0.054
R40299 S.n19063 S.n19062 0.054
R40300 S.n18905 S.n18904 0.054
R40301 S.n18197 S.n18196 0.054
R40302 S.n18022 S.n18021 0.054
R40303 S.n17308 S.n17307 0.054
R40304 S.n17113 S.n17112 0.054
R40305 S.n16406 S.n16405 0.054
R40306 S.n16195 S.n16194 0.054
R40307 S.n15482 S.n15481 0.054
R40308 S.n15251 S.n15250 0.054
R40309 S.n14545 S.n14544 0.054
R40310 S.n14298 S.n14297 0.054
R40311 S.n13586 S.n13585 0.054
R40312 S.n13319 S.n13318 0.054
R40313 S.n12614 S.n12613 0.054
R40314 S.n12331 S.n12330 0.054
R40315 S.n11620 S.n11619 0.054
R40316 S.n11317 S.n11316 0.054
R40317 S.n10613 S.n10612 0.054
R40318 S.n10294 S.n10293 0.054
R40319 S.n9584 S.n9583 0.054
R40320 S.n9245 S.n9244 0.054
R40321 S.n8542 S.n8541 0.054
R40322 S.n8187 S.n8186 0.054
R40323 S.n7478 S.n7477 0.054
R40324 S.n7103 S.n7102 0.054
R40325 S.n6401 S.n6400 0.054
R40326 S.n6010 S.n6009 0.054
R40327 S.n5301 S.n5300 0.054
R40328 S.n4890 S.n4889 0.054
R40329 S.n4188 S.n4187 0.054
R40330 S.n1894 S.n1893 0.054
R40331 S.n2631 S.n2630 0.054
R40332 S.n22374 S.n22373 0.054
R40333 S.n22697 S.n22696 0.054
R40334 S.n21647 S.n21646 0.054
R40335 S.n21662 S.n21661 0.054
R40336 S.n20513 S.n20512 0.054
R40337 S.n20867 S.n20866 0.054
R40338 S.n19902 S.n19901 0.054
R40339 S.n19793 S.n19792 0.054
R40340 S.n19048 S.n19047 0.054
R40341 S.n18921 S.n18920 0.054
R40342 S.n18182 S.n18181 0.054
R40343 S.n18038 S.n18037 0.054
R40344 S.n17293 S.n17292 0.054
R40345 S.n17129 S.n17128 0.054
R40346 S.n16391 S.n16390 0.054
R40347 S.n16211 S.n16210 0.054
R40348 S.n15467 S.n15466 0.054
R40349 S.n15267 S.n15266 0.054
R40350 S.n14530 S.n14529 0.054
R40351 S.n14314 S.n14313 0.054
R40352 S.n13571 S.n13570 0.054
R40353 S.n13335 S.n13334 0.054
R40354 S.n12599 S.n12598 0.054
R40355 S.n12347 S.n12346 0.054
R40356 S.n11605 S.n11604 0.054
R40357 S.n11333 S.n11332 0.054
R40358 S.n10598 S.n10597 0.054
R40359 S.n10310 S.n10309 0.054
R40360 S.n9569 S.n9568 0.054
R40361 S.n9261 S.n9260 0.054
R40362 S.n8527 S.n8526 0.054
R40363 S.n8203 S.n8202 0.054
R40364 S.n7463 S.n7462 0.054
R40365 S.n7119 S.n7118 0.054
R40366 S.n6386 S.n6385 0.054
R40367 S.n6026 S.n6025 0.054
R40368 S.n5286 S.n5285 0.054
R40369 S.n4906 S.n4905 0.054
R40370 S.n4173 S.n4172 0.054
R40371 S.n3778 S.n3777 0.054
R40372 S.n3047 S.n3046 0.054
R40373 S.n917 S.n916 0.054
R40374 S.n1991 S.n1990 0.054
R40375 S.n22744 S.n22743 0.054
R40376 S.n21317 S.n21316 0.054
R40377 S.n21220 S.n21219 0.054
R40378 S.n20494 S.n20493 0.054
R40379 S.n20401 S.n20400 0.054
R40380 S.n19883 S.n19882 0.054
R40381 S.n20277 S.n20276 0.054
R40382 S.n19029 S.n19028 0.054
R40383 S.n19409 S.n19408 0.054
R40384 S.n18163 S.n18162 0.054
R40385 S.n18522 S.n18521 0.054
R40386 S.n17274 S.n17273 0.054
R40387 S.n17622 S.n17621 0.054
R40388 S.n16372 S.n16371 0.054
R40389 S.n16699 S.n16698 0.054
R40390 S.n15448 S.n15447 0.054
R40391 S.n15764 S.n15763 0.054
R40392 S.n14511 S.n14510 0.054
R40393 S.n14806 S.n14805 0.054
R40394 S.n13552 S.n13551 0.054
R40395 S.n13836 S.n13835 0.054
R40396 S.n12580 S.n12579 0.054
R40397 S.n12843 S.n12842 0.054
R40398 S.n11586 S.n11585 0.054
R40399 S.n11838 S.n11837 0.054
R40400 S.n10579 S.n10578 0.054
R40401 S.n10810 S.n10809 0.054
R40402 S.n9550 S.n9549 0.054
R40403 S.n9770 S.n9769 0.054
R40404 S.n8508 S.n8507 0.054
R40405 S.n8707 S.n8706 0.054
R40406 S.n7444 S.n7443 0.054
R40407 S.n7632 S.n7631 0.054
R40408 S.n6367 S.n6366 0.054
R40409 S.n6534 S.n6533 0.054
R40410 S.n5267 S.n5266 0.054
R40411 S.n5423 S.n5422 0.054
R40412 S.n4154 S.n4153 0.054
R40413 S.n4289 S.n4288 0.054
R40414 S.n3028 S.n3027 0.054
R40415 S.n3152 S.n3151 0.054
R40416 S.n1868 S.n1867 0.054
R40417 S.n880 S.n879 0.054
R40418 S.n812 S.n811 0.054
R40419 S.n22357 S.n22356 0.054
R40420 S.n22716 S.n22715 0.054
R40421 S.n21351 S.n21350 0.054
R40422 S.n21267 S.n21266 0.054
R40423 S.n20830 S.n20829 0.054
R40424 S.n20851 S.n20850 0.054
R40425 S.n20195 S.n20194 0.054
R40426 S.n20213 S.n20212 0.054
R40427 S.n19325 S.n19324 0.054
R40428 S.n19343 S.n19342 0.054
R40429 S.n18443 S.n18442 0.054
R40430 S.n18461 S.n18460 0.054
R40431 S.n17538 S.n17537 0.054
R40432 S.n17556 S.n17555 0.054
R40433 S.n16620 S.n16619 0.054
R40434 S.n16638 S.n16637 0.054
R40435 S.n15680 S.n15679 0.054
R40436 S.n15698 S.n15697 0.054
R40437 S.n14727 S.n14726 0.054
R40438 S.n14745 S.n14744 0.054
R40439 S.n13752 S.n13751 0.054
R40440 S.n13770 S.n13769 0.054
R40441 S.n12764 S.n12763 0.054
R40442 S.n12782 S.n12781 0.054
R40443 S.n11754 S.n11753 0.054
R40444 S.n11772 S.n11771 0.054
R40445 S.n10731 S.n10730 0.054
R40446 S.n10749 S.n10748 0.054
R40447 S.n9686 S.n9685 0.054
R40448 S.n9704 S.n9703 0.054
R40449 S.n8628 S.n8627 0.054
R40450 S.n8646 S.n8645 0.054
R40451 S.n7548 S.n7547 0.054
R40452 S.n7566 S.n7565 0.054
R40453 S.n6455 S.n6454 0.054
R40454 S.n6473 S.n6472 0.054
R40455 S.n5339 S.n5338 0.054
R40456 S.n5357 S.n5356 0.054
R40457 S.n4210 S.n4209 0.054
R40458 S.n4228 S.n4227 0.054
R40459 S.n3069 S.n3068 0.054
R40460 S.n3087 S.n3086 0.054
R40461 S.n1888 S.n1887 0.054
R40462 S.n1934 S.n1933 0.054
R40463 S.n409 S.n408 0.054
R40464 S.n2143 S.n2142 0.054
R40465 S.n18486 S.n18485 0.054
R40466 S.n17172 S.n17171 0.054
R40467 S.n17771 S.n17770 0.054
R40468 S.n16272 S.n16271 0.054
R40469 S.n16844 S.n16843 0.054
R40470 S.n15348 S.n15347 0.054
R40471 S.n15909 S.n15908 0.054
R40472 S.n14411 S.n14410 0.054
R40473 S.n14951 S.n14950 0.054
R40474 S.n13452 S.n13451 0.054
R40475 S.n13981 S.n13980 0.054
R40476 S.n12480 S.n12479 0.054
R40477 S.n12988 S.n12987 0.054
R40478 S.n11486 S.n11485 0.054
R40479 S.n11983 S.n11982 0.054
R40480 S.n10479 S.n10478 0.054
R40481 S.n10955 S.n10954 0.054
R40482 S.n9450 S.n9449 0.054
R40483 S.n9915 S.n9914 0.054
R40484 S.n8408 S.n8407 0.054
R40485 S.n8852 S.n8851 0.054
R40486 S.n7344 S.n7343 0.054
R40487 S.n7777 S.n7776 0.054
R40488 S.n6267 S.n6266 0.054
R40489 S.n6679 S.n6678 0.054
R40490 S.n5167 S.n5166 0.054
R40491 S.n5569 S.n5568 0.054
R40492 S.n4055 S.n4054 0.054
R40493 S.n4434 S.n4433 0.054
R40494 S.n2928 S.n2927 0.054
R40495 S.n3296 S.n3295 0.054
R40496 S.n1760 S.n1759 0.054
R40497 S.n19 S.n18 0.054
R40498 S.n19373 S.n19372 0.054
R40499 S.n18080 S.n18079 0.054
R40500 S.n18639 S.n18638 0.054
R40501 S.n17191 S.n17190 0.054
R40502 S.n17739 S.n17738 0.054
R40503 S.n16289 S.n16288 0.054
R40504 S.n16812 S.n16811 0.054
R40505 S.n15365 S.n15364 0.054
R40506 S.n15877 S.n15876 0.054
R40507 S.n14428 S.n14427 0.054
R40508 S.n14919 S.n14918 0.054
R40509 S.n13469 S.n13468 0.054
R40510 S.n13949 S.n13948 0.054
R40511 S.n12497 S.n12496 0.054
R40512 S.n12956 S.n12955 0.054
R40513 S.n11503 S.n11502 0.054
R40514 S.n11951 S.n11950 0.054
R40515 S.n10496 S.n10495 0.054
R40516 S.n10923 S.n10922 0.054
R40517 S.n9467 S.n9466 0.054
R40518 S.n9883 S.n9882 0.054
R40519 S.n8425 S.n8424 0.054
R40520 S.n8820 S.n8819 0.054
R40521 S.n7361 S.n7360 0.054
R40522 S.n7745 S.n7744 0.054
R40523 S.n6284 S.n6283 0.054
R40524 S.n6647 S.n6646 0.054
R40525 S.n5184 S.n5183 0.054
R40526 S.n5537 S.n5536 0.054
R40527 S.n4072 S.n4071 0.054
R40528 S.n4402 S.n4401 0.054
R40529 S.n2945 S.n2944 0.054
R40530 S.n3265 S.n3264 0.054
R40531 S.n1779 S.n1778 0.054
R40532 S.n1802 S.n1801 0.054
R40533 S.n2085 S.n2084 0.054
R40534 S.n818 S.n817 0.054
R40535 S.n841 S.n840 0.054
R40536 S.n3236 S.n3235 0.054
R40537 S.n4373 S.n4372 0.054
R40538 S.n5508 S.n5507 0.054
R40539 S.n6618 S.n6617 0.054
R40540 S.n7716 S.n7715 0.054
R40541 S.n8791 S.n8790 0.054
R40542 S.n9854 S.n9853 0.054
R40543 S.n10894 S.n10893 0.054
R40544 S.n11922 S.n11921 0.054
R40545 S.n12927 S.n12926 0.054
R40546 S.n13920 S.n13919 0.054
R40547 S.n14890 S.n14889 0.054
R40548 S.n15848 S.n15847 0.054
R40549 S.n16783 S.n16782 0.054
R40550 S.n17706 S.n17705 0.054
R40551 S.n18606 S.n18605 0.054
R40552 S.n19496 S.n19495 0.054
R40553 S.n20241 S.n20240 0.054
R40554 S.n18964 S.n18963 0.054
R40555 S.n18099 S.n18098 0.054
R40556 S.n17210 S.n17209 0.054
R40557 S.n16308 S.n16307 0.054
R40558 S.n15384 S.n15383 0.054
R40559 S.n14447 S.n14446 0.054
R40560 S.n13488 S.n13487 0.054
R40561 S.n12516 S.n12515 0.054
R40562 S.n11522 S.n11521 0.054
R40563 S.n10515 S.n10514 0.054
R40564 S.n9486 S.n9485 0.054
R40565 S.n8444 S.n8443 0.054
R40566 S.n7380 S.n7379 0.054
R40567 S.n6303 S.n6302 0.054
R40568 S.n5203 S.n5202 0.054
R40569 S.n4091 S.n4090 0.054
R40570 S.n2964 S.n2963 0.054
R40571 S.n2051 S.n2050 0.054
R40572 S.n770 S.n769 0.054
R40573 S.n1331 S.n1330 0.054
R40574 S.n20430 S.n20429 0.054
R40575 S.n19842 S.n19841 0.054
R40576 S.n20336 S.n20335 0.054
R40577 S.n18990 S.n18989 0.054
R40578 S.n19464 S.n19463 0.054
R40579 S.n18124 S.n18123 0.054
R40580 S.n18574 S.n18573 0.054
R40581 S.n17235 S.n17234 0.054
R40582 S.n17674 S.n17673 0.054
R40583 S.n16333 S.n16332 0.054
R40584 S.n16751 S.n16750 0.054
R40585 S.n15409 S.n15408 0.054
R40586 S.n15816 S.n15815 0.054
R40587 S.n14472 S.n14471 0.054
R40588 S.n14858 S.n14857 0.054
R40589 S.n13513 S.n13512 0.054
R40590 S.n13888 S.n13887 0.054
R40591 S.n12541 S.n12540 0.054
R40592 S.n12895 S.n12894 0.054
R40593 S.n11547 S.n11546 0.054
R40594 S.n11890 S.n11889 0.054
R40595 S.n10540 S.n10539 0.054
R40596 S.n10862 S.n10861 0.054
R40597 S.n9511 S.n9510 0.054
R40598 S.n9822 S.n9821 0.054
R40599 S.n8469 S.n8468 0.054
R40600 S.n8759 S.n8758 0.054
R40601 S.n7405 S.n7404 0.054
R40602 S.n7684 S.n7683 0.054
R40603 S.n6328 S.n6327 0.054
R40604 S.n6586 S.n6585 0.054
R40605 S.n5228 S.n5227 0.054
R40606 S.n5476 S.n5475 0.054
R40607 S.n4116 S.n4115 0.054
R40608 S.n4341 S.n4340 0.054
R40609 S.n2989 S.n2988 0.054
R40610 S.n3204 S.n3203 0.054
R40611 S.n1826 S.n1825 0.054
R40612 S.n2018 S.n2017 0.054
R40613 S.n789 S.n788 0.054
R40614 S.n1848 S.n1847 0.054
R40615 S.n3172 S.n3171 0.054
R40616 S.n3009 S.n3008 0.054
R40617 S.n4309 S.n4308 0.054
R40618 S.n4135 S.n4134 0.054
R40619 S.n5444 S.n5443 0.054
R40620 S.n5248 S.n5247 0.054
R40621 S.n6554 S.n6553 0.054
R40622 S.n6348 S.n6347 0.054
R40623 S.n7652 S.n7651 0.054
R40624 S.n7425 S.n7424 0.054
R40625 S.n8727 S.n8726 0.054
R40626 S.n8489 S.n8488 0.054
R40627 S.n9790 S.n9789 0.054
R40628 S.n9531 S.n9530 0.054
R40629 S.n10830 S.n10829 0.054
R40630 S.n10560 S.n10559 0.054
R40631 S.n11858 S.n11857 0.054
R40632 S.n11567 S.n11566 0.054
R40633 S.n12863 S.n12862 0.054
R40634 S.n12561 S.n12560 0.054
R40635 S.n13856 S.n13855 0.054
R40636 S.n13533 S.n13532 0.054
R40637 S.n14826 S.n14825 0.054
R40638 S.n14492 S.n14491 0.054
R40639 S.n15784 S.n15783 0.054
R40640 S.n15429 S.n15428 0.054
R40641 S.n16719 S.n16718 0.054
R40642 S.n16353 S.n16352 0.054
R40643 S.n17642 S.n17641 0.054
R40644 S.n17255 S.n17254 0.054
R40645 S.n18542 S.n18541 0.054
R40646 S.n18144 S.n18143 0.054
R40647 S.n19429 S.n19428 0.054
R40648 S.n19010 S.n19009 0.054
R40649 S.n20301 S.n20300 0.054
R40650 S.n19864 S.n19863 0.054
R40651 S.n20369 S.n20368 0.054
R40652 S.n20475 S.n20474 0.054
R40653 S.n21248 S.n21247 0.054
R40654 S.n867 S.n866 0.054
R40655 S.n2113 S.n2112 0.054
R40656 S.n746 S.n745 0.054
R40657 S.n729 S.n728 0.054
R40658 S.n377 S.n376 0.054
R40659 S.n2202 S.n2201 0.054
R40660 S.n16663 S.n16662 0.054
R40661 S.n15310 S.n15309 0.054
R40662 S.n15974 S.n15973 0.054
R40663 S.n14375 S.n14374 0.054
R40664 S.n15012 S.n15011 0.054
R40665 S.n13416 S.n13415 0.054
R40666 S.n14042 S.n14041 0.054
R40667 S.n12444 S.n12443 0.054
R40668 S.n13049 S.n13048 0.054
R40669 S.n11450 S.n11449 0.054
R40670 S.n12044 S.n12043 0.054
R40671 S.n10443 S.n10442 0.054
R40672 S.n11016 S.n11015 0.054
R40673 S.n9414 S.n9413 0.054
R40674 S.n9976 S.n9975 0.054
R40675 S.n8372 S.n8371 0.054
R40676 S.n8913 S.n8912 0.054
R40677 S.n7308 S.n7307 0.054
R40678 S.n7838 S.n7837 0.054
R40679 S.n6231 S.n6230 0.054
R40680 S.n6740 S.n6739 0.054
R40681 S.n5131 S.n5130 0.054
R40682 S.n5630 S.n5629 0.054
R40683 S.n4019 S.n4018 0.054
R40684 S.n4495 S.n4494 0.054
R40685 S.n2892 S.n2891 0.054
R40686 S.n3356 S.n3355 0.054
R40687 S.n1723 S.n1722 0.054
R40688 S.n66 S.n65 0.054
R40689 S.n17586 S.n17585 0.054
R40690 S.n16253 S.n16252 0.054
R40691 S.n16877 S.n16876 0.054
R40692 S.n15329 S.n15328 0.054
R40693 S.n15942 S.n15941 0.054
R40694 S.n14392 S.n14391 0.054
R40695 S.n14980 S.n14979 0.054
R40696 S.n13433 S.n13432 0.054
R40697 S.n14010 S.n14009 0.054
R40698 S.n12461 S.n12460 0.054
R40699 S.n13017 S.n13016 0.054
R40700 S.n11467 S.n11466 0.054
R40701 S.n12012 S.n12011 0.054
R40702 S.n10460 S.n10459 0.054
R40703 S.n10984 S.n10983 0.054
R40704 S.n9431 S.n9430 0.054
R40705 S.n9944 S.n9943 0.054
R40706 S.n8389 S.n8388 0.054
R40707 S.n8881 S.n8880 0.054
R40708 S.n7325 S.n7324 0.054
R40709 S.n7806 S.n7805 0.054
R40710 S.n6248 S.n6247 0.054
R40711 S.n6708 S.n6707 0.054
R40712 S.n5148 S.n5147 0.054
R40713 S.n5598 S.n5597 0.054
R40714 S.n4036 S.n4035 0.054
R40715 S.n4463 S.n4462 0.054
R40716 S.n2909 S.n2908 0.054
R40717 S.n3325 S.n3324 0.054
R40718 S.n1740 S.n1739 0.054
R40719 S.n2172 S.n2171 0.054
R40720 S.n711 S.n710 0.054
R40721 S.n694 S.n693 0.054
R40722 S.n345 S.n344 0.054
R40723 S.n2261 S.n2260 0.054
R40724 S.n14770 S.n14769 0.054
R40725 S.n13378 S.n13377 0.054
R40726 S.n14107 S.n14106 0.054
R40727 S.n12408 S.n12407 0.054
R40728 S.n13110 S.n13109 0.054
R40729 S.n11414 S.n11413 0.054
R40730 S.n12105 S.n12104 0.054
R40731 S.n10407 S.n10406 0.054
R40732 S.n11077 S.n11076 0.054
R40733 S.n9378 S.n9377 0.054
R40734 S.n10037 S.n10036 0.054
R40735 S.n8336 S.n8335 0.054
R40736 S.n8974 S.n8973 0.054
R40737 S.n7272 S.n7271 0.054
R40738 S.n7899 S.n7898 0.054
R40739 S.n6195 S.n6194 0.054
R40740 S.n6801 S.n6800 0.054
R40741 S.n5095 S.n5094 0.054
R40742 S.n5691 S.n5690 0.054
R40743 S.n3983 S.n3982 0.054
R40744 S.n4556 S.n4555 0.054
R40745 S.n2856 S.n2855 0.054
R40746 S.n3416 S.n3415 0.054
R40747 S.n1686 S.n1685 0.054
R40748 S.n98 S.n97 0.054
R40749 S.n15728 S.n15727 0.054
R40750 S.n14356 S.n14355 0.054
R40751 S.n15045 S.n15044 0.054
R40752 S.n13397 S.n13396 0.054
R40753 S.n14075 S.n14074 0.054
R40754 S.n12425 S.n12424 0.054
R40755 S.n13078 S.n13077 0.054
R40756 S.n11431 S.n11430 0.054
R40757 S.n12073 S.n12072 0.054
R40758 S.n10424 S.n10423 0.054
R40759 S.n11045 S.n11044 0.054
R40760 S.n9395 S.n9394 0.054
R40761 S.n10005 S.n10004 0.054
R40762 S.n8353 S.n8352 0.054
R40763 S.n8942 S.n8941 0.054
R40764 S.n7289 S.n7288 0.054
R40765 S.n7867 S.n7866 0.054
R40766 S.n6212 S.n6211 0.054
R40767 S.n6769 S.n6768 0.054
R40768 S.n5112 S.n5111 0.054
R40769 S.n5659 S.n5658 0.054
R40770 S.n4000 S.n3999 0.054
R40771 S.n4524 S.n4523 0.054
R40772 S.n2873 S.n2872 0.054
R40773 S.n3385 S.n3384 0.054
R40774 S.n1703 S.n1702 0.054
R40775 S.n2231 S.n2230 0.054
R40776 S.n676 S.n675 0.054
R40777 S.n659 S.n658 0.054
R40778 S.n313 S.n312 0.054
R40779 S.n2320 S.n2319 0.054
R40780 S.n12807 S.n12806 0.054
R40781 S.n11376 S.n11375 0.054
R40782 S.n12170 S.n12169 0.054
R40783 S.n10371 S.n10370 0.054
R40784 S.n11138 S.n11137 0.054
R40785 S.n9342 S.n9341 0.054
R40786 S.n10098 S.n10097 0.054
R40787 S.n8300 S.n8299 0.054
R40788 S.n9035 S.n9034 0.054
R40789 S.n7236 S.n7235 0.054
R40790 S.n7960 S.n7959 0.054
R40791 S.n6159 S.n6158 0.054
R40792 S.n6862 S.n6861 0.054
R40793 S.n5059 S.n5058 0.054
R40794 S.n5752 S.n5751 0.054
R40795 S.n3947 S.n3946 0.054
R40796 S.n4617 S.n4616 0.054
R40797 S.n2820 S.n2819 0.054
R40798 S.n3476 S.n3475 0.054
R40799 S.n1649 S.n1648 0.054
R40800 S.n985 S.n984 0.054
R40801 S.n13800 S.n13799 0.054
R40802 S.n12389 S.n12388 0.054
R40803 S.n13143 S.n13142 0.054
R40804 S.n11395 S.n11394 0.054
R40805 S.n12138 S.n12137 0.054
R40806 S.n10388 S.n10387 0.054
R40807 S.n11106 S.n11105 0.054
R40808 S.n9359 S.n9358 0.054
R40809 S.n10066 S.n10065 0.054
R40810 S.n8317 S.n8316 0.054
R40811 S.n9003 S.n9002 0.054
R40812 S.n7253 S.n7252 0.054
R40813 S.n7928 S.n7927 0.054
R40814 S.n6176 S.n6175 0.054
R40815 S.n6830 S.n6829 0.054
R40816 S.n5076 S.n5075 0.054
R40817 S.n5720 S.n5719 0.054
R40818 S.n3964 S.n3963 0.054
R40819 S.n4585 S.n4584 0.054
R40820 S.n2837 S.n2836 0.054
R40821 S.n3445 S.n3444 0.054
R40822 S.n1666 S.n1665 0.054
R40823 S.n2290 S.n2289 0.054
R40824 S.n641 S.n640 0.054
R40825 S.n624 S.n623 0.054
R40826 S.n281 S.n280 0.054
R40827 S.n2379 S.n2378 0.054
R40828 S.n10774 S.n10773 0.054
R40829 S.n9304 S.n9303 0.054
R40830 S.n10163 S.n10162 0.054
R40831 S.n8264 S.n8263 0.054
R40832 S.n9096 S.n9095 0.054
R40833 S.n7200 S.n7199 0.054
R40834 S.n8021 S.n8020 0.054
R40835 S.n6123 S.n6122 0.054
R40836 S.n6923 S.n6922 0.054
R40837 S.n5023 S.n5022 0.054
R40838 S.n5813 S.n5812 0.054
R40839 S.n3911 S.n3910 0.054
R40840 S.n4678 S.n4677 0.054
R40841 S.n2784 S.n2783 0.054
R40842 S.n3536 S.n3535 0.054
R40843 S.n1612 S.n1611 0.054
R40844 S.n1017 S.n1016 0.054
R40845 S.n11802 S.n11801 0.054
R40846 S.n10352 S.n10351 0.054
R40847 S.n11171 S.n11170 0.054
R40848 S.n9323 S.n9322 0.054
R40849 S.n10131 S.n10130 0.054
R40850 S.n8281 S.n8280 0.054
R40851 S.n9064 S.n9063 0.054
R40852 S.n7217 S.n7216 0.054
R40853 S.n7989 S.n7988 0.054
R40854 S.n6140 S.n6139 0.054
R40855 S.n6891 S.n6890 0.054
R40856 S.n5040 S.n5039 0.054
R40857 S.n5781 S.n5780 0.054
R40858 S.n3928 S.n3927 0.054
R40859 S.n4646 S.n4645 0.054
R40860 S.n2801 S.n2800 0.054
R40861 S.n3505 S.n3504 0.054
R40862 S.n1629 S.n1628 0.054
R40863 S.n2349 S.n2348 0.054
R40864 S.n606 S.n605 0.054
R40865 S.n589 S.n588 0.054
R40866 S.n223 S.n222 0.054
R40867 S.n2438 S.n2437 0.054
R40868 S.n8671 S.n8670 0.054
R40869 S.n7162 S.n7161 0.054
R40870 S.n8086 S.n8085 0.054
R40871 S.n6087 S.n6086 0.054
R40872 S.n6984 S.n6983 0.054
R40873 S.n4987 S.n4986 0.054
R40874 S.n5874 S.n5873 0.054
R40875 S.n3875 S.n3874 0.054
R40876 S.n4739 S.n4738 0.054
R40877 S.n2748 S.n2747 0.054
R40878 S.n3596 S.n3595 0.054
R40879 S.n1575 S.n1574 0.054
R40880 S.n1049 S.n1048 0.054
R40881 S.n9734 S.n9733 0.054
R40882 S.n8245 S.n8244 0.054
R40883 S.n9129 S.n9128 0.054
R40884 S.n7181 S.n7180 0.054
R40885 S.n8054 S.n8053 0.054
R40886 S.n6104 S.n6103 0.054
R40887 S.n6952 S.n6951 0.054
R40888 S.n5004 S.n5003 0.054
R40889 S.n5842 S.n5841 0.054
R40890 S.n3892 S.n3891 0.054
R40891 S.n4707 S.n4706 0.054
R40892 S.n2765 S.n2764 0.054
R40893 S.n3565 S.n3564 0.054
R40894 S.n1592 S.n1591 0.054
R40895 S.n2408 S.n2407 0.054
R40896 S.n571 S.n570 0.054
R40897 S.n554 S.n553 0.054
R40898 S.n217 S.n216 0.054
R40899 S.n2497 S.n2496 0.054
R40900 S.n6498 S.n6497 0.054
R40901 S.n4949 S.n4948 0.054
R40902 S.n5939 S.n5938 0.054
R40903 S.n3839 S.n3838 0.054
R40904 S.n4800 S.n4799 0.054
R40905 S.n2712 S.n2711 0.054
R40906 S.n3656 S.n3655 0.054
R40907 S.n1538 S.n1537 0.054
R40908 S.n1081 S.n1080 0.054
R40909 S.n7596 S.n7595 0.054
R40910 S.n6068 S.n6067 0.054
R40911 S.n7017 S.n7016 0.054
R40912 S.n4968 S.n4967 0.054
R40913 S.n5907 S.n5906 0.054
R40914 S.n3856 S.n3855 0.054
R40915 S.n4768 S.n4767 0.054
R40916 S.n2729 S.n2728 0.054
R40917 S.n3625 S.n3624 0.054
R40918 S.n1555 S.n1554 0.054
R40919 S.n2467 S.n2466 0.054
R40920 S.n536 S.n535 0.054
R40921 S.n519 S.n518 0.054
R40922 S.n185 S.n184 0.054
R40923 S.n2556 S.n2555 0.054
R40924 S.n4253 S.n4252 0.054
R40925 S.n2674 S.n2673 0.054
R40926 S.n3720 S.n3719 0.054
R40927 S.n1501 S.n1500 0.054
R40928 S.n1113 S.n1112 0.054
R40929 S.n5387 S.n5386 0.054
R40930 S.n3820 S.n3819 0.054
R40931 S.n4833 S.n4832 0.054
R40932 S.n2693 S.n2692 0.054
R40933 S.n3689 S.n3688 0.054
R40934 S.n1518 S.n1517 0.054
R40935 S.n2526 S.n2525 0.054
R40936 S.n501 S.n500 0.054
R40937 S.n484 S.n483 0.054
R40938 S.n153 S.n152 0.054
R40939 S.n1957 S.n1956 0.054
R40940 S.n1151 S.n1150 0.054
R40941 S.n3117 S.n3116 0.054
R40942 S.n1481 S.n1480 0.054
R40943 S.n2589 S.n2588 0.054
R40944 S.n466 S.n465 0.054
R40945 S.n450 S.n449 0.054
R40946 S.n948 S.n947 0.054
R40947 S.n22771 S.n22770 0.054
R40948 S.n21331 S.n21330 0.054
R40949 S.n1377 S.n1376 0.053
R40950 S.n22981 S.n22980 0.053
R40951 S.n23008 S.n22805 0.053
R40952 S.n22285 S.n22283 0.052
R40953 S.n428 S.n427 0.052
R40954 S.n1456 S.n1455 0.052
R40955 S.n2650 S.n2649 0.052
R40956 S.n3795 S.n3794 0.052
R40957 S.n4925 S.n4924 0.052
R40958 S.n6043 S.n6042 0.052
R40959 S.n7138 S.n7137 0.052
R40960 S.n8220 S.n8219 0.052
R40961 S.n9280 S.n9279 0.052
R40962 S.n10327 S.n10326 0.052
R40963 S.n11352 S.n11351 0.052
R40964 S.n12364 S.n12363 0.052
R40965 S.n13354 S.n13353 0.052
R40966 S.n14331 S.n14330 0.052
R40967 S.n15286 S.n15285 0.052
R40968 S.n16228 S.n16227 0.052
R40969 S.n17148 S.n17147 0.052
R40970 S.n18055 S.n18054 0.052
R40971 S.n18940 S.n18939 0.052
R40972 S.n19810 S.n19809 0.052
R40973 S.n20448 S.n20447 0.052
R40974 S.n21292 S.n21291 0.052
R40975 S.n2617 S.n2616 0.052
R40976 S.n1917 S.n1916 0.052
R40977 S.n909 S.n907 0.051
R40978 S.n20236 S.n20234 0.051
R40979 S.n19349 S.n19348 0.051
R40980 S.n18481 S.n18479 0.051
R40981 S.n17562 S.n17561 0.051
R40982 S.n16658 S.n16656 0.051
R40983 S.n15704 S.n15703 0.051
R40984 S.n14765 S.n14763 0.051
R40985 S.n13776 S.n13775 0.051
R40986 S.n12802 S.n12800 0.051
R40987 S.n11778 S.n11777 0.051
R40988 S.n10769 S.n10767 0.051
R40989 S.n9710 S.n9709 0.051
R40990 S.n8666 S.n8664 0.051
R40991 S.n7572 S.n7571 0.051
R40992 S.n6493 S.n6491 0.051
R40993 S.n5363 S.n5362 0.051
R40994 S.n4248 S.n4246 0.051
R40995 S.n1952 S.n1950 0.051
R40996 S.n3093 S.n3092 0.051
R40997 S.n925 S.n923 0.051
R40998 S.n22987 S.n22986 0.051
R40999 S.n22989 S.n22988 0.051
R41000 S.n957 S.n956 0.051
R41001 S.n23003 S.n23002 0.051
R41002 S.n23005 S.n23004 0.051
R41003 S.n959 S.n958 0.051
R41004 S.n1809 S.n1808 0.051
R41005 S.n2971 S.n2970 0.051
R41006 S.n4098 S.n4097 0.051
R41007 S.n5210 S.n5209 0.051
R41008 S.n6310 S.n6309 0.051
R41009 S.n7387 S.n7386 0.051
R41010 S.n8451 S.n8450 0.051
R41011 S.n9493 S.n9492 0.051
R41012 S.n10522 S.n10521 0.051
R41013 S.n11529 S.n11528 0.051
R41014 S.n12523 S.n12522 0.051
R41015 S.n13495 S.n13494 0.051
R41016 S.n14454 S.n14453 0.051
R41017 S.n15391 S.n15390 0.051
R41018 S.n16315 S.n16314 0.051
R41019 S.n17217 S.n17216 0.051
R41020 S.n18106 S.n18105 0.051
R41021 S.n18971 S.n18970 0.051
R41022 S.n19823 S.n19822 0.051
R41023 S.n765 S.n764 0.051
R41024 S.n20398 S.n20397 0.05
R41025 S.n21217 S.n21216 0.05
R41026 S.n22741 S.n22740 0.05
R41027 S.n18600 S.n18599 0.05
R41028 S.n19490 S.n19489 0.05
R41029 S.n20238 S.n20237 0.05
R41030 S.n20295 S.n20282 0.05
R41031 S.n20366 S.n20353 0.05
R41032 S.n21242 S.n21229 0.05
R41033 S.n858 S.n857 0.05
R41034 S.n19367 S.n19364 0.05
R41035 S.n19370 S.n19351 0.05
R41036 S.n18633 S.n18611 0.05
R41037 S.n17733 S.n17711 0.05
R41038 S.n16838 S.n16837 0.05
R41039 S.n17765 S.n17764 0.05
R41040 S.n18483 S.n18482 0.05
R41041 S.n17580 S.n17577 0.05
R41042 S.n17583 S.n17564 0.05
R41043 S.n16871 S.n16849 0.05
R41044 S.n15936 S.n15914 0.05
R41045 S.n15006 S.n15005 0.05
R41046 S.n15968 S.n15967 0.05
R41047 S.n16660 S.n16659 0.05
R41048 S.n15720 S.n15719 0.05
R41049 S.n15725 S.n15706 0.05
R41050 S.n15039 S.n15017 0.05
R41051 S.n14069 S.n14047 0.05
R41052 S.n13104 S.n13103 0.05
R41053 S.n14101 S.n14100 0.05
R41054 S.n14767 S.n14766 0.05
R41055 S.n13792 S.n13791 0.05
R41056 S.n13797 S.n13778 0.05
R41057 S.n13137 S.n13115 0.05
R41058 S.n12132 S.n12110 0.05
R41059 S.n11132 S.n11131 0.05
R41060 S.n12164 S.n12163 0.05
R41061 S.n12804 S.n12803 0.05
R41062 S.n11794 S.n11793 0.05
R41063 S.n11799 S.n11780 0.05
R41064 S.n11165 S.n11143 0.05
R41065 S.n10125 S.n10103 0.05
R41066 S.n9090 S.n9089 0.05
R41067 S.n10157 S.n10156 0.05
R41068 S.n10771 S.n10770 0.05
R41069 S.n9728 S.n9725 0.05
R41070 S.n9731 S.n9712 0.05
R41071 S.n9123 S.n9101 0.05
R41072 S.n8048 S.n8026 0.05
R41073 S.n6978 S.n6977 0.05
R41074 S.n8080 S.n8079 0.05
R41075 S.n8668 S.n8667 0.05
R41076 S.n7590 S.n7587 0.05
R41077 S.n7593 S.n7574 0.05
R41078 S.n7011 S.n6989 0.05
R41079 S.n5901 S.n5879 0.05
R41080 S.n4794 S.n4793 0.05
R41081 S.n5933 S.n5932 0.05
R41082 S.n6495 S.n6494 0.05
R41083 S.n5381 S.n5378 0.05
R41084 S.n5384 S.n5365 0.05
R41085 S.n4827 S.n4805 0.05
R41086 S.n3683 S.n3661 0.05
R41087 S.n2550 S.n2549 0.05
R41088 S.n3714 S.n3713 0.05
R41089 S.n4250 S.n4249 0.05
R41090 S.n1954 S.n1953 0.05
R41091 S.n3111 S.n3108 0.05
R41092 S.n3114 S.n3095 0.05
R41093 S.n2583 S.n2561 0.05
R41094 S.n942 S.n926 0.05
R41095 S.n825 S.n824 0.05
R41096 S.n22332 S.n22331 0.05
R41097 S.n21190 S.n21189 0.05
R41098 S.n892 S.n891 0.049
R41099 S.n803 S.n802 0.049
R41100 S.n1815 S.n1814 0.049
R41101 S.n2978 S.n2977 0.049
R41102 S.n4105 S.n4104 0.049
R41103 S.n5217 S.n5216 0.049
R41104 S.n6317 S.n6316 0.049
R41105 S.n7394 S.n7393 0.049
R41106 S.n8458 S.n8457 0.049
R41107 S.n9500 S.n9499 0.049
R41108 S.n10529 S.n10528 0.049
R41109 S.n11536 S.n11535 0.049
R41110 S.n12530 S.n12529 0.049
R41111 S.n13502 S.n13501 0.049
R41112 S.n14461 S.n14460 0.049
R41113 S.n15398 S.n15397 0.049
R41114 S.n16322 S.n16321 0.049
R41115 S.n17224 S.n17223 0.049
R41116 S.n18113 S.n18112 0.049
R41117 S.n18978 S.n18977 0.049
R41118 S.n19830 S.n19829 0.049
R41119 S.n763 S.n762 0.049
R41120 S.n783 S.n782 0.049
R41121 S.n22756 S.n22751 0.049
R41122 S.n21170 S.n21169 0.048
R41123 S.n1913 S.n1912 0.048
R41124 S.n21980 S.n21191 0.048
R41125 S.n2073 S.n2068 0.048
R41126 S.n19474 S.n19473 0.048
R41127 S.n18584 S.n18583 0.048
R41128 S.n17684 S.n17683 0.048
R41129 S.n16761 S.n16760 0.048
R41130 S.n15826 S.n15825 0.048
R41131 S.n14868 S.n14867 0.048
R41132 S.n13898 S.n13897 0.048
R41133 S.n12905 S.n12904 0.048
R41134 S.n11900 S.n11899 0.048
R41135 S.n10872 S.n10871 0.048
R41136 S.n9832 S.n9831 0.048
R41137 S.n8769 S.n8768 0.048
R41138 S.n7694 S.n7693 0.048
R41139 S.n6596 S.n6595 0.048
R41140 S.n5486 S.n5485 0.048
R41141 S.n4351 S.n4350 0.048
R41142 S.n3215 S.n3214 0.048
R41143 S.n20183 S.n20181 0.047
R41144 S.n21133 S.n21129 0.047
R41145 S.n22640 S.n22635 0.047
R41146 S.n22010 S.n22006 0.047
R41147 S.n21617 S.n21612 0.047
R41148 S.n21942 S.n21938 0.047
R41149 S.n20794 S.n20789 0.047
R41150 S.n21172 S.n21146 0.047
R41151 S.n22656 S.n22654 0.047
R41152 S.n21995 S.n21993 0.047
R41153 S.n21638 S.n21636 0.047
R41154 S.n21962 S.n21959 0.047
R41155 S.n20818 S.n20813 0.047
R41156 S.n20344 S.n20341 0.047
R41157 S.n19313 S.n19311 0.047
R41158 S.n19533 S.n19529 0.047
R41159 S.n22624 S.n22619 0.047
R41160 S.n22025 S.n22021 0.047
R41161 S.n21601 S.n21596 0.047
R41162 S.n21927 S.n21923 0.047
R41163 S.n20778 S.n20773 0.047
R41164 S.n21117 S.n21113 0.047
R41165 S.n20167 S.n20162 0.047
R41166 S.n19504 S.n19501 0.047
R41167 S.n18431 S.n18429 0.047
R41168 S.n18676 S.n18672 0.047
R41169 S.n22608 S.n22603 0.047
R41170 S.n22040 S.n22036 0.047
R41171 S.n21585 S.n21580 0.047
R41172 S.n21912 S.n21908 0.047
R41173 S.n20762 S.n20757 0.047
R41174 S.n21102 S.n21098 0.047
R41175 S.n20151 S.n20146 0.047
R41176 S.n19548 S.n19544 0.047
R41177 S.n19297 S.n19292 0.047
R41178 S.n18647 S.n18644 0.047
R41179 S.n17526 S.n17524 0.047
R41180 S.n17808 S.n17804 0.047
R41181 S.n22592 S.n22587 0.047
R41182 S.n22055 S.n22051 0.047
R41183 S.n21569 S.n21564 0.047
R41184 S.n21897 S.n21893 0.047
R41185 S.n20746 S.n20741 0.047
R41186 S.n21087 S.n21083 0.047
R41187 S.n20135 S.n20130 0.047
R41188 S.n19563 S.n19559 0.047
R41189 S.n19281 S.n19276 0.047
R41190 S.n18691 S.n18687 0.047
R41191 S.n18415 S.n18410 0.047
R41192 S.n17779 S.n17776 0.047
R41193 S.n16608 S.n16606 0.047
R41194 S.n16914 S.n16910 0.047
R41195 S.n22576 S.n22571 0.047
R41196 S.n22070 S.n22066 0.047
R41197 S.n21553 S.n21548 0.047
R41198 S.n21882 S.n21878 0.047
R41199 S.n20730 S.n20725 0.047
R41200 S.n21072 S.n21068 0.047
R41201 S.n20119 S.n20114 0.047
R41202 S.n19578 S.n19574 0.047
R41203 S.n19265 S.n19260 0.047
R41204 S.n18706 S.n18702 0.047
R41205 S.n18399 S.n18394 0.047
R41206 S.n17823 S.n17819 0.047
R41207 S.n17510 S.n17505 0.047
R41208 S.n16885 S.n16882 0.047
R41209 S.n15668 S.n15666 0.047
R41210 S.n16011 S.n16007 0.047
R41211 S.n22560 S.n22555 0.047
R41212 S.n22085 S.n22081 0.047
R41213 S.n21537 S.n21532 0.047
R41214 S.n21867 S.n21863 0.047
R41215 S.n20714 S.n20709 0.047
R41216 S.n21057 S.n21053 0.047
R41217 S.n20103 S.n20098 0.047
R41218 S.n19593 S.n19589 0.047
R41219 S.n19249 S.n19244 0.047
R41220 S.n18721 S.n18717 0.047
R41221 S.n18383 S.n18378 0.047
R41222 S.n17838 S.n17834 0.047
R41223 S.n17494 S.n17489 0.047
R41224 S.n16929 S.n16925 0.047
R41225 S.n16592 S.n16587 0.047
R41226 S.n15982 S.n15979 0.047
R41227 S.n14715 S.n14713 0.047
R41228 S.n15082 S.n15078 0.047
R41229 S.n22544 S.n22539 0.047
R41230 S.n22100 S.n22096 0.047
R41231 S.n21521 S.n21516 0.047
R41232 S.n21852 S.n21848 0.047
R41233 S.n20698 S.n20693 0.047
R41234 S.n21042 S.n21038 0.047
R41235 S.n20087 S.n20082 0.047
R41236 S.n19608 S.n19604 0.047
R41237 S.n19233 S.n19228 0.047
R41238 S.n18736 S.n18732 0.047
R41239 S.n18367 S.n18362 0.047
R41240 S.n17853 S.n17849 0.047
R41241 S.n17478 S.n17473 0.047
R41242 S.n16944 S.n16940 0.047
R41243 S.n16576 S.n16571 0.047
R41244 S.n16026 S.n16022 0.047
R41245 S.n15652 S.n15647 0.047
R41246 S.n15053 S.n15050 0.047
R41247 S.n13740 S.n13738 0.047
R41248 S.n14144 S.n14140 0.047
R41249 S.n22528 S.n22523 0.047
R41250 S.n22115 S.n22111 0.047
R41251 S.n21505 S.n21500 0.047
R41252 S.n21837 S.n21833 0.047
R41253 S.n20682 S.n20677 0.047
R41254 S.n21027 S.n21023 0.047
R41255 S.n20071 S.n20066 0.047
R41256 S.n19623 S.n19619 0.047
R41257 S.n19217 S.n19212 0.047
R41258 S.n18751 S.n18747 0.047
R41259 S.n18351 S.n18346 0.047
R41260 S.n17868 S.n17864 0.047
R41261 S.n17462 S.n17457 0.047
R41262 S.n16959 S.n16955 0.047
R41263 S.n16560 S.n16555 0.047
R41264 S.n16041 S.n16037 0.047
R41265 S.n15636 S.n15631 0.047
R41266 S.n15097 S.n15093 0.047
R41267 S.n14699 S.n14694 0.047
R41268 S.n14115 S.n14112 0.047
R41269 S.n12752 S.n12750 0.047
R41270 S.n13180 S.n13176 0.047
R41271 S.n22512 S.n22507 0.047
R41272 S.n22130 S.n22126 0.047
R41273 S.n21489 S.n21484 0.047
R41274 S.n21822 S.n21818 0.047
R41275 S.n20666 S.n20661 0.047
R41276 S.n21012 S.n21008 0.047
R41277 S.n20055 S.n20050 0.047
R41278 S.n19638 S.n19634 0.047
R41279 S.n19201 S.n19196 0.047
R41280 S.n18766 S.n18762 0.047
R41281 S.n18335 S.n18330 0.047
R41282 S.n17883 S.n17879 0.047
R41283 S.n17446 S.n17441 0.047
R41284 S.n16974 S.n16970 0.047
R41285 S.n16544 S.n16539 0.047
R41286 S.n16056 S.n16052 0.047
R41287 S.n15620 S.n15615 0.047
R41288 S.n15112 S.n15108 0.047
R41289 S.n14683 S.n14678 0.047
R41290 S.n14159 S.n14155 0.047
R41291 S.n13724 S.n13719 0.047
R41292 S.n13151 S.n13148 0.047
R41293 S.n11742 S.n11740 0.047
R41294 S.n12207 S.n12203 0.047
R41295 S.n22496 S.n22491 0.047
R41296 S.n22145 S.n22141 0.047
R41297 S.n21473 S.n21468 0.047
R41298 S.n21807 S.n21803 0.047
R41299 S.n20650 S.n20645 0.047
R41300 S.n20997 S.n20993 0.047
R41301 S.n20039 S.n20034 0.047
R41302 S.n19653 S.n19649 0.047
R41303 S.n19185 S.n19180 0.047
R41304 S.n18781 S.n18777 0.047
R41305 S.n18319 S.n18314 0.047
R41306 S.n17898 S.n17894 0.047
R41307 S.n17430 S.n17425 0.047
R41308 S.n16989 S.n16985 0.047
R41309 S.n16528 S.n16523 0.047
R41310 S.n16071 S.n16067 0.047
R41311 S.n15604 S.n15599 0.047
R41312 S.n15127 S.n15123 0.047
R41313 S.n14667 S.n14662 0.047
R41314 S.n14174 S.n14170 0.047
R41315 S.n13708 S.n13703 0.047
R41316 S.n13195 S.n13191 0.047
R41317 S.n12736 S.n12731 0.047
R41318 S.n12178 S.n12175 0.047
R41319 S.n10719 S.n10717 0.047
R41320 S.n11208 S.n11204 0.047
R41321 S.n22480 S.n22475 0.047
R41322 S.n22160 S.n22156 0.047
R41323 S.n21457 S.n21452 0.047
R41324 S.n21792 S.n21788 0.047
R41325 S.n20634 S.n20629 0.047
R41326 S.n20982 S.n20978 0.047
R41327 S.n20023 S.n20018 0.047
R41328 S.n19668 S.n19664 0.047
R41329 S.n19169 S.n19164 0.047
R41330 S.n18796 S.n18792 0.047
R41331 S.n18303 S.n18298 0.047
R41332 S.n17913 S.n17909 0.047
R41333 S.n17414 S.n17409 0.047
R41334 S.n17004 S.n17000 0.047
R41335 S.n16512 S.n16507 0.047
R41336 S.n16086 S.n16082 0.047
R41337 S.n15588 S.n15583 0.047
R41338 S.n15142 S.n15138 0.047
R41339 S.n14651 S.n14646 0.047
R41340 S.n14189 S.n14185 0.047
R41341 S.n13692 S.n13687 0.047
R41342 S.n13210 S.n13206 0.047
R41343 S.n12720 S.n12715 0.047
R41344 S.n12222 S.n12218 0.047
R41345 S.n11726 S.n11721 0.047
R41346 S.n11179 S.n11176 0.047
R41347 S.n9674 S.n9672 0.047
R41348 S.n10200 S.n10196 0.047
R41349 S.n22464 S.n22459 0.047
R41350 S.n22175 S.n22171 0.047
R41351 S.n21441 S.n21436 0.047
R41352 S.n21777 S.n21773 0.047
R41353 S.n20618 S.n20613 0.047
R41354 S.n20967 S.n20963 0.047
R41355 S.n20007 S.n20002 0.047
R41356 S.n19683 S.n19679 0.047
R41357 S.n19153 S.n19148 0.047
R41358 S.n18811 S.n18807 0.047
R41359 S.n18287 S.n18282 0.047
R41360 S.n17928 S.n17924 0.047
R41361 S.n17398 S.n17393 0.047
R41362 S.n17019 S.n17015 0.047
R41363 S.n16496 S.n16491 0.047
R41364 S.n16101 S.n16097 0.047
R41365 S.n15572 S.n15567 0.047
R41366 S.n15157 S.n15153 0.047
R41367 S.n14635 S.n14630 0.047
R41368 S.n14204 S.n14200 0.047
R41369 S.n13676 S.n13671 0.047
R41370 S.n13225 S.n13221 0.047
R41371 S.n12704 S.n12699 0.047
R41372 S.n12237 S.n12233 0.047
R41373 S.n11710 S.n11705 0.047
R41374 S.n11223 S.n11219 0.047
R41375 S.n10703 S.n10698 0.047
R41376 S.n10171 S.n10168 0.047
R41377 S.n8616 S.n8614 0.047
R41378 S.n9166 S.n9162 0.047
R41379 S.n22448 S.n22443 0.047
R41380 S.n22190 S.n22186 0.047
R41381 S.n21425 S.n21420 0.047
R41382 S.n21762 S.n21758 0.047
R41383 S.n20602 S.n20597 0.047
R41384 S.n20952 S.n20948 0.047
R41385 S.n19991 S.n19986 0.047
R41386 S.n19698 S.n19694 0.047
R41387 S.n19137 S.n19132 0.047
R41388 S.n18826 S.n18822 0.047
R41389 S.n18271 S.n18266 0.047
R41390 S.n17943 S.n17939 0.047
R41391 S.n17382 S.n17377 0.047
R41392 S.n17034 S.n17030 0.047
R41393 S.n16480 S.n16475 0.047
R41394 S.n16116 S.n16112 0.047
R41395 S.n15556 S.n15551 0.047
R41396 S.n15172 S.n15168 0.047
R41397 S.n14619 S.n14614 0.047
R41398 S.n14219 S.n14215 0.047
R41399 S.n13660 S.n13655 0.047
R41400 S.n13240 S.n13236 0.047
R41401 S.n12688 S.n12683 0.047
R41402 S.n12252 S.n12248 0.047
R41403 S.n11694 S.n11689 0.047
R41404 S.n11238 S.n11234 0.047
R41405 S.n10687 S.n10682 0.047
R41406 S.n10215 S.n10211 0.047
R41407 S.n9658 S.n9653 0.047
R41408 S.n9137 S.n9134 0.047
R41409 S.n7536 S.n7534 0.047
R41410 S.n8123 S.n8119 0.047
R41411 S.n22432 S.n22427 0.047
R41412 S.n22205 S.n22201 0.047
R41413 S.n21409 S.n21404 0.047
R41414 S.n21747 S.n21743 0.047
R41415 S.n20586 S.n20581 0.047
R41416 S.n20937 S.n20933 0.047
R41417 S.n19975 S.n19970 0.047
R41418 S.n19713 S.n19709 0.047
R41419 S.n19121 S.n19116 0.047
R41420 S.n18841 S.n18837 0.047
R41421 S.n18255 S.n18250 0.047
R41422 S.n17958 S.n17954 0.047
R41423 S.n17366 S.n17361 0.047
R41424 S.n17049 S.n17045 0.047
R41425 S.n16464 S.n16459 0.047
R41426 S.n16131 S.n16127 0.047
R41427 S.n15540 S.n15535 0.047
R41428 S.n15187 S.n15183 0.047
R41429 S.n14603 S.n14598 0.047
R41430 S.n14234 S.n14230 0.047
R41431 S.n13644 S.n13639 0.047
R41432 S.n13255 S.n13251 0.047
R41433 S.n12672 S.n12667 0.047
R41434 S.n12267 S.n12263 0.047
R41435 S.n11678 S.n11673 0.047
R41436 S.n11253 S.n11249 0.047
R41437 S.n10671 S.n10666 0.047
R41438 S.n10230 S.n10226 0.047
R41439 S.n9642 S.n9637 0.047
R41440 S.n9181 S.n9177 0.047
R41441 S.n8600 S.n8595 0.047
R41442 S.n8094 S.n8091 0.047
R41443 S.n6443 S.n6441 0.047
R41444 S.n7054 S.n7050 0.047
R41445 S.n22416 S.n22411 0.047
R41446 S.n22220 S.n22216 0.047
R41447 S.n21393 S.n21388 0.047
R41448 S.n21732 S.n21728 0.047
R41449 S.n20570 S.n20565 0.047
R41450 S.n20922 S.n20918 0.047
R41451 S.n19959 S.n19954 0.047
R41452 S.n19728 S.n19724 0.047
R41453 S.n19105 S.n19100 0.047
R41454 S.n18856 S.n18852 0.047
R41455 S.n18239 S.n18234 0.047
R41456 S.n17973 S.n17969 0.047
R41457 S.n17350 S.n17345 0.047
R41458 S.n17064 S.n17060 0.047
R41459 S.n16448 S.n16443 0.047
R41460 S.n16146 S.n16142 0.047
R41461 S.n15524 S.n15519 0.047
R41462 S.n15202 S.n15198 0.047
R41463 S.n14587 S.n14582 0.047
R41464 S.n14249 S.n14245 0.047
R41465 S.n13628 S.n13623 0.047
R41466 S.n13270 S.n13266 0.047
R41467 S.n12656 S.n12651 0.047
R41468 S.n12282 S.n12278 0.047
R41469 S.n11662 S.n11657 0.047
R41470 S.n11268 S.n11264 0.047
R41471 S.n10655 S.n10650 0.047
R41472 S.n10245 S.n10241 0.047
R41473 S.n9626 S.n9621 0.047
R41474 S.n9196 S.n9192 0.047
R41475 S.n8584 S.n8579 0.047
R41476 S.n8138 S.n8134 0.047
R41477 S.n7520 S.n7515 0.047
R41478 S.n7025 S.n7022 0.047
R41479 S.n5327 S.n5325 0.047
R41480 S.n5976 S.n5972 0.047
R41481 S.n22400 S.n22395 0.047
R41482 S.n22235 S.n22231 0.047
R41483 S.n21377 S.n21372 0.047
R41484 S.n21717 S.n21713 0.047
R41485 S.n20554 S.n20549 0.047
R41486 S.n20907 S.n20903 0.047
R41487 S.n19943 S.n19938 0.047
R41488 S.n19743 S.n19739 0.047
R41489 S.n19089 S.n19084 0.047
R41490 S.n18871 S.n18867 0.047
R41491 S.n18223 S.n18218 0.047
R41492 S.n17988 S.n17984 0.047
R41493 S.n17334 S.n17329 0.047
R41494 S.n17079 S.n17075 0.047
R41495 S.n16432 S.n16427 0.047
R41496 S.n16161 S.n16157 0.047
R41497 S.n15508 S.n15503 0.047
R41498 S.n15217 S.n15213 0.047
R41499 S.n14571 S.n14566 0.047
R41500 S.n14264 S.n14260 0.047
R41501 S.n13612 S.n13607 0.047
R41502 S.n13285 S.n13281 0.047
R41503 S.n12640 S.n12635 0.047
R41504 S.n12297 S.n12293 0.047
R41505 S.n11646 S.n11641 0.047
R41506 S.n11283 S.n11279 0.047
R41507 S.n10639 S.n10634 0.047
R41508 S.n10260 S.n10256 0.047
R41509 S.n9610 S.n9605 0.047
R41510 S.n9211 S.n9207 0.047
R41511 S.n8568 S.n8563 0.047
R41512 S.n8153 S.n8149 0.047
R41513 S.n7504 S.n7499 0.047
R41514 S.n7069 S.n7065 0.047
R41515 S.n6427 S.n6422 0.047
R41516 S.n5947 S.n5944 0.047
R41517 S.n4198 S.n4196 0.047
R41518 S.n4871 S.n4867 0.047
R41519 S.n22384 S.n22379 0.047
R41520 S.n22250 S.n22246 0.047
R41521 S.n21361 S.n21356 0.047
R41522 S.n21702 S.n21698 0.047
R41523 S.n20538 S.n20533 0.047
R41524 S.n20892 S.n20888 0.047
R41525 S.n19927 S.n19922 0.047
R41526 S.n19758 S.n19754 0.047
R41527 S.n19073 S.n19068 0.047
R41528 S.n18886 S.n18882 0.047
R41529 S.n18207 S.n18202 0.047
R41530 S.n18003 S.n17999 0.047
R41531 S.n17318 S.n17313 0.047
R41532 S.n17094 S.n17090 0.047
R41533 S.n16416 S.n16411 0.047
R41534 S.n16176 S.n16172 0.047
R41535 S.n15492 S.n15487 0.047
R41536 S.n15232 S.n15228 0.047
R41537 S.n14555 S.n14550 0.047
R41538 S.n14279 S.n14275 0.047
R41539 S.n13596 S.n13591 0.047
R41540 S.n13300 S.n13296 0.047
R41541 S.n12624 S.n12619 0.047
R41542 S.n12312 S.n12308 0.047
R41543 S.n11630 S.n11625 0.047
R41544 S.n11298 S.n11294 0.047
R41545 S.n10623 S.n10618 0.047
R41546 S.n10275 S.n10271 0.047
R41547 S.n9594 S.n9589 0.047
R41548 S.n9229 S.n9225 0.047
R41549 S.n8552 S.n8547 0.047
R41550 S.n8168 S.n8164 0.047
R41551 S.n7488 S.n7483 0.047
R41552 S.n7084 S.n7080 0.047
R41553 S.n6411 S.n6406 0.047
R41554 S.n5991 S.n5987 0.047
R41555 S.n5311 S.n5306 0.047
R41556 S.n4841 S.n4838 0.047
R41557 S.n3057 S.n3055 0.047
R41558 S.n3759 S.n3754 0.047
R41559 S.n22672 S.n22269 0.047
R41560 S.n22675 S.n22261 0.047
R41561 S.n21685 S.n21675 0.047
R41562 S.n21687 S.n21667 0.047
R41563 S.n20522 S.n20518 0.047
R41564 S.n20877 S.n20872 0.047
R41565 S.n19911 S.n19907 0.047
R41566 S.n19774 S.n19769 0.047
R41567 S.n19057 S.n19053 0.047
R41568 S.n18902 S.n18897 0.047
R41569 S.n18191 S.n18187 0.047
R41570 S.n18019 S.n18014 0.047
R41571 S.n17302 S.n17298 0.047
R41572 S.n17110 S.n17105 0.047
R41573 S.n16400 S.n16396 0.047
R41574 S.n16192 S.n16187 0.047
R41575 S.n15476 S.n15472 0.047
R41576 S.n15248 S.n15243 0.047
R41577 S.n14539 S.n14535 0.047
R41578 S.n14295 S.n14290 0.047
R41579 S.n13580 S.n13576 0.047
R41580 S.n13316 S.n13311 0.047
R41581 S.n12608 S.n12604 0.047
R41582 S.n12328 S.n12323 0.047
R41583 S.n11614 S.n11610 0.047
R41584 S.n11314 S.n11309 0.047
R41585 S.n10607 S.n10603 0.047
R41586 S.n10291 S.n10286 0.047
R41587 S.n9578 S.n9574 0.047
R41588 S.n9242 S.n9237 0.047
R41589 S.n8536 S.n8532 0.047
R41590 S.n8184 S.n8179 0.047
R41591 S.n7472 S.n7468 0.047
R41592 S.n7100 S.n7095 0.047
R41593 S.n6395 S.n6391 0.047
R41594 S.n6007 S.n6002 0.047
R41595 S.n5295 S.n5291 0.047
R41596 S.n4887 S.n4882 0.047
R41597 S.n4182 S.n4178 0.047
R41598 S.n3728 S.n3725 0.047
R41599 S.n1899 S.n1897 0.047
R41600 S.n2628 S.n2623 0.047
R41601 S.n22368 S.n22362 0.047
R41602 S.n22694 S.n22686 0.047
R41603 S.n21654 S.n21280 0.047
R41604 S.n21656 S.n21272 0.047
R41605 S.n20507 S.n20503 0.047
R41606 S.n20861 S.n20856 0.047
R41607 S.n19896 S.n19892 0.047
R41608 S.n19790 S.n19785 0.047
R41609 S.n19042 S.n19038 0.047
R41610 S.n18918 S.n18913 0.047
R41611 S.n18176 S.n18172 0.047
R41612 S.n18035 S.n18030 0.047
R41613 S.n17287 S.n17283 0.047
R41614 S.n17126 S.n17121 0.047
R41615 S.n16385 S.n16381 0.047
R41616 S.n16208 S.n16203 0.047
R41617 S.n15461 S.n15457 0.047
R41618 S.n15264 S.n15259 0.047
R41619 S.n14524 S.n14520 0.047
R41620 S.n14311 S.n14306 0.047
R41621 S.n13565 S.n13561 0.047
R41622 S.n13332 S.n13327 0.047
R41623 S.n12593 S.n12589 0.047
R41624 S.n12344 S.n12339 0.047
R41625 S.n11599 S.n11595 0.047
R41626 S.n11330 S.n11325 0.047
R41627 S.n10592 S.n10588 0.047
R41628 S.n10307 S.n10302 0.047
R41629 S.n9563 S.n9559 0.047
R41630 S.n9258 S.n9253 0.047
R41631 S.n8521 S.n8517 0.047
R41632 S.n8200 S.n8195 0.047
R41633 S.n7457 S.n7453 0.047
R41634 S.n7116 S.n7111 0.047
R41635 S.n6380 S.n6376 0.047
R41636 S.n6023 S.n6018 0.047
R41637 S.n5280 S.n5276 0.047
R41638 S.n4903 S.n4898 0.047
R41639 S.n4167 S.n4163 0.047
R41640 S.n3775 S.n3770 0.047
R41641 S.n3041 S.n3037 0.047
R41642 S.n2597 S.n2594 0.047
R41643 S.n914 S.n899 0.047
R41644 S.n1985 S.n1975 0.047
R41645 S.n22741 S.n22726 0.047
R41646 S.n21314 S.n21306 0.047
R41647 S.n21217 S.n21205 0.047
R41648 S.n20491 S.n20483 0.047
R41649 S.n20398 S.n20386 0.047
R41650 S.n19880 S.n19872 0.047
R41651 S.n20271 S.n20259 0.047
R41652 S.n19026 S.n19018 0.047
R41653 S.n19403 S.n19391 0.047
R41654 S.n18160 S.n18152 0.047
R41655 S.n18516 S.n18504 0.047
R41656 S.n17271 S.n17263 0.047
R41657 S.n17616 S.n17604 0.047
R41658 S.n16369 S.n16361 0.047
R41659 S.n16693 S.n16681 0.047
R41660 S.n15445 S.n15437 0.047
R41661 S.n15758 S.n15746 0.047
R41662 S.n14508 S.n14500 0.047
R41663 S.n14800 S.n14788 0.047
R41664 S.n13549 S.n13541 0.047
R41665 S.n13830 S.n13818 0.047
R41666 S.n12577 S.n12569 0.047
R41667 S.n12837 S.n12825 0.047
R41668 S.n11583 S.n11575 0.047
R41669 S.n11832 S.n11820 0.047
R41670 S.n10576 S.n10568 0.047
R41671 S.n10804 S.n10792 0.047
R41672 S.n9547 S.n9539 0.047
R41673 S.n9764 S.n9752 0.047
R41674 S.n8505 S.n8497 0.047
R41675 S.n8701 S.n8689 0.047
R41676 S.n7441 S.n7433 0.047
R41677 S.n7626 S.n7614 0.047
R41678 S.n6364 S.n6356 0.047
R41679 S.n6528 S.n6516 0.047
R41680 S.n5264 S.n5256 0.047
R41681 S.n5417 S.n5405 0.047
R41682 S.n4151 S.n4143 0.047
R41683 S.n4283 S.n4271 0.047
R41684 S.n3025 S.n3017 0.047
R41685 S.n3146 S.n3135 0.047
R41686 S.n1865 S.n1856 0.047
R41687 S.n890 S.n883 0.047
R41688 S.n806 S.n801 0.047
R41689 S.n974 S.n954 0.047
R41690 S.n22351 S.n22349 0.047
R41691 S.n22713 S.n22711 0.047
R41692 S.n21345 S.n21343 0.047
R41693 S.n21261 S.n21259 0.047
R41694 S.n20835 S.n20833 0.047
R41695 S.n20845 S.n20843 0.047
R41696 S.n20200 S.n20198 0.047
R41697 S.n20210 S.n20208 0.047
R41698 S.n19330 S.n19328 0.047
R41699 S.n19340 S.n19338 0.047
R41700 S.n18448 S.n18446 0.047
R41701 S.n18458 S.n18456 0.047
R41702 S.n17543 S.n17541 0.047
R41703 S.n17553 S.n17551 0.047
R41704 S.n16625 S.n16623 0.047
R41705 S.n16635 S.n16633 0.047
R41706 S.n15685 S.n15683 0.047
R41707 S.n15695 S.n15693 0.047
R41708 S.n14732 S.n14730 0.047
R41709 S.n14742 S.n14740 0.047
R41710 S.n13757 S.n13755 0.047
R41711 S.n13767 S.n13765 0.047
R41712 S.n12769 S.n12767 0.047
R41713 S.n12779 S.n12777 0.047
R41714 S.n11759 S.n11757 0.047
R41715 S.n11769 S.n11767 0.047
R41716 S.n10736 S.n10734 0.047
R41717 S.n10746 S.n10744 0.047
R41718 S.n9691 S.n9689 0.047
R41719 S.n9701 S.n9699 0.047
R41720 S.n8633 S.n8631 0.047
R41721 S.n8643 S.n8641 0.047
R41722 S.n7553 S.n7551 0.047
R41723 S.n7563 S.n7561 0.047
R41724 S.n6460 S.n6458 0.047
R41725 S.n6470 S.n6468 0.047
R41726 S.n5344 S.n5342 0.047
R41727 S.n5354 S.n5352 0.047
R41728 S.n4215 S.n4213 0.047
R41729 S.n4225 S.n4223 0.047
R41730 S.n3074 S.n3072 0.047
R41731 S.n3084 S.n3082 0.047
R41732 S.n1882 S.n1880 0.047
R41733 S.n1931 S.n1925 0.047
R41734 S.n406 S.n404 0.047
R41735 S.n2137 S.n2127 0.047
R41736 S.n18483 S.n18469 0.047
R41737 S.n17169 S.n17161 0.047
R41738 S.n17765 S.n17753 0.047
R41739 S.n16269 S.n16261 0.047
R41740 S.n16838 S.n16826 0.047
R41741 S.n15345 S.n15337 0.047
R41742 S.n15903 S.n15891 0.047
R41743 S.n14408 S.n14400 0.047
R41744 S.n14945 S.n14933 0.047
R41745 S.n13449 S.n13441 0.047
R41746 S.n13975 S.n13963 0.047
R41747 S.n12477 S.n12469 0.047
R41748 S.n12982 S.n12970 0.047
R41749 S.n11483 S.n11475 0.047
R41750 S.n11977 S.n11965 0.047
R41751 S.n10476 S.n10468 0.047
R41752 S.n10949 S.n10937 0.047
R41753 S.n9447 S.n9439 0.047
R41754 S.n9909 S.n9897 0.047
R41755 S.n8405 S.n8397 0.047
R41756 S.n8846 S.n8834 0.047
R41757 S.n7341 S.n7333 0.047
R41758 S.n7771 S.n7759 0.047
R41759 S.n6264 S.n6256 0.047
R41760 S.n6673 S.n6661 0.047
R41761 S.n5164 S.n5156 0.047
R41762 S.n5563 S.n5551 0.047
R41763 S.n4052 S.n4044 0.047
R41764 S.n4428 S.n4416 0.047
R41765 S.n2925 S.n2917 0.047
R41766 S.n3290 S.n3279 0.047
R41767 S.n1757 S.n1748 0.047
R41768 S.n24 S.n22 0.047
R41769 S.n19370 S.n19361 0.047
R41770 S.n18077 S.n18075 0.047
R41771 S.n18633 S.n18622 0.047
R41772 S.n17188 S.n17186 0.047
R41773 S.n17733 S.n17722 0.047
R41774 S.n16286 S.n16284 0.047
R41775 S.n16806 S.n16795 0.047
R41776 S.n15362 S.n15360 0.047
R41777 S.n15871 S.n15860 0.047
R41778 S.n14425 S.n14423 0.047
R41779 S.n14913 S.n14902 0.047
R41780 S.n13466 S.n13464 0.047
R41781 S.n13943 S.n13932 0.047
R41782 S.n12494 S.n12492 0.047
R41783 S.n12950 S.n12939 0.047
R41784 S.n11500 S.n11498 0.047
R41785 S.n11945 S.n11934 0.047
R41786 S.n10493 S.n10491 0.047
R41787 S.n10917 S.n10906 0.047
R41788 S.n9464 S.n9462 0.047
R41789 S.n9877 S.n9866 0.047
R41790 S.n8422 S.n8420 0.047
R41791 S.n8814 S.n8803 0.047
R41792 S.n7358 S.n7356 0.047
R41793 S.n7739 S.n7728 0.047
R41794 S.n6281 S.n6279 0.047
R41795 S.n6641 S.n6630 0.047
R41796 S.n5181 S.n5179 0.047
R41797 S.n5531 S.n5520 0.047
R41798 S.n4069 S.n4067 0.047
R41799 S.n4396 S.n4385 0.047
R41800 S.n2942 S.n2940 0.047
R41801 S.n3259 S.n3248 0.047
R41802 S.n1776 S.n1772 0.047
R41803 S.n1799 S.n1794 0.047
R41804 S.n2079 S.n2064 0.047
R41805 S.n823 S.n821 0.047
R41806 S.n838 S.n832 0.047
R41807 S.n3230 S.n3219 0.047
R41808 S.n4367 S.n4355 0.047
R41809 S.n5502 S.n5490 0.047
R41810 S.n6612 S.n6600 0.047
R41811 S.n7710 S.n7698 0.047
R41812 S.n8785 S.n8773 0.047
R41813 S.n9848 S.n9836 0.047
R41814 S.n10888 S.n10876 0.047
R41815 S.n11916 S.n11904 0.047
R41816 S.n12921 S.n12909 0.047
R41817 S.n13914 S.n13902 0.047
R41818 S.n14884 S.n14872 0.047
R41819 S.n15842 S.n15830 0.047
R41820 S.n16777 S.n16765 0.047
R41821 S.n17700 S.n17688 0.047
R41822 S.n18600 S.n18588 0.047
R41823 S.n19490 S.n19478 0.047
R41824 S.n20238 S.n20224 0.047
R41825 S.n18961 S.n18953 0.047
R41826 S.n18096 S.n18088 0.047
R41827 S.n17207 S.n17199 0.047
R41828 S.n16305 S.n16297 0.047
R41829 S.n15381 S.n15373 0.047
R41830 S.n14444 S.n14436 0.047
R41831 S.n13485 S.n13477 0.047
R41832 S.n12513 S.n12505 0.047
R41833 S.n11519 S.n11511 0.047
R41834 S.n10512 S.n10504 0.047
R41835 S.n9483 S.n9475 0.047
R41836 S.n8441 S.n8433 0.047
R41837 S.n7377 S.n7369 0.047
R41838 S.n6300 S.n6292 0.047
R41839 S.n5200 S.n5192 0.047
R41840 S.n4088 S.n4080 0.047
R41841 S.n2961 S.n2953 0.047
R41842 S.n2045 S.n2036 0.047
R41843 S.n767 S.n757 0.047
R41844 S.n1337 S.n1334 0.047
R41845 S.n20424 S.n20416 0.047
R41846 S.n19839 S.n19833 0.047
R41847 S.n20330 S.n20312 0.047
R41848 S.n18987 S.n18981 0.047
R41849 S.n19458 S.n19440 0.047
R41850 S.n18121 S.n18116 0.047
R41851 S.n18568 S.n18553 0.047
R41852 S.n17232 S.n17227 0.047
R41853 S.n17668 S.n17653 0.047
R41854 S.n16330 S.n16325 0.047
R41855 S.n16745 S.n16730 0.047
R41856 S.n15406 S.n15401 0.047
R41857 S.n15810 S.n15795 0.047
R41858 S.n14469 S.n14464 0.047
R41859 S.n14852 S.n14837 0.047
R41860 S.n13510 S.n13505 0.047
R41861 S.n13882 S.n13867 0.047
R41862 S.n12538 S.n12533 0.047
R41863 S.n12889 S.n12874 0.047
R41864 S.n11544 S.n11539 0.047
R41865 S.n11884 S.n11869 0.047
R41866 S.n10537 S.n10532 0.047
R41867 S.n10856 S.n10841 0.047
R41868 S.n9508 S.n9503 0.047
R41869 S.n9816 S.n9801 0.047
R41870 S.n8466 S.n8461 0.047
R41871 S.n8753 S.n8738 0.047
R41872 S.n7402 S.n7397 0.047
R41873 S.n7678 S.n7663 0.047
R41874 S.n6325 S.n6320 0.047
R41875 S.n6580 S.n6565 0.047
R41876 S.n5225 S.n5220 0.047
R41877 S.n5470 S.n5455 0.047
R41878 S.n4113 S.n4108 0.047
R41879 S.n4335 S.n4320 0.047
R41880 S.n2986 S.n2981 0.047
R41881 S.n3198 S.n3183 0.047
R41882 S.n1823 S.n1818 0.047
R41883 S.n2012 S.n2003 0.047
R41884 S.n786 S.n781 0.047
R41885 S.n1845 S.n1839 0.047
R41886 S.n3166 S.n3164 0.047
R41887 S.n3006 S.n3001 0.047
R41888 S.n4303 S.n4301 0.047
R41889 S.n4132 S.n4128 0.047
R41890 S.n5438 S.n5435 0.047
R41891 S.n5245 S.n5240 0.047
R41892 S.n6548 S.n6546 0.047
R41893 S.n6345 S.n6340 0.047
R41894 S.n7646 S.n7644 0.047
R41895 S.n7422 S.n7417 0.047
R41896 S.n8721 S.n8719 0.047
R41897 S.n8486 S.n8481 0.047
R41898 S.n9784 S.n9782 0.047
R41899 S.n9528 S.n9523 0.047
R41900 S.n10824 S.n10822 0.047
R41901 S.n10557 S.n10552 0.047
R41902 S.n11852 S.n11850 0.047
R41903 S.n11564 S.n11559 0.047
R41904 S.n12857 S.n12855 0.047
R41905 S.n12558 S.n12553 0.047
R41906 S.n13850 S.n13848 0.047
R41907 S.n13530 S.n13525 0.047
R41908 S.n14820 S.n14818 0.047
R41909 S.n14489 S.n14484 0.047
R41910 S.n15778 S.n15776 0.047
R41911 S.n15426 S.n15421 0.047
R41912 S.n16713 S.n16711 0.047
R41913 S.n16350 S.n16345 0.047
R41914 S.n17636 S.n17634 0.047
R41915 S.n17252 S.n17247 0.047
R41916 S.n18536 S.n18534 0.047
R41917 S.n18141 S.n18136 0.047
R41918 S.n19423 S.n19421 0.047
R41919 S.n19007 S.n19002 0.047
R41920 S.n20295 S.n20293 0.047
R41921 S.n19861 S.n19856 0.047
R41922 S.n20366 S.n20364 0.047
R41923 S.n20472 S.n20467 0.047
R41924 S.n21242 S.n21240 0.047
R41925 S.n864 S.n856 0.047
R41926 S.n2107 S.n2097 0.047
R41927 S.n743 S.n741 0.047
R41928 S.n726 S.n724 0.047
R41929 S.n374 S.n372 0.047
R41930 S.n2196 S.n2186 0.047
R41931 S.n16660 S.n16646 0.047
R41932 S.n15307 S.n15299 0.047
R41933 S.n15968 S.n15956 0.047
R41934 S.n14372 S.n14364 0.047
R41935 S.n15006 S.n14994 0.047
R41936 S.n13413 S.n13405 0.047
R41937 S.n14036 S.n14024 0.047
R41938 S.n12441 S.n12433 0.047
R41939 S.n13043 S.n13031 0.047
R41940 S.n11447 S.n11439 0.047
R41941 S.n12038 S.n12026 0.047
R41942 S.n10440 S.n10432 0.047
R41943 S.n11010 S.n10998 0.047
R41944 S.n9411 S.n9403 0.047
R41945 S.n9970 S.n9958 0.047
R41946 S.n8369 S.n8361 0.047
R41947 S.n8907 S.n8895 0.047
R41948 S.n7305 S.n7297 0.047
R41949 S.n7832 S.n7820 0.047
R41950 S.n6228 S.n6220 0.047
R41951 S.n6734 S.n6722 0.047
R41952 S.n5128 S.n5120 0.047
R41953 S.n5624 S.n5612 0.047
R41954 S.n4016 S.n4008 0.047
R41955 S.n4489 S.n4477 0.047
R41956 S.n2889 S.n2881 0.047
R41957 S.n3350 S.n3339 0.047
R41958 S.n1720 S.n1711 0.047
R41959 S.n71 S.n69 0.047
R41960 S.n17583 S.n17574 0.047
R41961 S.n16250 S.n16248 0.047
R41962 S.n16871 S.n16860 0.047
R41963 S.n15326 S.n15324 0.047
R41964 S.n15936 S.n15925 0.047
R41965 S.n14389 S.n14387 0.047
R41966 S.n14974 S.n14963 0.047
R41967 S.n13430 S.n13428 0.047
R41968 S.n14004 S.n13993 0.047
R41969 S.n12458 S.n12456 0.047
R41970 S.n13011 S.n13000 0.047
R41971 S.n11464 S.n11462 0.047
R41972 S.n12006 S.n11995 0.047
R41973 S.n10457 S.n10455 0.047
R41974 S.n10978 S.n10967 0.047
R41975 S.n9428 S.n9426 0.047
R41976 S.n9938 S.n9927 0.047
R41977 S.n8386 S.n8384 0.047
R41978 S.n8875 S.n8864 0.047
R41979 S.n7322 S.n7320 0.047
R41980 S.n7800 S.n7789 0.047
R41981 S.n6245 S.n6243 0.047
R41982 S.n6702 S.n6691 0.047
R41983 S.n5145 S.n5143 0.047
R41984 S.n5592 S.n5581 0.047
R41985 S.n4033 S.n4031 0.047
R41986 S.n4457 S.n4446 0.047
R41987 S.n2906 S.n2904 0.047
R41988 S.n3319 S.n3308 0.047
R41989 S.n1737 S.n1735 0.047
R41990 S.n2166 S.n2155 0.047
R41991 S.n708 S.n706 0.047
R41992 S.n691 S.n689 0.047
R41993 S.n342 S.n340 0.047
R41994 S.n2255 S.n2245 0.047
R41995 S.n14767 S.n14753 0.047
R41996 S.n13375 S.n13367 0.047
R41997 S.n14101 S.n14089 0.047
R41998 S.n12405 S.n12397 0.047
R41999 S.n13104 S.n13092 0.047
R42000 S.n11411 S.n11403 0.047
R42001 S.n12099 S.n12087 0.047
R42002 S.n10404 S.n10396 0.047
R42003 S.n11071 S.n11059 0.047
R42004 S.n9375 S.n9367 0.047
R42005 S.n10031 S.n10019 0.047
R42006 S.n8333 S.n8325 0.047
R42007 S.n8968 S.n8956 0.047
R42008 S.n7269 S.n7261 0.047
R42009 S.n7893 S.n7881 0.047
R42010 S.n6192 S.n6184 0.047
R42011 S.n6795 S.n6783 0.047
R42012 S.n5092 S.n5084 0.047
R42013 S.n5685 S.n5673 0.047
R42014 S.n3980 S.n3972 0.047
R42015 S.n4550 S.n4538 0.047
R42016 S.n2853 S.n2845 0.047
R42017 S.n3410 S.n3399 0.047
R42018 S.n1683 S.n1674 0.047
R42019 S.n103 S.n101 0.047
R42020 S.n15725 S.n15716 0.047
R42021 S.n14353 S.n14351 0.047
R42022 S.n15039 S.n15028 0.047
R42023 S.n13394 S.n13392 0.047
R42024 S.n14069 S.n14058 0.047
R42025 S.n12422 S.n12420 0.047
R42026 S.n13072 S.n13061 0.047
R42027 S.n11428 S.n11426 0.047
R42028 S.n12067 S.n12056 0.047
R42029 S.n10421 S.n10419 0.047
R42030 S.n11039 S.n11028 0.047
R42031 S.n9392 S.n9390 0.047
R42032 S.n9999 S.n9988 0.047
R42033 S.n8350 S.n8348 0.047
R42034 S.n8936 S.n8925 0.047
R42035 S.n7286 S.n7284 0.047
R42036 S.n7861 S.n7850 0.047
R42037 S.n6209 S.n6207 0.047
R42038 S.n6763 S.n6752 0.047
R42039 S.n5109 S.n5107 0.047
R42040 S.n5653 S.n5642 0.047
R42041 S.n3997 S.n3995 0.047
R42042 S.n4518 S.n4507 0.047
R42043 S.n2870 S.n2868 0.047
R42044 S.n3379 S.n3368 0.047
R42045 S.n1700 S.n1698 0.047
R42046 S.n2225 S.n2214 0.047
R42047 S.n673 S.n671 0.047
R42048 S.n656 S.n654 0.047
R42049 S.n310 S.n308 0.047
R42050 S.n2314 S.n2304 0.047
R42051 S.n12804 S.n12790 0.047
R42052 S.n11373 S.n11365 0.047
R42053 S.n12164 S.n12152 0.047
R42054 S.n10368 S.n10360 0.047
R42055 S.n11132 S.n11120 0.047
R42056 S.n9339 S.n9331 0.047
R42057 S.n10092 S.n10080 0.047
R42058 S.n8297 S.n8289 0.047
R42059 S.n9029 S.n9017 0.047
R42060 S.n7233 S.n7225 0.047
R42061 S.n7954 S.n7942 0.047
R42062 S.n6156 S.n6148 0.047
R42063 S.n6856 S.n6844 0.047
R42064 S.n5056 S.n5048 0.047
R42065 S.n5746 S.n5734 0.047
R42066 S.n3944 S.n3936 0.047
R42067 S.n4611 S.n4599 0.047
R42068 S.n2817 S.n2809 0.047
R42069 S.n3470 S.n3459 0.047
R42070 S.n1646 S.n1637 0.047
R42071 S.n990 S.n988 0.047
R42072 S.n13797 S.n13788 0.047
R42073 S.n12386 S.n12384 0.047
R42074 S.n13137 S.n13126 0.047
R42075 S.n11392 S.n11390 0.047
R42076 S.n12132 S.n12121 0.047
R42077 S.n10385 S.n10383 0.047
R42078 S.n11100 S.n11089 0.047
R42079 S.n9356 S.n9354 0.047
R42080 S.n10060 S.n10049 0.047
R42081 S.n8314 S.n8312 0.047
R42082 S.n8997 S.n8986 0.047
R42083 S.n7250 S.n7248 0.047
R42084 S.n7922 S.n7911 0.047
R42085 S.n6173 S.n6171 0.047
R42086 S.n6824 S.n6813 0.047
R42087 S.n5073 S.n5071 0.047
R42088 S.n5714 S.n5703 0.047
R42089 S.n3961 S.n3959 0.047
R42090 S.n4579 S.n4568 0.047
R42091 S.n2834 S.n2832 0.047
R42092 S.n3439 S.n3428 0.047
R42093 S.n1663 S.n1661 0.047
R42094 S.n2284 S.n2273 0.047
R42095 S.n638 S.n636 0.047
R42096 S.n621 S.n619 0.047
R42097 S.n278 S.n276 0.047
R42098 S.n2373 S.n2363 0.047
R42099 S.n10771 S.n10757 0.047
R42100 S.n9301 S.n9293 0.047
R42101 S.n10157 S.n10145 0.047
R42102 S.n8261 S.n8253 0.047
R42103 S.n9090 S.n9078 0.047
R42104 S.n7197 S.n7189 0.047
R42105 S.n8015 S.n8003 0.047
R42106 S.n6120 S.n6112 0.047
R42107 S.n6917 S.n6905 0.047
R42108 S.n5020 S.n5012 0.047
R42109 S.n5807 S.n5795 0.047
R42110 S.n3908 S.n3900 0.047
R42111 S.n4672 S.n4660 0.047
R42112 S.n2781 S.n2773 0.047
R42113 S.n3530 S.n3519 0.047
R42114 S.n1609 S.n1600 0.047
R42115 S.n1022 S.n1020 0.047
R42116 S.n11799 S.n11790 0.047
R42117 S.n10349 S.n10347 0.047
R42118 S.n11165 S.n11154 0.047
R42119 S.n9320 S.n9318 0.047
R42120 S.n10125 S.n10114 0.047
R42121 S.n8278 S.n8276 0.047
R42122 S.n9058 S.n9047 0.047
R42123 S.n7214 S.n7212 0.047
R42124 S.n7983 S.n7972 0.047
R42125 S.n6137 S.n6135 0.047
R42126 S.n6885 S.n6874 0.047
R42127 S.n5037 S.n5035 0.047
R42128 S.n5775 S.n5764 0.047
R42129 S.n3925 S.n3923 0.047
R42130 S.n4640 S.n4629 0.047
R42131 S.n2798 S.n2796 0.047
R42132 S.n3499 S.n3488 0.047
R42133 S.n1626 S.n1624 0.047
R42134 S.n2343 S.n2332 0.047
R42135 S.n603 S.n601 0.047
R42136 S.n586 S.n584 0.047
R42137 S.n249 S.n247 0.047
R42138 S.n2432 S.n2422 0.047
R42139 S.n8668 S.n8654 0.047
R42140 S.n7159 S.n7151 0.047
R42141 S.n8080 S.n8068 0.047
R42142 S.n6084 S.n6076 0.047
R42143 S.n6978 S.n6966 0.047
R42144 S.n4984 S.n4976 0.047
R42145 S.n5868 S.n5856 0.047
R42146 S.n3872 S.n3864 0.047
R42147 S.n4733 S.n4721 0.047
R42148 S.n2745 S.n2737 0.047
R42149 S.n3590 S.n3579 0.047
R42150 S.n1572 S.n1563 0.047
R42151 S.n1054 S.n1052 0.047
R42152 S.n9731 S.n9722 0.047
R42153 S.n8242 S.n8240 0.047
R42154 S.n9123 S.n9112 0.047
R42155 S.n7178 S.n7176 0.047
R42156 S.n8048 S.n8037 0.047
R42157 S.n6101 S.n6099 0.047
R42158 S.n6946 S.n6935 0.047
R42159 S.n5001 S.n4999 0.047
R42160 S.n5836 S.n5825 0.047
R42161 S.n3889 S.n3887 0.047
R42162 S.n4701 S.n4690 0.047
R42163 S.n2762 S.n2760 0.047
R42164 S.n3559 S.n3548 0.047
R42165 S.n1589 S.n1587 0.047
R42166 S.n2402 S.n2391 0.047
R42167 S.n568 S.n566 0.047
R42168 S.n551 S.n549 0.047
R42169 S.n214 S.n212 0.047
R42170 S.n2491 S.n2481 0.047
R42171 S.n6495 S.n6481 0.047
R42172 S.n4946 S.n4938 0.047
R42173 S.n5933 S.n5921 0.047
R42174 S.n3836 S.n3828 0.047
R42175 S.n4794 S.n4782 0.047
R42176 S.n2709 S.n2701 0.047
R42177 S.n3650 S.n3639 0.047
R42178 S.n1535 S.n1526 0.047
R42179 S.n1086 S.n1084 0.047
R42180 S.n7593 S.n7584 0.047
R42181 S.n6065 S.n6063 0.047
R42182 S.n7011 S.n7000 0.047
R42183 S.n4965 S.n4963 0.047
R42184 S.n5901 S.n5890 0.047
R42185 S.n3853 S.n3851 0.047
R42186 S.n4762 S.n4751 0.047
R42187 S.n2726 S.n2724 0.047
R42188 S.n3619 S.n3608 0.047
R42189 S.n1552 S.n1550 0.047
R42190 S.n2461 S.n2450 0.047
R42191 S.n533 S.n531 0.047
R42192 S.n516 S.n514 0.047
R42193 S.n182 S.n180 0.047
R42194 S.n2550 S.n2540 0.047
R42195 S.n4250 S.n4236 0.047
R42196 S.n2671 S.n2663 0.047
R42197 S.n3714 S.n3703 0.047
R42198 S.n1498 S.n1489 0.047
R42199 S.n1118 S.n1116 0.047
R42200 S.n5384 S.n5375 0.047
R42201 S.n3817 S.n3815 0.047
R42202 S.n4827 S.n4816 0.047
R42203 S.n2690 S.n2688 0.047
R42204 S.n3683 S.n3672 0.047
R42205 S.n1515 S.n1513 0.047
R42206 S.n2520 S.n2509 0.047
R42207 S.n498 S.n496 0.047
R42208 S.n481 S.n479 0.047
R42209 S.n150 S.n148 0.047
R42210 S.n1954 S.n1942 0.047
R42211 S.n1156 S.n1154 0.047
R42212 S.n3114 S.n3105 0.047
R42213 S.n1478 S.n1476 0.047
R42214 S.n2583 S.n2572 0.047
R42215 S.n463 S.n461 0.047
R42216 S.n447 S.n445 0.047
R42217 S.n942 S.n935 0.047
R42218 S.n21980 S.n21975 0.047
R42219 S.n22765 S.n22763 0.047
R42220 S.n21328 S.n21326 0.047
R42221 S.n22307 S.n22303 0.047
R42222 S.n1365 S.n1364 0.046
R42223 S.t158 S.n1306 0.046
R42224 S.t158 S.n1296 0.046
R42225 S.t158 S.n1284 0.046
R42226 S.t158 S.n1272 0.046
R42227 S.t158 S.n1259 0.046
R42228 S.t158 S.n1246 0.046
R42229 S.t158 S.n1233 0.046
R42230 S.t158 S.n1220 0.046
R42231 S.t158 S.n1207 0.046
R42232 S.t158 S.n1194 0.046
R42233 S.n21961 S.n21960 0.046
R42234 S.n1313 S.n1311 0.045
R42235 S.n22999 S.n22998 0.045
R42236 S.n885 S.n884 0.045
R42237 S.n1321 S.n1320 0.045
R42238 S.n2027 S.n2019 0.045
R42239 S.n3195 S.n3187 0.045
R42240 S.n4332 S.n4324 0.045
R42241 S.n5467 S.n5459 0.045
R42242 S.n6577 S.n6569 0.045
R42243 S.n7675 S.n7667 0.045
R42244 S.n8750 S.n8742 0.045
R42245 S.n9813 S.n9805 0.045
R42246 S.n10853 S.n10845 0.045
R42247 S.n11881 S.n11873 0.045
R42248 S.n12886 S.n12878 0.045
R42249 S.n13879 S.n13871 0.045
R42250 S.n14849 S.n14841 0.045
R42251 S.n15807 S.n15799 0.045
R42252 S.n16742 S.n16734 0.045
R42253 S.n17665 S.n17657 0.045
R42254 S.n18565 S.n18557 0.045
R42255 S.n19446 S.n19445 0.045
R42256 S.n20318 S.n20317 0.045
R42257 S.n22984 S.n22983 0.045
R42258 S.n2546 S.n2545 0.045
R42259 S.n1353 S.n1352 0.044
R42260 S.n3759 S.n3758 0.044
R42261 S.n4887 S.n4886 0.044
R42262 S.n6007 S.n6006 0.044
R42263 S.n7100 S.n7099 0.044
R42264 S.n8184 S.n8183 0.044
R42265 S.n9242 S.n9241 0.044
R42266 S.n10291 S.n10290 0.044
R42267 S.n11314 S.n11313 0.044
R42268 S.n12328 S.n12327 0.044
R42269 S.n13316 S.n13315 0.044
R42270 S.n14295 S.n14294 0.044
R42271 S.n15248 S.n15247 0.044
R42272 S.n16192 S.n16191 0.044
R42273 S.n17110 S.n17109 0.044
R42274 S.n18019 S.n18018 0.044
R42275 S.n18902 S.n18901 0.044
R42276 S.n19774 S.n19773 0.044
R42277 S.n20877 S.n20876 0.044
R42278 S.n21687 S.n21686 0.044
R42279 S.n22675 S.n22674 0.044
R42280 S.n2628 S.n2627 0.044
R42281 S.n3775 S.n3774 0.044
R42282 S.n4903 S.n4902 0.044
R42283 S.n6023 S.n6022 0.044
R42284 S.n7116 S.n7115 0.044
R42285 S.n8200 S.n8199 0.044
R42286 S.n9258 S.n9257 0.044
R42287 S.n10307 S.n10306 0.044
R42288 S.n11330 S.n11329 0.044
R42289 S.n12344 S.n12343 0.044
R42290 S.n13332 S.n13331 0.044
R42291 S.n14311 S.n14310 0.044
R42292 S.n15264 S.n15263 0.044
R42293 S.n16208 S.n16207 0.044
R42294 S.n17126 S.n17125 0.044
R42295 S.n18035 S.n18034 0.044
R42296 S.n18918 S.n18917 0.044
R42297 S.n19790 S.n19789 0.044
R42298 S.n20861 S.n20860 0.044
R42299 S.n21656 S.n21655 0.044
R42300 S.n22982 S.n22981 0.044
R42301 S.n22807 S.n22806 0.044
R42302 S.n20845 S.n20836 0.043
R42303 S.n20210 S.n20201 0.043
R42304 S.n19340 S.n19331 0.043
R42305 S.n18458 S.n18449 0.043
R42306 S.n17553 S.n17544 0.043
R42307 S.n16635 S.n16626 0.043
R42308 S.n15695 S.n15686 0.043
R42309 S.n14742 S.n14733 0.043
R42310 S.n13767 S.n13758 0.043
R42311 S.n12779 S.n12770 0.043
R42312 S.n11769 S.n11760 0.043
R42313 S.n10746 S.n10737 0.043
R42314 S.n9701 S.n9692 0.043
R42315 S.n8643 S.n8634 0.043
R42316 S.n7563 S.n7554 0.043
R42317 S.n6470 S.n6461 0.043
R42318 S.n5354 S.n5345 0.043
R42319 S.n4225 S.n4216 0.043
R42320 S.n3084 S.n3075 0.043
R42321 S.n425 S.n424 0.043
R42322 S.n22740 S.n22739 0.043
R42323 S.n835 S.n834 0.043
R42324 S.n20282 S.n20281 0.043
R42325 S.n20353 S.n20352 0.043
R42326 S.n21229 S.n21228 0.043
R42327 S.n18611 S.n18608 0.043
R42328 S.n17711 S.n17708 0.043
R42329 S.n16849 S.n16846 0.043
R42330 S.n15914 S.n15911 0.043
R42331 S.n15017 S.n15014 0.043
R42332 S.n14047 S.n14044 0.043
R42333 S.n13115 S.n13112 0.043
R42334 S.n12110 S.n12107 0.043
R42335 S.n11143 S.n11140 0.043
R42336 S.n10103 S.n10100 0.043
R42337 S.n268 S.n267 0.043
R42338 S.n9101 S.n9098 0.043
R42339 S.n8026 S.n8023 0.043
R42340 S.n239 S.n238 0.043
R42341 S.n6989 S.n6986 0.043
R42342 S.n5879 S.n5876 0.043
R42343 S.n4805 S.n4802 0.043
R42344 S.n3661 S.n3658 0.043
R42345 S.n140 S.n139 0.043
R42346 S.n2561 S.n2558 0.043
R42347 S.n21213 S.n21210 0.043
R42348 S.n20394 S.n20391 0.043
R42349 S.n17761 S.n17758 0.043
R42350 S.n16834 S.n16831 0.043
R42351 S.n19486 S.n19483 0.043
R42352 S.n18596 S.n18593 0.043
R42353 S.n15964 S.n15961 0.043
R42354 S.n15002 S.n14999 0.043
R42355 S.n14097 S.n14094 0.043
R42356 S.n13100 S.n13097 0.043
R42357 S.n12160 S.n12157 0.043
R42358 S.n11128 S.n11125 0.043
R42359 S.n10153 S.n10150 0.043
R42360 S.n9086 S.n9083 0.043
R42361 S.n8076 S.n8073 0.043
R42362 S.n6974 S.n6971 0.043
R42363 S.n5929 S.n5926 0.043
R42364 S.n4790 S.n4787 0.043
R42365 S.n3710 S.n3708 0.043
R42366 S.n1981 S.n1980 0.043
R42367 S.n2133 S.n2132 0.043
R42368 S.n2192 S.n2191 0.043
R42369 S.n2251 S.n2250 0.043
R42370 S.n2310 S.n2309 0.043
R42371 S.n2369 S.n2368 0.043
R42372 S.n2428 S.n2427 0.043
R42373 S.n2487 S.n2486 0.043
R42374 S.n2056 S.n2055 0.043
R42375 S.n1170 S.n1169 0.043
R42376 S.n1369 S.n1368 0.043
R42377 S.n1494 S.n1493 0.042
R42378 S.n2090 S.n2089 0.042
R42379 S.n3240 S.n3239 0.042
R42380 S.n4377 S.n4376 0.042
R42381 S.n5512 S.n5511 0.042
R42382 S.n6622 S.n6621 0.042
R42383 S.n7720 S.n7719 0.042
R42384 S.n8795 S.n8794 0.042
R42385 S.n9858 S.n9857 0.042
R42386 S.n10898 S.n10897 0.042
R42387 S.n11926 S.n11925 0.042
R42388 S.n12931 S.n12930 0.042
R42389 S.n13924 S.n13923 0.042
R42390 S.n14894 S.n14893 0.042
R42391 S.n15852 S.n15851 0.042
R42392 S.n16787 S.n16786 0.042
R42393 S.n2148 S.n2147 0.042
R42394 S.n3300 S.n3299 0.042
R42395 S.n4438 S.n4437 0.042
R42396 S.n5573 S.n5572 0.042
R42397 S.n6683 S.n6682 0.042
R42398 S.n7781 S.n7780 0.042
R42399 S.n8856 S.n8855 0.042
R42400 S.n9919 S.n9918 0.042
R42401 S.n10959 S.n10958 0.042
R42402 S.n11987 S.n11986 0.042
R42403 S.n12992 S.n12991 0.042
R42404 S.n13985 S.n13984 0.042
R42405 S.n14955 S.n14954 0.042
R42406 S.n2207 S.n2206 0.042
R42407 S.n3360 S.n3359 0.042
R42408 S.n4499 S.n4498 0.042
R42409 S.n5634 S.n5633 0.042
R42410 S.n6744 S.n6743 0.042
R42411 S.n7842 S.n7841 0.042
R42412 S.n8917 S.n8916 0.042
R42413 S.n9980 S.n9979 0.042
R42414 S.n11020 S.n11019 0.042
R42415 S.n12048 S.n12047 0.042
R42416 S.n13053 S.n13052 0.042
R42417 S.n2266 S.n2265 0.042
R42418 S.n3420 S.n3419 0.042
R42419 S.n4560 S.n4559 0.042
R42420 S.n5695 S.n5694 0.042
R42421 S.n6805 S.n6804 0.042
R42422 S.n7903 S.n7902 0.042
R42423 S.n8978 S.n8977 0.042
R42424 S.n10041 S.n10040 0.042
R42425 S.n11081 S.n11080 0.042
R42426 S.n2325 S.n2324 0.042
R42427 S.n3480 S.n3479 0.042
R42428 S.n4621 S.n4620 0.042
R42429 S.n5756 S.n5755 0.042
R42430 S.n6866 S.n6865 0.042
R42431 S.n7964 S.n7963 0.042
R42432 S.n9039 S.n9038 0.042
R42433 S.n2384 S.n2383 0.042
R42434 S.n3540 S.n3539 0.042
R42435 S.n4682 S.n4681 0.042
R42436 S.n5817 S.n5816 0.042
R42437 S.n6927 S.n6926 0.042
R42438 S.n2443 S.n2442 0.042
R42439 S.n3600 S.n3599 0.042
R42440 S.n4743 S.n4742 0.042
R42441 S.n2502 S.n2501 0.042
R42442 S.n938 S.n937 0.042
R42443 S.n20267 S.n20264 0.042
R42444 S.n19399 S.n19396 0.042
R42445 S.n18512 S.n18509 0.042
R42446 S.n17612 S.n17609 0.042
R42447 S.n16689 S.n16686 0.042
R42448 S.n15754 S.n15751 0.042
R42449 S.n14796 S.n14793 0.042
R42450 S.n13826 S.n13823 0.042
R42451 S.n12833 S.n12830 0.042
R42452 S.n11828 S.n11825 0.042
R42453 S.n10800 S.n10797 0.042
R42454 S.n9760 S.n9757 0.042
R42455 S.n8697 S.n8694 0.042
R42456 S.n7622 S.n7619 0.042
R42457 S.n6524 S.n6521 0.042
R42458 S.n5413 S.n5410 0.042
R42459 S.n4279 S.n4276 0.042
R42460 S.n3142 S.n3140 0.042
R42461 S.n1861 S.n1860 0.042
R42462 S.n15899 S.n15896 0.042
R42463 S.n14941 S.n14938 0.042
R42464 S.n13971 S.n13968 0.042
R42465 S.n12978 S.n12975 0.042
R42466 S.n11973 S.n11970 0.042
R42467 S.n10945 S.n10942 0.042
R42468 S.n9905 S.n9902 0.042
R42469 S.n8842 S.n8839 0.042
R42470 S.n7767 S.n7764 0.042
R42471 S.n6669 S.n6666 0.042
R42472 S.n5559 S.n5556 0.042
R42473 S.n4424 S.n4421 0.042
R42474 S.n3286 S.n3284 0.042
R42475 S.n1753 S.n1752 0.042
R42476 S.n17696 S.n17693 0.042
R42477 S.n16773 S.n16770 0.042
R42478 S.n15838 S.n15835 0.042
R42479 S.n14880 S.n14877 0.042
R42480 S.n13910 S.n13907 0.042
R42481 S.n12917 S.n12914 0.042
R42482 S.n11912 S.n11909 0.042
R42483 S.n10884 S.n10881 0.042
R42484 S.n9844 S.n9841 0.042
R42485 S.n8781 S.n8778 0.042
R42486 S.n7706 S.n7703 0.042
R42487 S.n6608 S.n6605 0.042
R42488 S.n5498 S.n5495 0.042
R42489 S.n4363 S.n4360 0.042
R42490 S.n3226 S.n3224 0.042
R42491 S.n1786 S.n1785 0.042
R42492 S.n14032 S.n14029 0.042
R42493 S.n13039 S.n13036 0.042
R42494 S.n12034 S.n12031 0.042
R42495 S.n11006 S.n11003 0.042
R42496 S.n9966 S.n9963 0.042
R42497 S.n8903 S.n8900 0.042
R42498 S.n7828 S.n7825 0.042
R42499 S.n6730 S.n6727 0.042
R42500 S.n5620 S.n5617 0.042
R42501 S.n4485 S.n4482 0.042
R42502 S.n3346 S.n3344 0.042
R42503 S.n1716 S.n1715 0.042
R42504 S.n12095 S.n12092 0.042
R42505 S.n11067 S.n11064 0.042
R42506 S.n10027 S.n10024 0.042
R42507 S.n8964 S.n8961 0.042
R42508 S.n7889 S.n7886 0.042
R42509 S.n6791 S.n6788 0.042
R42510 S.n5681 S.n5678 0.042
R42511 S.n4546 S.n4543 0.042
R42512 S.n3406 S.n3404 0.042
R42513 S.n1679 S.n1678 0.042
R42514 S.n10088 S.n10085 0.042
R42515 S.n9025 S.n9022 0.042
R42516 S.n7950 S.n7947 0.042
R42517 S.n6852 S.n6849 0.042
R42518 S.n5742 S.n5739 0.042
R42519 S.n4607 S.n4604 0.042
R42520 S.n3466 S.n3464 0.042
R42521 S.n1642 S.n1641 0.042
R42522 S.n8011 S.n8008 0.042
R42523 S.n6913 S.n6910 0.042
R42524 S.n5803 S.n5800 0.042
R42525 S.n4668 S.n4665 0.042
R42526 S.n3526 S.n3524 0.042
R42527 S.n1605 S.n1604 0.042
R42528 S.n5864 S.n5861 0.042
R42529 S.n4729 S.n4726 0.042
R42530 S.n3586 S.n3584 0.042
R42531 S.n1568 S.n1567 0.042
R42532 S.n3646 S.n3644 0.042
R42533 S.n1531 S.n1530 0.042
R42534 S.n26 S.n25 0.042
R42535 S.n1339 S.n1338 0.042
R42536 S.n73 S.n72 0.042
R42537 S.n105 S.n104 0.042
R42538 S.n992 S.n991 0.042
R42539 S.n1024 S.n1023 0.042
R42540 S.n1056 S.n1055 0.042
R42541 S.n1088 S.n1087 0.042
R42542 S.n1120 S.n1119 0.042
R42543 S.n1158 S.n1157 0.042
R42544 S.n19413 S.n19412 0.042
R42545 S.n18526 S.n18525 0.042
R42546 S.n17626 S.n17625 0.042
R42547 S.n16703 S.n16702 0.042
R42548 S.n15768 S.n15767 0.042
R42549 S.n14810 S.n14809 0.042
R42550 S.n13840 S.n13839 0.042
R42551 S.n12847 S.n12846 0.042
R42552 S.n11842 S.n11841 0.042
R42553 S.n10814 S.n10813 0.042
R42554 S.n9774 S.n9773 0.042
R42555 S.n8711 S.n8710 0.042
R42556 S.n7636 S.n7635 0.042
R42557 S.n6538 S.n6537 0.042
R42558 S.n5427 S.n5426 0.042
R42559 S.n4293 S.n4292 0.042
R42560 S.n3156 S.n3155 0.042
R42561 S.n1995 S.n1994 0.042
R42562 S.n20221 S.n20220 0.041
R42563 S.n1373 S.n1372 0.041
R42564 S.n4 S.n3 0.041
R42565 S.n51 S.n50 0.041
R42566 S.n82 S.n81 0.041
R42567 S.n114 S.n113 0.041
R42568 S.n1001 S.n1000 0.041
R42569 S.n1033 S.n1032 0.041
R42570 S.n1065 S.n1064 0.041
R42571 S.n1097 S.n1096 0.041
R42572 S.n1129 S.n1128 0.041
R42573 S.n1167 S.n1166 0.041
R42574 S.n1182 S.n1180 0.041
R42575 S.n952 S.n951 0.041
R42576 S.n1356 S.n1355 0.04
R42577 S.n88 S.n87 0.04
R42578 S.n1039 S.n1038 0.04
R42579 S.n428 S.n419 0.04
R42580 S.n1456 S.n1448 0.04
R42581 S.n2650 S.n2643 0.04
R42582 S.n3795 S.n3788 0.04
R42583 S.n4925 S.n4918 0.04
R42584 S.n6043 S.n6036 0.04
R42585 S.n7138 S.n7131 0.04
R42586 S.n8220 S.n8213 0.04
R42587 S.n9280 S.n9273 0.04
R42588 S.n10327 S.n10320 0.04
R42589 S.n11352 S.n11345 0.04
R42590 S.n12364 S.n12357 0.04
R42591 S.n13354 S.n13347 0.04
R42592 S.n14331 S.n14324 0.04
R42593 S.n15286 S.n15279 0.04
R42594 S.n16228 S.n16221 0.04
R42595 S.n17148 S.n17141 0.04
R42596 S.n18055 S.n18048 0.04
R42597 S.n18940 S.n18933 0.04
R42598 S.n19810 S.n19803 0.04
R42599 S.n20448 S.n20441 0.04
R42600 S.n21292 S.n21285 0.04
R42601 S.n22285 S.n22284 0.04
R42602 S.n1179 S.n1178 0.039
R42603 S.n427 S.n420 0.039
R42604 S.n1455 S.n1450 0.039
R42605 S.n2649 S.n2644 0.039
R42606 S.n3794 S.n3789 0.039
R42607 S.n4924 S.n4919 0.039
R42608 S.n6042 S.n6037 0.039
R42609 S.n7137 S.n7132 0.039
R42610 S.n8219 S.n8214 0.039
R42611 S.n9279 S.n9274 0.039
R42612 S.n10326 S.n10321 0.039
R42613 S.n11351 S.n11346 0.039
R42614 S.n12363 S.n12358 0.039
R42615 S.n13353 S.n13348 0.039
R42616 S.n14330 S.n14325 0.039
R42617 S.n15285 S.n15280 0.039
R42618 S.n16227 S.n16222 0.039
R42619 S.n17147 S.n17142 0.039
R42620 S.n18054 S.n18049 0.039
R42621 S.n18939 S.n18934 0.039
R42622 S.n19809 S.n19804 0.039
R42623 S.n20447 S.n20442 0.039
R42624 S.n21291 S.n21286 0.039
R42625 S.n22283 S.n22282 0.039
R42626 S.n22980 S.n22967 0.039
R42627 S.n22970 S.n22969 0.039
R42628 S.n22274 S.n22272 0.038
R42629 S.n19848 S.n19846 0.038
R42630 S.n20459 S.n20457 0.038
R42631 S.n21284 S.n21282 0.038
R42632 S.n18067 S.n18066 0.038
R42633 S.n17178 S.n17177 0.038
R42634 S.n16240 S.n16239 0.038
R42635 S.n15316 S.n15315 0.038
R42636 S.n14343 S.n14342 0.038
R42637 S.n13384 S.n13383 0.038
R42638 S.n12376 S.n12375 0.038
R42639 S.n11382 S.n11381 0.038
R42640 S.n10339 S.n10338 0.038
R42641 S.n9310 S.n9309 0.038
R42642 S.n8232 S.n8231 0.038
R42643 S.n7168 S.n7167 0.038
R42644 S.n6055 S.n6054 0.038
R42645 S.n4955 S.n4954 0.038
R42646 S.n3807 S.n3806 0.038
R42647 S.n2680 S.n2679 0.038
R42648 S.n1468 S.n1467 0.038
R42649 S.n21201 S.n21200 0.038
R42650 S.n20382 S.n20381 0.038
R42651 S.n20255 S.n20254 0.038
R42652 S.n19387 S.n19386 0.038
R42653 S.n18500 S.n18499 0.038
R42654 S.n17600 S.n17599 0.038
R42655 S.n16677 S.n16676 0.038
R42656 S.n15742 S.n15741 0.038
R42657 S.n14784 S.n14783 0.038
R42658 S.n13814 S.n13813 0.038
R42659 S.n12821 S.n12820 0.038
R42660 S.n11816 S.n11815 0.038
R42661 S.n10788 S.n10787 0.038
R42662 S.n9748 S.n9747 0.038
R42663 S.n8685 S.n8684 0.038
R42664 S.n7610 S.n7609 0.038
R42665 S.n6512 S.n6511 0.038
R42666 S.n5401 S.n5400 0.038
R42667 S.n4267 S.n4266 0.038
R42668 S.n3131 S.n3130 0.038
R42669 S.n1971 S.n1970 0.038
R42670 S.n17749 S.n17748 0.038
R42671 S.n16822 S.n16821 0.038
R42672 S.n15887 S.n15886 0.038
R42673 S.n14929 S.n14928 0.038
R42674 S.n13959 S.n13958 0.038
R42675 S.n12966 S.n12965 0.038
R42676 S.n11961 S.n11960 0.038
R42677 S.n10933 S.n10932 0.038
R42678 S.n9893 S.n9892 0.038
R42679 S.n8830 S.n8829 0.038
R42680 S.n7755 S.n7754 0.038
R42681 S.n6657 S.n6656 0.038
R42682 S.n5547 S.n5546 0.038
R42683 S.n4412 S.n4411 0.038
R42684 S.n3275 S.n3274 0.038
R42685 S.n2123 S.n2122 0.038
R42686 S.n18631 S.n18626 0.038
R42687 S.n17731 S.n17726 0.038
R42688 S.n16804 S.n16799 0.038
R42689 S.n15869 S.n15864 0.038
R42690 S.n14911 S.n14906 0.038
R42691 S.n13941 S.n13936 0.038
R42692 S.n12948 S.n12943 0.038
R42693 S.n11943 S.n11938 0.038
R42694 S.n10915 S.n10910 0.038
R42695 S.n9875 S.n9870 0.038
R42696 S.n8812 S.n8807 0.038
R42697 S.n7737 S.n7732 0.038
R42698 S.n6639 S.n6634 0.038
R42699 S.n5529 S.n5524 0.038
R42700 S.n4394 S.n4389 0.038
R42701 S.n3257 S.n3252 0.038
R42702 S.n2105 S.n2101 0.038
R42703 S.n15952 S.n15951 0.038
R42704 S.n14990 S.n14989 0.038
R42705 S.n14020 S.n14019 0.038
R42706 S.n13027 S.n13026 0.038
R42707 S.n12022 S.n12021 0.038
R42708 S.n10994 S.n10993 0.038
R42709 S.n9954 S.n9953 0.038
R42710 S.n8891 S.n8890 0.038
R42711 S.n7816 S.n7815 0.038
R42712 S.n6718 S.n6717 0.038
R42713 S.n5608 S.n5607 0.038
R42714 S.n4473 S.n4472 0.038
R42715 S.n3335 S.n3334 0.038
R42716 S.n2182 S.n2181 0.038
R42717 S.n16869 S.n16864 0.038
R42718 S.n15934 S.n15929 0.038
R42719 S.n14972 S.n14967 0.038
R42720 S.n14002 S.n13997 0.038
R42721 S.n13009 S.n13004 0.038
R42722 S.n12004 S.n11999 0.038
R42723 S.n10976 S.n10971 0.038
R42724 S.n9936 S.n9931 0.038
R42725 S.n8873 S.n8868 0.038
R42726 S.n7798 S.n7793 0.038
R42727 S.n6700 S.n6695 0.038
R42728 S.n5590 S.n5585 0.038
R42729 S.n4455 S.n4450 0.038
R42730 S.n3317 S.n3312 0.038
R42731 S.n2164 S.n2159 0.038
R42732 S.n14085 S.n14084 0.038
R42733 S.n13088 S.n13087 0.038
R42734 S.n12083 S.n12082 0.038
R42735 S.n11055 S.n11054 0.038
R42736 S.n10015 S.n10014 0.038
R42737 S.n8952 S.n8951 0.038
R42738 S.n7877 S.n7876 0.038
R42739 S.n6779 S.n6778 0.038
R42740 S.n5669 S.n5668 0.038
R42741 S.n4534 S.n4533 0.038
R42742 S.n3395 S.n3394 0.038
R42743 S.n2241 S.n2240 0.038
R42744 S.n15037 S.n15032 0.038
R42745 S.n14067 S.n14062 0.038
R42746 S.n13070 S.n13065 0.038
R42747 S.n12065 S.n12060 0.038
R42748 S.n11037 S.n11032 0.038
R42749 S.n9997 S.n9992 0.038
R42750 S.n8934 S.n8929 0.038
R42751 S.n7859 S.n7854 0.038
R42752 S.n6761 S.n6756 0.038
R42753 S.n5651 S.n5646 0.038
R42754 S.n4516 S.n4511 0.038
R42755 S.n3377 S.n3372 0.038
R42756 S.n2223 S.n2218 0.038
R42757 S.n12148 S.n12147 0.038
R42758 S.n11116 S.n11115 0.038
R42759 S.n10076 S.n10075 0.038
R42760 S.n9013 S.n9012 0.038
R42761 S.n7938 S.n7937 0.038
R42762 S.n6840 S.n6839 0.038
R42763 S.n5730 S.n5729 0.038
R42764 S.n4595 S.n4594 0.038
R42765 S.n3455 S.n3454 0.038
R42766 S.n2300 S.n2299 0.038
R42767 S.n13135 S.n13130 0.038
R42768 S.n12130 S.n12125 0.038
R42769 S.n11098 S.n11093 0.038
R42770 S.n10058 S.n10053 0.038
R42771 S.n8995 S.n8990 0.038
R42772 S.n7920 S.n7915 0.038
R42773 S.n6822 S.n6817 0.038
R42774 S.n5712 S.n5707 0.038
R42775 S.n4577 S.n4572 0.038
R42776 S.n3437 S.n3432 0.038
R42777 S.n2282 S.n2277 0.038
R42778 S.n10141 S.n10140 0.038
R42779 S.n9074 S.n9073 0.038
R42780 S.n7999 S.n7998 0.038
R42781 S.n6901 S.n6900 0.038
R42782 S.n5791 S.n5790 0.038
R42783 S.n4656 S.n4655 0.038
R42784 S.n3515 S.n3514 0.038
R42785 S.n2359 S.n2358 0.038
R42786 S.n11163 S.n11158 0.038
R42787 S.n10123 S.n10118 0.038
R42788 S.n9056 S.n9051 0.038
R42789 S.n7981 S.n7976 0.038
R42790 S.n6883 S.n6878 0.038
R42791 S.n5773 S.n5768 0.038
R42792 S.n4638 S.n4633 0.038
R42793 S.n3497 S.n3492 0.038
R42794 S.n2341 S.n2336 0.038
R42795 S.n8064 S.n8063 0.038
R42796 S.n6962 S.n6961 0.038
R42797 S.n5852 S.n5851 0.038
R42798 S.n4717 S.n4716 0.038
R42799 S.n3575 S.n3574 0.038
R42800 S.n2418 S.n2417 0.038
R42801 S.n9121 S.n9116 0.038
R42802 S.n8046 S.n8041 0.038
R42803 S.n6944 S.n6939 0.038
R42804 S.n5834 S.n5829 0.038
R42805 S.n4699 S.n4694 0.038
R42806 S.n3557 S.n3552 0.038
R42807 S.n2400 S.n2395 0.038
R42808 S.n5917 S.n5916 0.038
R42809 S.n4778 S.n4777 0.038
R42810 S.n3635 S.n3634 0.038
R42811 S.n2477 S.n2476 0.038
R42812 S.n7009 S.n7004 0.038
R42813 S.n5899 S.n5894 0.038
R42814 S.n4760 S.n4755 0.038
R42815 S.n3617 S.n3612 0.038
R42816 S.n2459 S.n2454 0.038
R42817 S.n3699 S.n3698 0.038
R42818 S.n2536 S.n2535 0.038
R42819 S.n4825 S.n4820 0.038
R42820 S.n3681 S.n3676 0.038
R42821 S.n2518 S.n2513 0.038
R42822 S.n2581 S.n2576 0.038
R42823 S.n3198 S.n3180 0.038
R42824 S.n4335 S.n4317 0.038
R42825 S.n5470 S.n5452 0.038
R42826 S.n6580 S.n6562 0.038
R42827 S.n7678 S.n7660 0.038
R42828 S.n8753 S.n8735 0.038
R42829 S.n9816 S.n9798 0.038
R42830 S.n10856 S.n10838 0.038
R42831 S.n11884 S.n11866 0.038
R42832 S.n12889 S.n12871 0.038
R42833 S.n13882 S.n13864 0.038
R42834 S.n14852 S.n14834 0.038
R42835 S.n15810 S.n15792 0.038
R42836 S.n16745 S.n16727 0.038
R42837 S.n17668 S.n17650 0.038
R42838 S.n18568 S.n18550 0.038
R42839 S.n19458 S.n19437 0.038
R42840 S.n20330 S.n20309 0.038
R42841 S.n20424 S.n20413 0.038
R42842 S.n2045 S.n2040 0.038
R42843 S.n2598 S.n1900 0.038
R42844 S.n20423 S.n20421 0.037
R42845 S.n2012 S.n2004 0.037
R42846 S.n21986 S.n21985 0.037
R42847 S.n21952 S.n21951 0.037
R42848 S.n1431 S.n1430 0.036
R42849 S.n974 S.n952 0.036
R42850 S.n1844 S.n1843 0.036
R42851 S.n2994 S.n2993 0.036
R42852 S.n4121 S.n4120 0.036
R42853 S.n5233 S.n5232 0.036
R42854 S.n6333 S.n6332 0.036
R42855 S.n7410 S.n7409 0.036
R42856 S.n8474 S.n8473 0.036
R42857 S.n9516 S.n9515 0.036
R42858 S.n10545 S.n10544 0.036
R42859 S.n11552 S.n11551 0.036
R42860 S.n12546 S.n12545 0.036
R42861 S.n13518 S.n13517 0.036
R42862 S.n14477 S.n14476 0.036
R42863 S.n15414 S.n15413 0.036
R42864 S.n16338 S.n16337 0.036
R42865 S.n17240 S.n17239 0.036
R42866 S.n18129 S.n18128 0.036
R42867 S.n18995 S.n18994 0.036
R42868 S.n22756 S.n22755 0.036
R42869 S.n16277 S.n16276 0.035
R42870 S.n15353 S.n15352 0.035
R42871 S.n14416 S.n14415 0.035
R42872 S.n13457 S.n13456 0.035
R42873 S.n12485 S.n12484 0.035
R42874 S.n11491 S.n11490 0.035
R42875 S.n10484 S.n10483 0.035
R42876 S.n9455 S.n9454 0.035
R42877 S.n8413 S.n8412 0.035
R42878 S.n7349 S.n7348 0.035
R42879 S.n6272 S.n6271 0.035
R42880 S.n5172 S.n5171 0.035
R42881 S.n4060 S.n4059 0.035
R42882 S.n2933 S.n2932 0.035
R42883 S.n1765 S.n1764 0.035
R42884 S.n14380 S.n14379 0.035
R42885 S.n13421 S.n13420 0.035
R42886 S.n12449 S.n12448 0.035
R42887 S.n11455 S.n11454 0.035
R42888 S.n10448 S.n10447 0.035
R42889 S.n9419 S.n9418 0.035
R42890 S.n8377 S.n8376 0.035
R42891 S.n7313 S.n7312 0.035
R42892 S.n6236 S.n6235 0.035
R42893 S.n5136 S.n5135 0.035
R42894 S.n4024 S.n4023 0.035
R42895 S.n2897 S.n2896 0.035
R42896 S.n1728 S.n1727 0.035
R42897 S.n12413 S.n12412 0.035
R42898 S.n11419 S.n11418 0.035
R42899 S.n10412 S.n10411 0.035
R42900 S.n9383 S.n9382 0.035
R42901 S.n8341 S.n8340 0.035
R42902 S.n7277 S.n7276 0.035
R42903 S.n6200 S.n6199 0.035
R42904 S.n5100 S.n5099 0.035
R42905 S.n3988 S.n3987 0.035
R42906 S.n2861 S.n2860 0.035
R42907 S.n1691 S.n1690 0.035
R42908 S.n10376 S.n10375 0.035
R42909 S.n9347 S.n9346 0.035
R42910 S.n8305 S.n8304 0.035
R42911 S.n7241 S.n7240 0.035
R42912 S.n6164 S.n6163 0.035
R42913 S.n5064 S.n5063 0.035
R42914 S.n3952 S.n3951 0.035
R42915 S.n2825 S.n2824 0.035
R42916 S.n1654 S.n1653 0.035
R42917 S.n8269 S.n8268 0.035
R42918 S.n7205 S.n7204 0.035
R42919 S.n6128 S.n6127 0.035
R42920 S.n5028 S.n5027 0.035
R42921 S.n3916 S.n3915 0.035
R42922 S.n2789 S.n2788 0.035
R42923 S.n1617 S.n1616 0.035
R42924 S.n6092 S.n6091 0.035
R42925 S.n4992 S.n4991 0.035
R42926 S.n3880 S.n3879 0.035
R42927 S.n2753 S.n2752 0.035
R42928 S.n1580 S.n1579 0.035
R42929 S.n3844 S.n3843 0.035
R42930 S.n2717 S.n2716 0.035
R42931 S.n1543 S.n1542 0.035
R42932 S.n1506 S.n1505 0.035
R42933 S.n22834 S.n22833 0.035
R42934 S.n22825 S.n22824 0.035
R42935 S.n22721 S.n22720 0.035
R42936 S.n22293 S.n22292 0.035
R42937 S.n18064 S.n18063 0.035
R42938 S.n18948 S.n18947 0.035
R42939 S.n19819 S.n19818 0.035
R42940 S.n20456 S.n20455 0.035
R42941 S.n21301 S.n21300 0.035
R42942 S.n16237 S.n16236 0.035
R42943 S.n17156 S.n17155 0.035
R42944 S.n14340 S.n14339 0.035
R42945 S.n15294 S.n15293 0.035
R42946 S.n12373 S.n12372 0.035
R42947 S.n13362 S.n13361 0.035
R42948 S.n10336 S.n10335 0.035
R42949 S.n11360 S.n11359 0.035
R42950 S.n8229 S.n8228 0.035
R42951 S.n9288 S.n9287 0.035
R42952 S.n6052 S.n6051 0.035
R42953 S.n7146 S.n7145 0.035
R42954 S.n3804 S.n3803 0.035
R42955 S.n4933 S.n4932 0.035
R42956 S.n1465 S.n1464 0.035
R42957 S.n2658 S.n2657 0.035
R42958 S.n437 S.n436 0.035
R42959 S.n21201 S.n21196 0.035
R42960 S.n20382 S.n20377 0.035
R42961 S.n20255 S.n20250 0.035
R42962 S.n19387 S.n19382 0.035
R42963 S.n18500 S.n18495 0.035
R42964 S.n17600 S.n17595 0.035
R42965 S.n16677 S.n16672 0.035
R42966 S.n15742 S.n15737 0.035
R42967 S.n14784 S.n14779 0.035
R42968 S.n13814 S.n13809 0.035
R42969 S.n12821 S.n12816 0.035
R42970 S.n11816 S.n11811 0.035
R42971 S.n10788 S.n10783 0.035
R42972 S.n9748 S.n9743 0.035
R42973 S.n8685 S.n8680 0.035
R42974 S.n7610 S.n7605 0.035
R42975 S.n6512 S.n6507 0.035
R42976 S.n5401 S.n5396 0.035
R42977 S.n4267 S.n4262 0.035
R42978 S.n3131 S.n3126 0.035
R42979 S.n1971 S.n1966 0.035
R42980 S.n17749 S.n17744 0.035
R42981 S.n16822 S.n16817 0.035
R42982 S.n15887 S.n15882 0.035
R42983 S.n14929 S.n14924 0.035
R42984 S.n13959 S.n13954 0.035
R42985 S.n12966 S.n12961 0.035
R42986 S.n11961 S.n11956 0.035
R42987 S.n10933 S.n10928 0.035
R42988 S.n9893 S.n9888 0.035
R42989 S.n8830 S.n8825 0.035
R42990 S.n7755 S.n7750 0.035
R42991 S.n6657 S.n6652 0.035
R42992 S.n5547 S.n5542 0.035
R42993 S.n4412 S.n4407 0.035
R42994 S.n3275 S.n3270 0.035
R42995 S.n2123 S.n2118 0.035
R42996 S.n20238 S.n20221 0.035
R42997 S.n20327 S.n20326 0.035
R42998 S.n19455 S.n19454 0.035
R42999 S.n2105 S.n2104 0.035
R43000 S.n3257 S.n3256 0.035
R43001 S.n4394 S.n4393 0.035
R43002 S.n5529 S.n5528 0.035
R43003 S.n6639 S.n6638 0.035
R43004 S.n7737 S.n7736 0.035
R43005 S.n8812 S.n8811 0.035
R43006 S.n9875 S.n9874 0.035
R43007 S.n10915 S.n10914 0.035
R43008 S.n11943 S.n11942 0.035
R43009 S.n12948 S.n12947 0.035
R43010 S.n13941 S.n13940 0.035
R43011 S.n14911 S.n14910 0.035
R43012 S.n15869 S.n15868 0.035
R43013 S.n16804 S.n16803 0.035
R43014 S.n17731 S.n17730 0.035
R43015 S.n18631 S.n18630 0.035
R43016 S.n15952 S.n15947 0.035
R43017 S.n14990 S.n14985 0.035
R43018 S.n14020 S.n14015 0.035
R43019 S.n13027 S.n13022 0.035
R43020 S.n12022 S.n12017 0.035
R43021 S.n10994 S.n10989 0.035
R43022 S.n9954 S.n9949 0.035
R43023 S.n8891 S.n8886 0.035
R43024 S.n7816 S.n7811 0.035
R43025 S.n6718 S.n6713 0.035
R43026 S.n5608 S.n5603 0.035
R43027 S.n4473 S.n4468 0.035
R43028 S.n3335 S.n3330 0.035
R43029 S.n2182 S.n2177 0.035
R43030 S.n2164 S.n2163 0.035
R43031 S.n3317 S.n3316 0.035
R43032 S.n4455 S.n4454 0.035
R43033 S.n5590 S.n5589 0.035
R43034 S.n6700 S.n6699 0.035
R43035 S.n7798 S.n7797 0.035
R43036 S.n8873 S.n8872 0.035
R43037 S.n9936 S.n9935 0.035
R43038 S.n10976 S.n10975 0.035
R43039 S.n12004 S.n12003 0.035
R43040 S.n13009 S.n13008 0.035
R43041 S.n14002 S.n14001 0.035
R43042 S.n14972 S.n14971 0.035
R43043 S.n15934 S.n15933 0.035
R43044 S.n16869 S.n16868 0.035
R43045 S.n14085 S.n14080 0.035
R43046 S.n13088 S.n13083 0.035
R43047 S.n12083 S.n12078 0.035
R43048 S.n11055 S.n11050 0.035
R43049 S.n10015 S.n10010 0.035
R43050 S.n8952 S.n8947 0.035
R43051 S.n7877 S.n7872 0.035
R43052 S.n6779 S.n6774 0.035
R43053 S.n5669 S.n5664 0.035
R43054 S.n4534 S.n4529 0.035
R43055 S.n3395 S.n3390 0.035
R43056 S.n2241 S.n2236 0.035
R43057 S.n2223 S.n2222 0.035
R43058 S.n3377 S.n3376 0.035
R43059 S.n4516 S.n4515 0.035
R43060 S.n5651 S.n5650 0.035
R43061 S.n6761 S.n6760 0.035
R43062 S.n7859 S.n7858 0.035
R43063 S.n8934 S.n8933 0.035
R43064 S.n9997 S.n9996 0.035
R43065 S.n11037 S.n11036 0.035
R43066 S.n12065 S.n12064 0.035
R43067 S.n13070 S.n13069 0.035
R43068 S.n14067 S.n14066 0.035
R43069 S.n15037 S.n15036 0.035
R43070 S.n12148 S.n12143 0.035
R43071 S.n11116 S.n11111 0.035
R43072 S.n10076 S.n10071 0.035
R43073 S.n9013 S.n9008 0.035
R43074 S.n7938 S.n7933 0.035
R43075 S.n6840 S.n6835 0.035
R43076 S.n5730 S.n5725 0.035
R43077 S.n4595 S.n4590 0.035
R43078 S.n3455 S.n3450 0.035
R43079 S.n2300 S.n2295 0.035
R43080 S.n2282 S.n2281 0.035
R43081 S.n3437 S.n3436 0.035
R43082 S.n4577 S.n4576 0.035
R43083 S.n5712 S.n5711 0.035
R43084 S.n6822 S.n6821 0.035
R43085 S.n7920 S.n7919 0.035
R43086 S.n8995 S.n8994 0.035
R43087 S.n10058 S.n10057 0.035
R43088 S.n11098 S.n11097 0.035
R43089 S.n12130 S.n12129 0.035
R43090 S.n13135 S.n13134 0.035
R43091 S.n10141 S.n10136 0.035
R43092 S.n9074 S.n9069 0.035
R43093 S.n7999 S.n7994 0.035
R43094 S.n6901 S.n6896 0.035
R43095 S.n5791 S.n5786 0.035
R43096 S.n4656 S.n4651 0.035
R43097 S.n3515 S.n3510 0.035
R43098 S.n2359 S.n2354 0.035
R43099 S.n2341 S.n2340 0.035
R43100 S.n3497 S.n3496 0.035
R43101 S.n4638 S.n4637 0.035
R43102 S.n5773 S.n5772 0.035
R43103 S.n6883 S.n6882 0.035
R43104 S.n7981 S.n7980 0.035
R43105 S.n9056 S.n9055 0.035
R43106 S.n10123 S.n10122 0.035
R43107 S.n11163 S.n11162 0.035
R43108 S.n8064 S.n8059 0.035
R43109 S.n6962 S.n6957 0.035
R43110 S.n5852 S.n5847 0.035
R43111 S.n4717 S.n4712 0.035
R43112 S.n3575 S.n3570 0.035
R43113 S.n2418 S.n2413 0.035
R43114 S.n2400 S.n2399 0.035
R43115 S.n3557 S.n3556 0.035
R43116 S.n4699 S.n4698 0.035
R43117 S.n5834 S.n5833 0.035
R43118 S.n6944 S.n6943 0.035
R43119 S.n8046 S.n8045 0.035
R43120 S.n9121 S.n9120 0.035
R43121 S.n5917 S.n5912 0.035
R43122 S.n4778 S.n4773 0.035
R43123 S.n3635 S.n3630 0.035
R43124 S.n2477 S.n2472 0.035
R43125 S.n2459 S.n2458 0.035
R43126 S.n3617 S.n3616 0.035
R43127 S.n4760 S.n4759 0.035
R43128 S.n5899 S.n5898 0.035
R43129 S.n7009 S.n7008 0.035
R43130 S.n3699 S.n3694 0.035
R43131 S.n2536 S.n2531 0.035
R43132 S.n2518 S.n2517 0.035
R43133 S.n3681 S.n3680 0.035
R43134 S.n4825 S.n4824 0.035
R43135 S.n2581 S.n2580 0.035
R43136 S.t41 S.n22955 0.035
R43137 S.t41 S.n22962 0.035
R43138 S.t41 S.n22948 0.035
R43139 S.t41 S.n22941 0.035
R43140 S.t41 S.n22934 0.035
R43141 S.t41 S.n22927 0.035
R43142 S.t41 S.n22920 0.035
R43143 S.t41 S.n22913 0.035
R43144 S.t41 S.n22906 0.035
R43145 S.t41 S.n22899 0.035
R43146 S.t41 S.n22892 0.035
R43147 S.t41 S.n22885 0.035
R43148 S.t41 S.n22878 0.035
R43149 S.t41 S.n22871 0.035
R43150 S.t41 S.n22864 0.035
R43151 S.t41 S.n22857 0.035
R43152 S.t41 S.n22850 0.035
R43153 S.t41 S.n22843 0.035
R43154 S.t41 S.n22836 0.035
R43155 S.t41 S.n22827 0.035
R43156 S.t41 S.n22816 0.035
R43157 S.t41 S.n22818 0.035
R43158 S.t158 S.n1294 0.035
R43159 S.t158 S.n1416 0.035
R43160 S.t158 S.n1308 0.035
R43161 S.t158 S.n1319 0.035
R43162 S.t158 S.n1367 0.035
R43163 S.t158 S.n1282 0.035
R43164 S.t158 S.n1412 0.035
R43165 S.t158 S.n1269 0.035
R43166 S.t158 S.n1408 0.035
R43167 S.t158 S.n1256 0.035
R43168 S.t158 S.n1404 0.035
R43169 S.t158 S.n1243 0.035
R43170 S.t158 S.n1400 0.035
R43171 S.t158 S.n1230 0.035
R43172 S.t158 S.n1396 0.035
R43173 S.t158 S.n1217 0.035
R43174 S.t158 S.n1392 0.035
R43175 S.t158 S.n1204 0.035
R43176 S.t158 S.n1388 0.035
R43177 S.t158 S.n1191 0.035
R43178 S.t158 S.n1384 0.035
R43179 S.t158 S.n1380 0.035
R43180 S.t41 S.n22993 0.035
R43181 S.n22810 S.n22809 0.035
R43182 S.n1305 S.n1301 0.034
R43183 S.n1298 S.n1297 0.034
R43184 S.n1286 S.n1285 0.034
R43185 S.n1274 S.n1273 0.034
R43186 S.n1261 S.n1260 0.034
R43187 S.n1248 S.n1247 0.034
R43188 S.n1235 S.n1234 0.034
R43189 S.n1222 S.n1221 0.034
R43190 S.n1209 S.n1208 0.034
R43191 S.n1196 S.n1195 0.034
R43192 S.n3728 S.n2618 0.034
R43193 S.n2597 S.n1918 0.034
R43194 S.n910 S.n909 0.034
R43195 S.n19812 S.n19802 0.034
R43196 S.n18942 S.n18932 0.034
R43197 S.n18057 S.n18047 0.034
R43198 S.n17150 S.n17140 0.034
R43199 S.n16230 S.n16220 0.034
R43200 S.n15288 S.n15278 0.034
R43201 S.n14333 S.n14323 0.034
R43202 S.n13356 S.n13346 0.034
R43203 S.n12366 S.n12356 0.034
R43204 S.n11354 S.n11344 0.034
R43205 S.n10329 S.n10319 0.034
R43206 S.n9282 S.n9272 0.034
R43207 S.n8222 S.n8212 0.034
R43208 S.n7140 S.n7130 0.034
R43209 S.n6045 S.n6035 0.034
R43210 S.n4927 S.n4917 0.034
R43211 S.n3797 S.n3787 0.034
R43212 S.n1458 S.n1447 0.034
R43213 S.n2652 S.n2642 0.034
R43214 S.n430 S.n418 0.034
R43215 S.t41 S.n22958 0.034
R43216 S.t41 S.n22965 0.034
R43217 S.t41 S.n22951 0.034
R43218 S.t41 S.n22944 0.034
R43219 S.t41 S.n22937 0.034
R43220 S.t41 S.n22930 0.034
R43221 S.t41 S.n22923 0.034
R43222 S.t41 S.n22916 0.034
R43223 S.t41 S.n22909 0.034
R43224 S.t41 S.n22902 0.034
R43225 S.t41 S.n22895 0.034
R43226 S.t41 S.n22888 0.034
R43227 S.t41 S.n22881 0.034
R43228 S.t41 S.n22874 0.034
R43229 S.t41 S.n22867 0.034
R43230 S.t41 S.n22860 0.034
R43231 S.t41 S.n22853 0.034
R43232 S.t41 S.n22846 0.034
R43233 S.t41 S.n22839 0.034
R43234 S.t41 S.n22830 0.034
R43235 S.t41 S.n22813 0.034
R43236 S.t41 S.n22821 0.034
R43237 S.t158 S.n1293 0.034
R43238 S.t158 S.n1419 0.034
R43239 S.t158 S.n1307 0.034
R43240 S.t158 S.n1318 0.034
R43241 S.t158 S.n1366 0.034
R43242 S.t158 S.n1281 0.034
R43243 S.t158 S.n1415 0.034
R43244 S.t158 S.n1268 0.034
R43245 S.t158 S.n1411 0.034
R43246 S.t158 S.n1255 0.034
R43247 S.t158 S.n1407 0.034
R43248 S.t158 S.n1242 0.034
R43249 S.t158 S.n1403 0.034
R43250 S.t158 S.n1229 0.034
R43251 S.t158 S.n1399 0.034
R43252 S.t158 S.n1216 0.034
R43253 S.t158 S.n1395 0.034
R43254 S.t158 S.n1203 0.034
R43255 S.t158 S.n1391 0.034
R43256 S.t158 S.n1190 0.034
R43257 S.t158 S.n1387 0.034
R43258 S.t158 S.n1383 0.034
R43259 S.t41 S.n22996 0.034
R43260 S.n1798 S.n1797 0.033
R43261 S.n22306 S.n22305 0.033
R43262 S.n1182 S.n1181 0.032
R43263 S.n22287 S.n22274 0.032
R43264 S.n19849 S.n19848 0.032
R43265 S.n20460 S.n20459 0.032
R43266 S.n21294 S.n21284 0.032
R43267 S.n1833 S.n1832 0.032
R43268 S.n1947 S.n1946 0.031
R43269 S.n18068 S.n18067 0.031
R43270 S.n17179 S.n17178 0.031
R43271 S.n16241 S.n16240 0.031
R43272 S.n15317 S.n15316 0.031
R43273 S.n14344 S.n14343 0.031
R43274 S.n13385 S.n13384 0.031
R43275 S.n12377 S.n12376 0.031
R43276 S.n11383 S.n11382 0.031
R43277 S.n10340 S.n10339 0.031
R43278 S.n9311 S.n9310 0.031
R43279 S.n8233 S.n8232 0.031
R43280 S.n7169 S.n7168 0.031
R43281 S.n6056 S.n6055 0.031
R43282 S.n4956 S.n4955 0.031
R43283 S.n3808 S.n3807 0.031
R43284 S.n2681 S.n2680 0.031
R43285 S.n1469 S.n1468 0.031
R43286 S.t88 S.n22721 0.031
R43287 S.t9 S.n22293 0.031
R43288 S.t79 S.n18064 0.031
R43289 S.t150 S.n18948 0.031
R43290 S.t209 S.n19819 0.031
R43291 S.t64 S.n20456 0.031
R43292 S.t100 S.n21301 0.031
R43293 S.t167 S.n16237 0.031
R43294 S.t218 S.n17156 0.031
R43295 S.t0 S.n14340 0.031
R43296 S.t60 S.n15294 0.031
R43297 S.t357 S.n12373 0.031
R43298 S.t73 S.n13362 0.031
R43299 S.t31 S.n10336 0.031
R43300 S.t54 S.n11360 0.031
R43301 S.t19 S.n8229 0.031
R43302 S.t366 S.n9288 0.031
R43303 S.t83 S.n6052 0.031
R43304 S.t47 S.n7146 0.031
R43305 S.t176 S.n3804 0.031
R43306 S.t214 S.n4933 0.031
R43307 S.t75 S.n1465 0.031
R43308 S.t14 S.n2658 0.031
R43309 S.t137 S.n437 0.031
R43310 S.n21196 S.n21195 0.031
R43311 S.n20377 S.n20376 0.031
R43312 S.n20250 S.n20249 0.031
R43313 S.n19382 S.n19381 0.031
R43314 S.n18495 S.n18494 0.031
R43315 S.n17595 S.n17594 0.031
R43316 S.n16672 S.n16671 0.031
R43317 S.n15737 S.n15736 0.031
R43318 S.n14779 S.n14778 0.031
R43319 S.n13809 S.n13808 0.031
R43320 S.n12816 S.n12815 0.031
R43321 S.n11811 S.n11810 0.031
R43322 S.n10783 S.n10782 0.031
R43323 S.n9743 S.n9742 0.031
R43324 S.n8680 S.n8679 0.031
R43325 S.n7605 S.n7604 0.031
R43326 S.n6507 S.n6506 0.031
R43327 S.n5396 S.n5395 0.031
R43328 S.n4262 S.n4261 0.031
R43329 S.n3126 S.n3125 0.031
R43330 S.n1966 S.n1965 0.031
R43331 S.n950 S.n949 0.031
R43332 S.n17744 S.n17743 0.031
R43333 S.n16817 S.n16816 0.031
R43334 S.n15882 S.n15881 0.031
R43335 S.n14924 S.n14923 0.031
R43336 S.n13954 S.n13953 0.031
R43337 S.n12961 S.n12960 0.031
R43338 S.n11956 S.n11955 0.031
R43339 S.n10928 S.n10927 0.031
R43340 S.n9888 S.n9887 0.031
R43341 S.n8825 S.n8824 0.031
R43342 S.n7750 S.n7749 0.031
R43343 S.n6652 S.n6651 0.031
R43344 S.n5542 S.n5541 0.031
R43345 S.n4407 S.n4406 0.031
R43346 S.n3270 S.n3269 0.031
R43347 S.n2118 S.n2117 0.031
R43348 S.n2104 S.n2103 0.031
R43349 S.n3256 S.n3255 0.031
R43350 S.n4393 S.n4392 0.031
R43351 S.n5528 S.n5527 0.031
R43352 S.n6638 S.n6637 0.031
R43353 S.n7736 S.n7735 0.031
R43354 S.n8811 S.n8810 0.031
R43355 S.n9874 S.n9873 0.031
R43356 S.n10914 S.n10913 0.031
R43357 S.n11942 S.n11941 0.031
R43358 S.n12947 S.n12946 0.031
R43359 S.n13940 S.n13939 0.031
R43360 S.n14910 S.n14909 0.031
R43361 S.n15868 S.n15867 0.031
R43362 S.n16803 S.n16802 0.031
R43363 S.n17730 S.n17729 0.031
R43364 S.n18630 S.n18629 0.031
R43365 S.n15947 S.n15946 0.031
R43366 S.n14985 S.n14984 0.031
R43367 S.n14015 S.n14014 0.031
R43368 S.n13022 S.n13021 0.031
R43369 S.n12017 S.n12016 0.031
R43370 S.n10989 S.n10988 0.031
R43371 S.n9949 S.n9948 0.031
R43372 S.n8886 S.n8885 0.031
R43373 S.n7811 S.n7810 0.031
R43374 S.n6713 S.n6712 0.031
R43375 S.n5603 S.n5602 0.031
R43376 S.n4468 S.n4467 0.031
R43377 S.n3330 S.n3329 0.031
R43378 S.n2177 S.n2176 0.031
R43379 S.n2163 S.n2162 0.031
R43380 S.n3316 S.n3315 0.031
R43381 S.n4454 S.n4453 0.031
R43382 S.n5589 S.n5588 0.031
R43383 S.n6699 S.n6698 0.031
R43384 S.n7797 S.n7796 0.031
R43385 S.n8872 S.n8871 0.031
R43386 S.n9935 S.n9934 0.031
R43387 S.n10975 S.n10974 0.031
R43388 S.n12003 S.n12002 0.031
R43389 S.n13008 S.n13007 0.031
R43390 S.n14001 S.n14000 0.031
R43391 S.n14971 S.n14970 0.031
R43392 S.n15933 S.n15932 0.031
R43393 S.n16868 S.n16867 0.031
R43394 S.n14080 S.n14079 0.031
R43395 S.n13083 S.n13082 0.031
R43396 S.n12078 S.n12077 0.031
R43397 S.n11050 S.n11049 0.031
R43398 S.n10010 S.n10009 0.031
R43399 S.n8947 S.n8946 0.031
R43400 S.n7872 S.n7871 0.031
R43401 S.n6774 S.n6773 0.031
R43402 S.n5664 S.n5663 0.031
R43403 S.n4529 S.n4528 0.031
R43404 S.n3390 S.n3389 0.031
R43405 S.n2236 S.n2235 0.031
R43406 S.n2222 S.n2221 0.031
R43407 S.n3376 S.n3375 0.031
R43408 S.n4515 S.n4514 0.031
R43409 S.n5650 S.n5649 0.031
R43410 S.n6760 S.n6759 0.031
R43411 S.n7858 S.n7857 0.031
R43412 S.n8933 S.n8932 0.031
R43413 S.n9996 S.n9995 0.031
R43414 S.n11036 S.n11035 0.031
R43415 S.n12064 S.n12063 0.031
R43416 S.n13069 S.n13068 0.031
R43417 S.n14066 S.n14065 0.031
R43418 S.n15036 S.n15035 0.031
R43419 S.n12143 S.n12142 0.031
R43420 S.n11111 S.n11110 0.031
R43421 S.n10071 S.n10070 0.031
R43422 S.n9008 S.n9007 0.031
R43423 S.n7933 S.n7932 0.031
R43424 S.n6835 S.n6834 0.031
R43425 S.n5725 S.n5724 0.031
R43426 S.n4590 S.n4589 0.031
R43427 S.n3450 S.n3449 0.031
R43428 S.n2295 S.n2294 0.031
R43429 S.n2281 S.n2280 0.031
R43430 S.n3436 S.n3435 0.031
R43431 S.n4576 S.n4575 0.031
R43432 S.n5711 S.n5710 0.031
R43433 S.n6821 S.n6820 0.031
R43434 S.n7919 S.n7918 0.031
R43435 S.n8994 S.n8993 0.031
R43436 S.n10057 S.n10056 0.031
R43437 S.n11097 S.n11096 0.031
R43438 S.n12129 S.n12128 0.031
R43439 S.n13134 S.n13133 0.031
R43440 S.n10136 S.n10135 0.031
R43441 S.n9069 S.n9068 0.031
R43442 S.n7994 S.n7993 0.031
R43443 S.n6896 S.n6895 0.031
R43444 S.n5786 S.n5785 0.031
R43445 S.n4651 S.n4650 0.031
R43446 S.n3510 S.n3509 0.031
R43447 S.n2354 S.n2353 0.031
R43448 S.n2340 S.n2339 0.031
R43449 S.n3496 S.n3495 0.031
R43450 S.n4637 S.n4636 0.031
R43451 S.n5772 S.n5771 0.031
R43452 S.n6882 S.n6881 0.031
R43453 S.n7980 S.n7979 0.031
R43454 S.n9055 S.n9054 0.031
R43455 S.n10122 S.n10121 0.031
R43456 S.n11162 S.n11161 0.031
R43457 S.n8059 S.n8058 0.031
R43458 S.n6957 S.n6956 0.031
R43459 S.n5847 S.n5846 0.031
R43460 S.n4712 S.n4711 0.031
R43461 S.n3570 S.n3569 0.031
R43462 S.n2413 S.n2412 0.031
R43463 S.n2399 S.n2398 0.031
R43464 S.n3556 S.n3555 0.031
R43465 S.n4698 S.n4697 0.031
R43466 S.n5833 S.n5832 0.031
R43467 S.n6943 S.n6942 0.031
R43468 S.n8045 S.n8044 0.031
R43469 S.n9120 S.n9119 0.031
R43470 S.n5912 S.n5911 0.031
R43471 S.n4773 S.n4772 0.031
R43472 S.n3630 S.n3629 0.031
R43473 S.n2472 S.n2471 0.031
R43474 S.n2458 S.n2457 0.031
R43475 S.n3616 S.n3615 0.031
R43476 S.n4759 S.n4758 0.031
R43477 S.n5898 S.n5897 0.031
R43478 S.n7008 S.n7007 0.031
R43479 S.n3694 S.n3693 0.031
R43480 S.n2531 S.n2530 0.031
R43481 S.n2517 S.n2516 0.031
R43482 S.n3680 S.n3679 0.031
R43483 S.n4824 S.n4823 0.031
R43484 S.n2580 S.n2579 0.031
R43485 S.n22333 S.n22317 0.031
R43486 S.n23033 S.n23032 0.031
R43487 S.n23032 S.n23031 0.031
R43488 S.n23031 S.n23030 0.031
R43489 S.n23030 S.n23029 0.031
R43490 S.n23029 S.n23028 0.031
R43491 S.n23028 S.n23027 0.031
R43492 S.n23027 S.n23026 0.031
R43493 S.n23026 S.n23025 0.031
R43494 S.n23025 S.n23024 0.031
R43495 S.n23024 S.n23023 0.031
R43496 S.n23023 S.n23022 0.031
R43497 S.n23022 S.n23021 0.031
R43498 S.n23021 S.n23020 0.031
R43499 S.n23020 S.n23019 0.031
R43500 S.n23019 S.n23018 0.031
R43501 S.n23018 S.n23017 0.031
R43502 S.n23017 S.n23016 0.031
R43503 S.n23016 S.n23015 0.031
R43504 S.n23015 S.n23014 0.031
R43505 S.n23014 S.n23013 0.031
R43506 S.n23013 S.n23012 0.031
R43507 S.n23012 S.n23011 0.031
R43508 S.n1435 S.n1434 0.031
R43509 S.n1436 S.n1435 0.031
R43510 S.n1437 S.n1436 0.031
R43511 S.n1438 S.n1437 0.031
R43512 S.n1439 S.n1438 0.031
R43513 S.n1440 S.n1439 0.031
R43514 S.n1441 S.n1440 0.031
R43515 S.n22317 S.n22316 0.031
R43516 S.n15723 S.n15722 0.031
R43517 S.n13795 S.n13794 0.031
R43518 S.n11797 S.n11796 0.031
R43519 S.n19353 S.n19352 0.03
R43520 S.n17566 S.n17565 0.03
R43521 S.n15708 S.n15707 0.03
R43522 S.n13780 S.n13779 0.03
R43523 S.n11782 S.n11781 0.03
R43524 S.n9714 S.n9713 0.03
R43525 S.n7576 S.n7575 0.03
R43526 S.n5367 S.n5366 0.03
R43527 S.n3097 S.n3096 0.03
R43528 S.n20322 S.n20321 0.03
R43529 S.n19450 S.n19449 0.03
R43530 S.n18562 S.n18561 0.03
R43531 S.n17662 S.n17661 0.03
R43532 S.n16739 S.n16738 0.03
R43533 S.n15804 S.n15803 0.03
R43534 S.n14846 S.n14845 0.03
R43535 S.n13876 S.n13875 0.03
R43536 S.n12883 S.n12882 0.03
R43537 S.n11878 S.n11877 0.03
R43538 S.n10850 S.n10849 0.03
R43539 S.n9810 S.n9809 0.03
R43540 S.n8747 S.n8746 0.03
R43541 S.n7672 S.n7671 0.03
R43542 S.n6574 S.n6573 0.03
R43543 S.n5464 S.n5463 0.03
R43544 S.n4329 S.n4328 0.03
R43545 S.n3192 S.n3191 0.03
R43546 S.n2024 S.n2023 0.03
R43547 S.n1347 S.n1346 0.03
R43548 S.n1432 S.n1429 0.029
R43549 S.n18476 S.n18473 0.029
R43550 S.n20231 S.n20228 0.029
R43551 S.n16653 S.n16650 0.029
R43552 S.n14760 S.n14757 0.029
R43553 S.n12797 S.n12794 0.029
R43554 S.n10764 S.n10761 0.029
R43555 S.n8661 S.n8658 0.029
R43556 S.n6488 S.n6485 0.029
R43557 S.n4243 S.n4240 0.029
R43558 S.n3142 S.n3141 0.029
R43559 S.n4279 S.n4278 0.029
R43560 S.n5413 S.n5412 0.029
R43561 S.n6524 S.n6523 0.029
R43562 S.n7622 S.n7621 0.029
R43563 S.n8697 S.n8696 0.029
R43564 S.n9760 S.n9759 0.029
R43565 S.n10800 S.n10799 0.029
R43566 S.n11828 S.n11827 0.029
R43567 S.n12833 S.n12832 0.029
R43568 S.n13826 S.n13825 0.029
R43569 S.n14796 S.n14795 0.029
R43570 S.n15754 S.n15753 0.029
R43571 S.n16689 S.n16688 0.029
R43572 S.n17612 S.n17611 0.029
R43573 S.n18512 S.n18511 0.029
R43574 S.n19399 S.n19398 0.029
R43575 S.n20267 S.n20266 0.029
R43576 S.n3226 S.n3225 0.029
R43577 S.n4363 S.n4362 0.029
R43578 S.n5498 S.n5497 0.029
R43579 S.n6608 S.n6607 0.029
R43580 S.n7706 S.n7705 0.029
R43581 S.n8781 S.n8780 0.029
R43582 S.n9844 S.n9843 0.029
R43583 S.n10884 S.n10883 0.029
R43584 S.n11912 S.n11911 0.029
R43585 S.n12917 S.n12916 0.029
R43586 S.n13910 S.n13909 0.029
R43587 S.n14880 S.n14879 0.029
R43588 S.n15838 S.n15837 0.029
R43589 S.n16773 S.n16772 0.029
R43590 S.n17696 S.n17695 0.029
R43591 S.n3286 S.n3285 0.029
R43592 S.n4424 S.n4423 0.029
R43593 S.n5559 S.n5558 0.029
R43594 S.n6669 S.n6668 0.029
R43595 S.n7767 S.n7766 0.029
R43596 S.n8842 S.n8841 0.029
R43597 S.n9905 S.n9904 0.029
R43598 S.n10945 S.n10944 0.029
R43599 S.n11973 S.n11972 0.029
R43600 S.n12978 S.n12977 0.029
R43601 S.n13971 S.n13970 0.029
R43602 S.n14941 S.n14940 0.029
R43603 S.n15899 S.n15898 0.029
R43604 S.n3346 S.n3345 0.029
R43605 S.n4485 S.n4484 0.029
R43606 S.n5620 S.n5619 0.029
R43607 S.n6730 S.n6729 0.029
R43608 S.n7828 S.n7827 0.029
R43609 S.n8903 S.n8902 0.029
R43610 S.n9966 S.n9965 0.029
R43611 S.n11006 S.n11005 0.029
R43612 S.n12034 S.n12033 0.029
R43613 S.n13039 S.n13038 0.029
R43614 S.n14032 S.n14031 0.029
R43615 S.n3406 S.n3405 0.029
R43616 S.n4546 S.n4545 0.029
R43617 S.n5681 S.n5680 0.029
R43618 S.n6791 S.n6790 0.029
R43619 S.n7889 S.n7888 0.029
R43620 S.n8964 S.n8963 0.029
R43621 S.n10027 S.n10026 0.029
R43622 S.n11067 S.n11066 0.029
R43623 S.n12095 S.n12094 0.029
R43624 S.n3466 S.n3465 0.029
R43625 S.n4607 S.n4606 0.029
R43626 S.n5742 S.n5741 0.029
R43627 S.n6852 S.n6851 0.029
R43628 S.n7950 S.n7949 0.029
R43629 S.n9025 S.n9024 0.029
R43630 S.n10088 S.n10087 0.029
R43631 S.n3526 S.n3525 0.029
R43632 S.n4668 S.n4667 0.029
R43633 S.n5803 S.n5802 0.029
R43634 S.n6913 S.n6912 0.029
R43635 S.n8011 S.n8010 0.029
R43636 S.n3586 S.n3585 0.029
R43637 S.n4729 S.n4728 0.029
R43638 S.n5864 S.n5863 0.029
R43639 S.n3646 S.n3645 0.029
R43640 S.n18561 S.n18560 0.029
R43641 S.n17661 S.n17660 0.029
R43642 S.n16738 S.n16737 0.029
R43643 S.n15803 S.n15802 0.029
R43644 S.n14845 S.n14844 0.029
R43645 S.n13875 S.n13874 0.029
R43646 S.n12882 S.n12881 0.029
R43647 S.n11877 S.n11876 0.029
R43648 S.n10849 S.n10848 0.029
R43649 S.n9809 S.n9808 0.029
R43650 S.n8746 S.n8745 0.029
R43651 S.n7671 S.n7670 0.029
R43652 S.n6573 S.n6572 0.029
R43653 S.n5463 S.n5462 0.029
R43654 S.n4328 S.n4327 0.029
R43655 S.n3191 S.n3190 0.029
R43656 S.n2023 S.n2022 0.029
R43657 S.n1346 S.n1345 0.029
R43658 S.n21126 S.n21125 0.029
R43659 S.n19475 S.n19474 0.028
R43660 S.n18585 S.n18584 0.028
R43661 S.n17685 S.n17684 0.028
R43662 S.n16762 S.n16761 0.028
R43663 S.n15827 S.n15826 0.028
R43664 S.n14869 S.n14868 0.028
R43665 S.n13899 S.n13898 0.028
R43666 S.n12906 S.n12905 0.028
R43667 S.n11901 S.n11900 0.028
R43668 S.n10873 S.n10872 0.028
R43669 S.n9833 S.n9832 0.028
R43670 S.n8770 S.n8769 0.028
R43671 S.n7695 S.n7694 0.028
R43672 S.n6597 S.n6596 0.028
R43673 S.n5487 S.n5486 0.028
R43674 S.n4352 S.n4351 0.028
R43675 S.n21196 S.n21193 0.028
R43676 S.n20377 S.n20374 0.028
R43677 S.n20250 S.n20247 0.028
R43678 S.n19382 S.n19379 0.028
R43679 S.n18495 S.n18492 0.028
R43680 S.n17595 S.n17592 0.028
R43681 S.n16672 S.n16669 0.028
R43682 S.n15737 S.n15734 0.028
R43683 S.n14779 S.n14776 0.028
R43684 S.n13809 S.n13806 0.028
R43685 S.n12816 S.n12813 0.028
R43686 S.n11811 S.n11808 0.028
R43687 S.n10783 S.n10780 0.028
R43688 S.n9743 S.n9740 0.028
R43689 S.n8680 S.n8677 0.028
R43690 S.n7605 S.n7602 0.028
R43691 S.n6507 S.n6504 0.028
R43692 S.n5396 S.n5393 0.028
R43693 S.n4262 S.n4259 0.028
R43694 S.n3126 S.n3123 0.028
R43695 S.n1966 S.n1963 0.028
R43696 S.n17744 S.n17741 0.028
R43697 S.n16817 S.n16814 0.028
R43698 S.n15882 S.n15879 0.028
R43699 S.n14924 S.n14921 0.028
R43700 S.n13954 S.n13951 0.028
R43701 S.n12961 S.n12958 0.028
R43702 S.n11956 S.n11953 0.028
R43703 S.n10928 S.n10925 0.028
R43704 S.n9888 S.n9885 0.028
R43705 S.n8825 S.n8822 0.028
R43706 S.n7750 S.n7747 0.028
R43707 S.n6652 S.n6649 0.028
R43708 S.n5542 S.n5539 0.028
R43709 S.n4407 S.n4404 0.028
R43710 S.n3270 S.n3267 0.028
R43711 S.n2118 S.n2115 0.028
R43712 S.n3256 S.n3253 0.028
R43713 S.n4393 S.n4390 0.028
R43714 S.n5528 S.n5525 0.028
R43715 S.n6638 S.n6635 0.028
R43716 S.n7736 S.n7733 0.028
R43717 S.n8811 S.n8808 0.028
R43718 S.n9874 S.n9871 0.028
R43719 S.n10914 S.n10911 0.028
R43720 S.n11942 S.n11939 0.028
R43721 S.n12947 S.n12944 0.028
R43722 S.n13940 S.n13937 0.028
R43723 S.n14910 S.n14907 0.028
R43724 S.n15868 S.n15865 0.028
R43725 S.n16803 S.n16800 0.028
R43726 S.n17730 S.n17727 0.028
R43727 S.n18630 S.n18627 0.028
R43728 S.n15947 S.n15944 0.028
R43729 S.n14985 S.n14982 0.028
R43730 S.n14015 S.n14012 0.028
R43731 S.n13022 S.n13019 0.028
R43732 S.n12017 S.n12014 0.028
R43733 S.n10989 S.n10986 0.028
R43734 S.n9949 S.n9946 0.028
R43735 S.n8886 S.n8883 0.028
R43736 S.n7811 S.n7808 0.028
R43737 S.n6713 S.n6710 0.028
R43738 S.n5603 S.n5600 0.028
R43739 S.n4468 S.n4465 0.028
R43740 S.n3330 S.n3327 0.028
R43741 S.n2177 S.n2174 0.028
R43742 S.n2163 S.n2160 0.028
R43743 S.n3316 S.n3313 0.028
R43744 S.n4454 S.n4451 0.028
R43745 S.n5589 S.n5586 0.028
R43746 S.n6699 S.n6696 0.028
R43747 S.n7797 S.n7794 0.028
R43748 S.n8872 S.n8869 0.028
R43749 S.n9935 S.n9932 0.028
R43750 S.n10975 S.n10972 0.028
R43751 S.n12003 S.n12000 0.028
R43752 S.n13008 S.n13005 0.028
R43753 S.n14001 S.n13998 0.028
R43754 S.n14971 S.n14968 0.028
R43755 S.n15933 S.n15930 0.028
R43756 S.n16868 S.n16865 0.028
R43757 S.n14080 S.n14077 0.028
R43758 S.n13083 S.n13080 0.028
R43759 S.n12078 S.n12075 0.028
R43760 S.n11050 S.n11047 0.028
R43761 S.n10010 S.n10007 0.028
R43762 S.n8947 S.n8944 0.028
R43763 S.n7872 S.n7869 0.028
R43764 S.n6774 S.n6771 0.028
R43765 S.n5664 S.n5661 0.028
R43766 S.n4529 S.n4526 0.028
R43767 S.n3390 S.n3387 0.028
R43768 S.n2236 S.n2233 0.028
R43769 S.n2222 S.n2219 0.028
R43770 S.n3376 S.n3373 0.028
R43771 S.n4515 S.n4512 0.028
R43772 S.n5650 S.n5647 0.028
R43773 S.n6760 S.n6757 0.028
R43774 S.n7858 S.n7855 0.028
R43775 S.n8933 S.n8930 0.028
R43776 S.n9996 S.n9993 0.028
R43777 S.n11036 S.n11033 0.028
R43778 S.n12064 S.n12061 0.028
R43779 S.n13069 S.n13066 0.028
R43780 S.n14066 S.n14063 0.028
R43781 S.n15036 S.n15033 0.028
R43782 S.n12143 S.n12140 0.028
R43783 S.n11111 S.n11108 0.028
R43784 S.n10071 S.n10068 0.028
R43785 S.n9008 S.n9005 0.028
R43786 S.n7933 S.n7930 0.028
R43787 S.n6835 S.n6832 0.028
R43788 S.n5725 S.n5722 0.028
R43789 S.n4590 S.n4587 0.028
R43790 S.n3450 S.n3447 0.028
R43791 S.n2295 S.n2292 0.028
R43792 S.n2281 S.n2278 0.028
R43793 S.n3436 S.n3433 0.028
R43794 S.n4576 S.n4573 0.028
R43795 S.n5711 S.n5708 0.028
R43796 S.n6821 S.n6818 0.028
R43797 S.n7919 S.n7916 0.028
R43798 S.n8994 S.n8991 0.028
R43799 S.n10057 S.n10054 0.028
R43800 S.n11097 S.n11094 0.028
R43801 S.n12129 S.n12126 0.028
R43802 S.n13134 S.n13131 0.028
R43803 S.n10136 S.n10133 0.028
R43804 S.n9069 S.n9066 0.028
R43805 S.n7994 S.n7991 0.028
R43806 S.n6896 S.n6893 0.028
R43807 S.n5786 S.n5783 0.028
R43808 S.n4651 S.n4648 0.028
R43809 S.n3510 S.n3507 0.028
R43810 S.n2354 S.n2351 0.028
R43811 S.n2340 S.n2337 0.028
R43812 S.n3496 S.n3493 0.028
R43813 S.n4637 S.n4634 0.028
R43814 S.n5772 S.n5769 0.028
R43815 S.n6882 S.n6879 0.028
R43816 S.n7980 S.n7977 0.028
R43817 S.n9055 S.n9052 0.028
R43818 S.n10122 S.n10119 0.028
R43819 S.n11162 S.n11159 0.028
R43820 S.n8059 S.n8056 0.028
R43821 S.n6957 S.n6954 0.028
R43822 S.n5847 S.n5844 0.028
R43823 S.n4712 S.n4709 0.028
R43824 S.n3570 S.n3567 0.028
R43825 S.n2413 S.n2410 0.028
R43826 S.n2399 S.n2396 0.028
R43827 S.n3556 S.n3553 0.028
R43828 S.n4698 S.n4695 0.028
R43829 S.n5833 S.n5830 0.028
R43830 S.n6943 S.n6940 0.028
R43831 S.n8045 S.n8042 0.028
R43832 S.n9120 S.n9117 0.028
R43833 S.n5912 S.n5909 0.028
R43834 S.n4773 S.n4770 0.028
R43835 S.n3630 S.n3627 0.028
R43836 S.n2472 S.n2469 0.028
R43837 S.n2458 S.n2455 0.028
R43838 S.n3616 S.n3613 0.028
R43839 S.n4759 S.n4756 0.028
R43840 S.n5898 S.n5895 0.028
R43841 S.n7008 S.n7005 0.028
R43842 S.n3694 S.n3691 0.028
R43843 S.n2531 S.n2528 0.028
R43844 S.n2517 S.n2514 0.028
R43845 S.n3680 S.n3677 0.028
R43846 S.n4824 S.n4821 0.028
R43847 S.n2580 S.n2577 0.028
R43848 S.n1927 S.n1926 0.028
R43849 S.n1929 S.n1927 0.028
R43850 S.n2039 S.n2038 0.028
R43851 S.n1813 S.n1812 0.028
R43852 S.n3179 S.n3178 0.028
R43853 S.n2976 S.n2975 0.028
R43854 S.n4316 S.n4315 0.028
R43855 S.n4103 S.n4102 0.028
R43856 S.n5451 S.n5450 0.028
R43857 S.n5215 S.n5214 0.028
R43858 S.n6561 S.n6560 0.028
R43859 S.n6315 S.n6314 0.028
R43860 S.n7659 S.n7658 0.028
R43861 S.n7392 S.n7391 0.028
R43862 S.n8734 S.n8733 0.028
R43863 S.n8456 S.n8455 0.028
R43864 S.n9797 S.n9796 0.028
R43865 S.n9498 S.n9497 0.028
R43866 S.n10837 S.n10836 0.028
R43867 S.n10527 S.n10526 0.028
R43868 S.n11865 S.n11864 0.028
R43869 S.n11534 S.n11533 0.028
R43870 S.n12870 S.n12869 0.028
R43871 S.n12528 S.n12527 0.028
R43872 S.n13863 S.n13862 0.028
R43873 S.n13500 S.n13499 0.028
R43874 S.n14833 S.n14832 0.028
R43875 S.n14459 S.n14458 0.028
R43876 S.n15791 S.n15790 0.028
R43877 S.n15396 S.n15395 0.028
R43878 S.n16726 S.n16725 0.028
R43879 S.n16320 S.n16319 0.028
R43880 S.n17649 S.n17648 0.028
R43881 S.n17222 S.n17221 0.028
R43882 S.n18549 S.n18548 0.028
R43883 S.n18111 S.n18110 0.028
R43884 S.n19436 S.n19435 0.028
R43885 S.n18976 S.n18975 0.028
R43886 S.n20308 S.n20307 0.028
R43887 S.n19828 S.n19827 0.028
R43888 S.n20412 S.n20411 0.028
R43889 S.n761 S.n760 0.028
R43890 S.n2006 S.n2005 0.028
R43891 S.n2008 S.n2006 0.028
R43892 S.n20394 S.n20393 0.028
R43893 S.n21213 S.n21212 0.028
R43894 S.n22734 S.n22733 0.028
R43895 S.n18596 S.n18595 0.028
R43896 S.n19486 S.n19485 0.028
R43897 S.n20231 S.n20230 0.028
R43898 S.n16834 S.n16833 0.028
R43899 S.n17761 S.n17760 0.028
R43900 S.n18476 S.n18475 0.028
R43901 S.n15002 S.n15001 0.028
R43902 S.n15964 S.n15963 0.028
R43903 S.n16653 S.n16652 0.028
R43904 S.n13100 S.n13099 0.028
R43905 S.n14097 S.n14096 0.028
R43906 S.n14760 S.n14759 0.028
R43907 S.n11128 S.n11127 0.028
R43908 S.n12160 S.n12159 0.028
R43909 S.n12797 S.n12796 0.028
R43910 S.n9086 S.n9085 0.028
R43911 S.n10153 S.n10152 0.028
R43912 S.n10764 S.n10763 0.028
R43913 S.n6974 S.n6973 0.028
R43914 S.n8076 S.n8075 0.028
R43915 S.n8661 S.n8660 0.028
R43916 S.n4790 S.n4789 0.028
R43917 S.n5929 S.n5928 0.028
R43918 S.n6488 S.n6487 0.028
R43919 S.n3710 S.n3709 0.028
R43920 S.n4243 S.n4242 0.028
R43921 S.n1812 S.n1811 0.028
R43922 S.n2975 S.n2974 0.028
R43923 S.n4102 S.n4101 0.028
R43924 S.n5214 S.n5213 0.028
R43925 S.n6314 S.n6313 0.028
R43926 S.n7391 S.n7390 0.028
R43927 S.n8455 S.n8454 0.028
R43928 S.n9497 S.n9496 0.028
R43929 S.n10526 S.n10525 0.028
R43930 S.n11533 S.n11532 0.028
R43931 S.n12527 S.n12526 0.028
R43932 S.n13499 S.n13498 0.028
R43933 S.n14458 S.n14457 0.028
R43934 S.n15395 S.n15394 0.028
R43935 S.n16319 S.n16318 0.028
R43936 S.n17221 S.n17220 0.028
R43937 S.n18110 S.n18109 0.028
R43938 S.n18975 S.n18974 0.028
R43939 S.n19827 S.n19826 0.028
R43940 S.n760 S.n759 0.028
R43941 S.n21986 S.n21984 0.027
R43942 S.n21952 S.n21950 0.027
R43943 S.n22674 S.n22673 0.027
R43944 S.n22367 S.n22366 0.027
R43945 S.n22342 S.n22341 0.027
R43946 S.n3216 S.n3215 0.027
R43947 S.n2597 S.n1902 0.027
R43948 S.n860 S.n859 0.027
R43949 S.n19366 S.n19365 0.027
R43950 S.n17579 S.n17578 0.027
R43951 S.n15722 S.n15721 0.027
R43952 S.n13794 S.n13793 0.027
R43953 S.n11796 S.n11795 0.027
R43954 S.n9727 S.n9726 0.027
R43955 S.n7589 S.n7588 0.027
R43956 S.n5380 S.n5379 0.027
R43957 S.n3110 S.n3109 0.027
R43958 S.n21980 S.n21979 0.027
R43959 S.n1774 S.n1773 0.027
R43960 S.n21172 S.n20346 0.026
R43961 S.n20344 S.n19524 0.026
R43962 S.n19504 S.n18667 0.026
R43963 S.n18647 S.n17799 0.026
R43964 S.n17779 S.n16905 0.026
R43965 S.n16885 S.n16002 0.026
R43966 S.n15982 S.n15073 0.026
R43967 S.n15053 S.n14135 0.026
R43968 S.n14115 S.n13171 0.026
R43969 S.n13151 S.n12198 0.026
R43970 S.n12178 S.n11199 0.026
R43971 S.n11179 S.n10191 0.026
R43972 S.n10171 S.n9157 0.026
R43973 S.n9137 S.n8114 0.026
R43974 S.n8094 S.n7045 0.026
R43975 S.n7025 S.n5967 0.026
R43976 S.n5947 S.n4862 0.026
R43977 S.n4841 S.n3749 0.026
R43978 S.n1985 S.n1982 0.026
R43979 S.n1865 S.n1862 0.026
R43980 S.n3146 S.n3143 0.026
R43981 S.n3025 S.n3022 0.026
R43982 S.n4283 S.n4280 0.026
R43983 S.n4151 S.n4148 0.026
R43984 S.n5417 S.n5414 0.026
R43985 S.n5264 S.n5261 0.026
R43986 S.n6528 S.n6525 0.026
R43987 S.n6364 S.n6361 0.026
R43988 S.n7626 S.n7623 0.026
R43989 S.n7441 S.n7438 0.026
R43990 S.n8701 S.n8698 0.026
R43991 S.n8505 S.n8502 0.026
R43992 S.n9764 S.n9761 0.026
R43993 S.n9547 S.n9544 0.026
R43994 S.n10804 S.n10801 0.026
R43995 S.n10576 S.n10573 0.026
R43996 S.n11832 S.n11829 0.026
R43997 S.n11583 S.n11580 0.026
R43998 S.n12837 S.n12834 0.026
R43999 S.n12577 S.n12574 0.026
R44000 S.n13830 S.n13827 0.026
R44001 S.n13549 S.n13546 0.026
R44002 S.n14800 S.n14797 0.026
R44003 S.n14508 S.n14505 0.026
R44004 S.n15758 S.n15755 0.026
R44005 S.n15445 S.n15442 0.026
R44006 S.n16693 S.n16690 0.026
R44007 S.n16369 S.n16366 0.026
R44008 S.n17616 S.n17613 0.026
R44009 S.n17271 S.n17268 0.026
R44010 S.n18516 S.n18513 0.026
R44011 S.n18160 S.n18157 0.026
R44012 S.n19403 S.n19400 0.026
R44013 S.n19026 S.n19023 0.026
R44014 S.n20271 S.n20268 0.026
R44015 S.n19880 S.n19877 0.026
R44016 S.n20398 S.n20395 0.026
R44017 S.n20491 S.n20488 0.026
R44018 S.n21217 S.n21214 0.026
R44019 S.n21314 S.n21311 0.026
R44020 S.n22741 S.n22735 0.026
R44021 S.n2079 S.n2057 0.026
R44022 S.n1799 S.n1787 0.026
R44023 S.n3230 S.n3227 0.026
R44024 S.n2961 S.n2958 0.026
R44025 S.n4367 S.n4364 0.026
R44026 S.n4088 S.n4085 0.026
R44027 S.n5502 S.n5499 0.026
R44028 S.n5200 S.n5197 0.026
R44029 S.n6612 S.n6609 0.026
R44030 S.n6300 S.n6297 0.026
R44031 S.n7710 S.n7707 0.026
R44032 S.n7377 S.n7374 0.026
R44033 S.n8785 S.n8782 0.026
R44034 S.n8441 S.n8438 0.026
R44035 S.n9848 S.n9845 0.026
R44036 S.n9483 S.n9480 0.026
R44037 S.n10888 S.n10885 0.026
R44038 S.n10512 S.n10509 0.026
R44039 S.n11916 S.n11913 0.026
R44040 S.n11519 S.n11516 0.026
R44041 S.n12921 S.n12918 0.026
R44042 S.n12513 S.n12510 0.026
R44043 S.n13914 S.n13911 0.026
R44044 S.n13485 S.n13482 0.026
R44045 S.n14884 S.n14881 0.026
R44046 S.n14444 S.n14441 0.026
R44047 S.n15842 S.n15839 0.026
R44048 S.n15381 S.n15378 0.026
R44049 S.n16777 S.n16774 0.026
R44050 S.n16305 S.n16302 0.026
R44051 S.n17700 S.n17697 0.026
R44052 S.n17207 S.n17204 0.026
R44053 S.n18600 S.n18597 0.026
R44054 S.n18096 S.n18093 0.026
R44055 S.n19490 S.n19487 0.026
R44056 S.n18961 S.n18958 0.026
R44057 S.n20238 S.n20232 0.026
R44058 S.n1810 S.n1807 0.026
R44059 S.n2972 S.n2969 0.026
R44060 S.n4099 S.n4096 0.026
R44061 S.n5211 S.n5208 0.026
R44062 S.n6311 S.n6308 0.026
R44063 S.n7388 S.n7385 0.026
R44064 S.n8452 S.n8449 0.026
R44065 S.n9494 S.n9491 0.026
R44066 S.n10523 S.n10520 0.026
R44067 S.n11530 S.n11527 0.026
R44068 S.n12524 S.n12521 0.026
R44069 S.n13496 S.n13493 0.026
R44070 S.n14455 S.n14452 0.026
R44071 S.n15392 S.n15389 0.026
R44072 S.n16316 S.n16313 0.026
R44073 S.n17218 S.n17215 0.026
R44074 S.n18107 S.n18104 0.026
R44075 S.n18972 S.n18969 0.026
R44076 S.n19824 S.n19821 0.026
R44077 S.n20471 S.n20470 0.026
R44078 S.n19860 S.n19859 0.026
R44079 S.n19006 S.n19005 0.026
R44080 S.n18140 S.n18139 0.026
R44081 S.n17251 S.n17250 0.026
R44082 S.n16349 S.n16348 0.026
R44083 S.n15425 S.n15424 0.026
R44084 S.n14488 S.n14487 0.026
R44085 S.n13529 S.n13528 0.026
R44086 S.n12557 S.n12556 0.026
R44087 S.n11563 S.n11562 0.026
R44088 S.n10556 S.n10555 0.026
R44089 S.n9527 S.n9526 0.026
R44090 S.n8485 S.n8484 0.026
R44091 S.n7421 S.n7420 0.026
R44092 S.n6344 S.n6343 0.026
R44093 S.n5244 S.n5243 0.026
R44094 S.n4131 S.n4130 0.026
R44095 S.n3005 S.n3004 0.026
R44096 S.n1834 S.n1833 0.026
R44097 S.n2012 S.n1996 0.026
R44098 S.n3166 S.n3157 0.026
R44099 S.n4303 S.n4294 0.026
R44100 S.n5438 S.n5428 0.026
R44101 S.n6548 S.n6539 0.026
R44102 S.n7646 S.n7637 0.026
R44103 S.n8721 S.n8712 0.026
R44104 S.n9784 S.n9775 0.026
R44105 S.n10824 S.n10815 0.026
R44106 S.n11852 S.n11843 0.026
R44107 S.n12857 S.n12848 0.026
R44108 S.n13850 S.n13841 0.026
R44109 S.n14820 S.n14811 0.026
R44110 S.n15778 S.n15769 0.026
R44111 S.n16713 S.n16704 0.026
R44112 S.n17636 S.n17627 0.026
R44113 S.n18536 S.n18527 0.026
R44114 S.n19423 S.n19414 0.026
R44115 S.n20295 S.n20286 0.026
R44116 S.n20366 S.n20357 0.026
R44117 S.n21242 S.n21233 0.026
R44118 S.n864 S.n850 0.026
R44119 S.n19370 S.n19354 0.026
R44120 S.n18633 S.n18615 0.026
R44121 S.n17733 S.n17715 0.026
R44122 S.n16806 S.n16788 0.026
R44123 S.n15871 S.n15853 0.026
R44124 S.n14913 S.n14895 0.026
R44125 S.n13943 S.n13925 0.026
R44126 S.n12950 S.n12932 0.026
R44127 S.n11945 S.n11927 0.026
R44128 S.n10917 S.n10899 0.026
R44129 S.n9877 S.n9859 0.026
R44130 S.n8814 S.n8796 0.026
R44131 S.n7739 S.n7721 0.026
R44132 S.n6641 S.n6623 0.026
R44133 S.n5531 S.n5513 0.026
R44134 S.n4396 S.n4378 0.026
R44135 S.n3259 S.n3241 0.026
R44136 S.n2107 S.n2091 0.026
R44137 S.n24 S.n10 0.026
R44138 S.n2137 S.n2134 0.026
R44139 S.n1757 S.n1754 0.026
R44140 S.n3290 S.n3287 0.026
R44141 S.n2925 S.n2922 0.026
R44142 S.n4428 S.n4425 0.026
R44143 S.n4052 S.n4049 0.026
R44144 S.n5563 S.n5560 0.026
R44145 S.n5164 S.n5161 0.026
R44146 S.n6673 S.n6670 0.026
R44147 S.n6264 S.n6261 0.026
R44148 S.n7771 S.n7768 0.026
R44149 S.n7341 S.n7338 0.026
R44150 S.n8846 S.n8843 0.026
R44151 S.n8405 S.n8402 0.026
R44152 S.n9909 S.n9906 0.026
R44153 S.n9447 S.n9444 0.026
R44154 S.n10949 S.n10946 0.026
R44155 S.n10476 S.n10473 0.026
R44156 S.n11977 S.n11974 0.026
R44157 S.n11483 S.n11480 0.026
R44158 S.n12982 S.n12979 0.026
R44159 S.n12477 S.n12474 0.026
R44160 S.n13975 S.n13972 0.026
R44161 S.n13449 S.n13446 0.026
R44162 S.n14945 S.n14942 0.026
R44163 S.n14408 S.n14405 0.026
R44164 S.n15903 S.n15900 0.026
R44165 S.n15345 S.n15342 0.026
R44166 S.n16838 S.n16835 0.026
R44167 S.n16269 S.n16266 0.026
R44168 S.n17765 S.n17762 0.026
R44169 S.n17169 S.n17166 0.026
R44170 S.n18483 S.n18477 0.026
R44171 S.n17583 S.n17567 0.026
R44172 S.n16871 S.n16853 0.026
R44173 S.n15936 S.n15918 0.026
R44174 S.n14974 S.n14956 0.026
R44175 S.n14004 S.n13986 0.026
R44176 S.n13011 S.n12993 0.026
R44177 S.n12006 S.n11988 0.026
R44178 S.n10978 S.n10960 0.026
R44179 S.n9938 S.n9920 0.026
R44180 S.n8875 S.n8857 0.026
R44181 S.n7800 S.n7782 0.026
R44182 S.n6702 S.n6684 0.026
R44183 S.n5592 S.n5574 0.026
R44184 S.n4457 S.n4439 0.026
R44185 S.n3319 S.n3301 0.026
R44186 S.n2166 S.n2149 0.026
R44187 S.n71 S.n57 0.026
R44188 S.n2196 S.n2193 0.026
R44189 S.n1720 S.n1717 0.026
R44190 S.n3350 S.n3347 0.026
R44191 S.n2889 S.n2886 0.026
R44192 S.n4489 S.n4486 0.026
R44193 S.n4016 S.n4013 0.026
R44194 S.n5624 S.n5621 0.026
R44195 S.n5128 S.n5125 0.026
R44196 S.n6734 S.n6731 0.026
R44197 S.n6228 S.n6225 0.026
R44198 S.n7832 S.n7829 0.026
R44199 S.n7305 S.n7302 0.026
R44200 S.n8907 S.n8904 0.026
R44201 S.n8369 S.n8366 0.026
R44202 S.n9970 S.n9967 0.026
R44203 S.n9411 S.n9408 0.026
R44204 S.n11010 S.n11007 0.026
R44205 S.n10440 S.n10437 0.026
R44206 S.n12038 S.n12035 0.026
R44207 S.n11447 S.n11444 0.026
R44208 S.n13043 S.n13040 0.026
R44209 S.n12441 S.n12438 0.026
R44210 S.n14036 S.n14033 0.026
R44211 S.n13413 S.n13410 0.026
R44212 S.n15006 S.n15003 0.026
R44213 S.n14372 S.n14369 0.026
R44214 S.n15968 S.n15965 0.026
R44215 S.n15307 S.n15304 0.026
R44216 S.n16660 S.n16654 0.026
R44217 S.n15725 S.n15709 0.026
R44218 S.n15039 S.n15021 0.026
R44219 S.n14069 S.n14051 0.026
R44220 S.n13072 S.n13054 0.026
R44221 S.n12067 S.n12049 0.026
R44222 S.n11039 S.n11021 0.026
R44223 S.n9999 S.n9981 0.026
R44224 S.n8936 S.n8918 0.026
R44225 S.n7861 S.n7843 0.026
R44226 S.n6763 S.n6745 0.026
R44227 S.n5653 S.n5635 0.026
R44228 S.n4518 S.n4500 0.026
R44229 S.n3379 S.n3361 0.026
R44230 S.n2225 S.n2208 0.026
R44231 S.n103 S.n89 0.026
R44232 S.n2255 S.n2252 0.026
R44233 S.n1683 S.n1680 0.026
R44234 S.n3410 S.n3407 0.026
R44235 S.n2853 S.n2850 0.026
R44236 S.n4550 S.n4547 0.026
R44237 S.n3980 S.n3977 0.026
R44238 S.n5685 S.n5682 0.026
R44239 S.n5092 S.n5089 0.026
R44240 S.n6795 S.n6792 0.026
R44241 S.n6192 S.n6189 0.026
R44242 S.n7893 S.n7890 0.026
R44243 S.n7269 S.n7266 0.026
R44244 S.n8968 S.n8965 0.026
R44245 S.n8333 S.n8330 0.026
R44246 S.n10031 S.n10028 0.026
R44247 S.n9375 S.n9372 0.026
R44248 S.n11071 S.n11068 0.026
R44249 S.n10404 S.n10401 0.026
R44250 S.n12099 S.n12096 0.026
R44251 S.n11411 S.n11408 0.026
R44252 S.n13104 S.n13101 0.026
R44253 S.n12405 S.n12402 0.026
R44254 S.n14101 S.n14098 0.026
R44255 S.n13375 S.n13372 0.026
R44256 S.n14767 S.n14761 0.026
R44257 S.n13797 S.n13781 0.026
R44258 S.n13137 S.n13119 0.026
R44259 S.n12132 S.n12114 0.026
R44260 S.n11100 S.n11082 0.026
R44261 S.n10060 S.n10042 0.026
R44262 S.n8997 S.n8979 0.026
R44263 S.n7922 S.n7904 0.026
R44264 S.n6824 S.n6806 0.026
R44265 S.n5714 S.n5696 0.026
R44266 S.n4579 S.n4561 0.026
R44267 S.n3439 S.n3421 0.026
R44268 S.n2284 S.n2267 0.026
R44269 S.n990 S.n121 0.026
R44270 S.n2314 S.n2311 0.026
R44271 S.n1646 S.n1643 0.026
R44272 S.n3470 S.n3467 0.026
R44273 S.n2817 S.n2814 0.026
R44274 S.n4611 S.n4608 0.026
R44275 S.n3944 S.n3941 0.026
R44276 S.n5746 S.n5743 0.026
R44277 S.n5056 S.n5053 0.026
R44278 S.n6856 S.n6853 0.026
R44279 S.n6156 S.n6153 0.026
R44280 S.n7954 S.n7951 0.026
R44281 S.n7233 S.n7230 0.026
R44282 S.n9029 S.n9026 0.026
R44283 S.n8297 S.n8294 0.026
R44284 S.n10092 S.n10089 0.026
R44285 S.n9339 S.n9336 0.026
R44286 S.n11132 S.n11129 0.026
R44287 S.n10368 S.n10365 0.026
R44288 S.n12164 S.n12161 0.026
R44289 S.n11373 S.n11370 0.026
R44290 S.n12804 S.n12798 0.026
R44291 S.n11799 S.n11783 0.026
R44292 S.n11165 S.n11147 0.026
R44293 S.n10125 S.n10107 0.026
R44294 S.n9058 S.n9040 0.026
R44295 S.n7983 S.n7965 0.026
R44296 S.n6885 S.n6867 0.026
R44297 S.n5775 S.n5757 0.026
R44298 S.n4640 S.n4622 0.026
R44299 S.n3499 S.n3481 0.026
R44300 S.n2343 S.n2326 0.026
R44301 S.n1022 S.n1008 0.026
R44302 S.n2373 S.n2370 0.026
R44303 S.n1609 S.n1606 0.026
R44304 S.n3530 S.n3527 0.026
R44305 S.n2781 S.n2778 0.026
R44306 S.n4672 S.n4669 0.026
R44307 S.n3908 S.n3905 0.026
R44308 S.n5807 S.n5804 0.026
R44309 S.n5020 S.n5017 0.026
R44310 S.n6917 S.n6914 0.026
R44311 S.n6120 S.n6117 0.026
R44312 S.n8015 S.n8012 0.026
R44313 S.n7197 S.n7194 0.026
R44314 S.n9090 S.n9087 0.026
R44315 S.n8261 S.n8258 0.026
R44316 S.n10157 S.n10154 0.026
R44317 S.n9301 S.n9298 0.026
R44318 S.n10771 S.n10765 0.026
R44319 S.n9731 S.n9715 0.026
R44320 S.n9123 S.n9105 0.026
R44321 S.n8048 S.n8030 0.026
R44322 S.n6946 S.n6928 0.026
R44323 S.n5836 S.n5818 0.026
R44324 S.n4701 S.n4683 0.026
R44325 S.n3559 S.n3541 0.026
R44326 S.n2402 S.n2385 0.026
R44327 S.n1054 S.n1040 0.026
R44328 S.n2432 S.n2429 0.026
R44329 S.n1572 S.n1569 0.026
R44330 S.n3590 S.n3587 0.026
R44331 S.n2745 S.n2742 0.026
R44332 S.n4733 S.n4730 0.026
R44333 S.n3872 S.n3869 0.026
R44334 S.n5868 S.n5865 0.026
R44335 S.n4984 S.n4981 0.026
R44336 S.n6978 S.n6975 0.026
R44337 S.n6084 S.n6081 0.026
R44338 S.n8080 S.n8077 0.026
R44339 S.n7159 S.n7156 0.026
R44340 S.n8668 S.n8662 0.026
R44341 S.n7593 S.n7577 0.026
R44342 S.n7011 S.n6993 0.026
R44343 S.n5901 S.n5883 0.026
R44344 S.n4762 S.n4744 0.026
R44345 S.n3619 S.n3601 0.026
R44346 S.n2461 S.n2444 0.026
R44347 S.n1086 S.n1072 0.026
R44348 S.n2491 S.n2488 0.026
R44349 S.n1535 S.n1532 0.026
R44350 S.n3650 S.n3647 0.026
R44351 S.n2709 S.n2706 0.026
R44352 S.n4794 S.n4791 0.026
R44353 S.n3836 S.n3833 0.026
R44354 S.n5933 S.n5930 0.026
R44355 S.n4946 S.n4943 0.026
R44356 S.n6495 S.n6489 0.026
R44357 S.n5384 S.n5368 0.026
R44358 S.n4827 S.n4809 0.026
R44359 S.n3683 S.n3665 0.026
R44360 S.n2520 S.n2503 0.026
R44361 S.n1118 S.n1104 0.026
R44362 S.n2550 S.n2547 0.026
R44363 S.n1498 S.n1495 0.026
R44364 S.n3714 S.n3711 0.026
R44365 S.n2671 S.n2668 0.026
R44366 S.n4250 S.n4244 0.026
R44367 S.n1954 S.n1948 0.026
R44368 S.n3114 S.n3098 0.026
R44369 S.n2583 S.n2565 0.026
R44370 S.n1156 S.n1142 0.026
R44371 S.n942 S.n929 0.026
R44372 S.n942 S.n939 0.026
R44373 S.n22325 S.n22324 0.026
R44374 S.n928 S.n927 0.026
R44375 S.n838 S.n837 0.026
R44376 S.n902 S.n901 0.026
R44377 S.n22751 S.n22750 0.025
R44378 S.n19474 S.n19469 0.025
R44379 S.n18584 S.n18579 0.025
R44380 S.n17684 S.n17679 0.025
R44381 S.n16761 S.n16756 0.025
R44382 S.n15826 S.n15821 0.025
R44383 S.n14868 S.n14863 0.025
R44384 S.n13898 S.n13893 0.025
R44385 S.n12905 S.n12900 0.025
R44386 S.n11900 S.n11895 0.025
R44387 S.n10872 S.n10867 0.025
R44388 S.n9832 S.n9827 0.025
R44389 S.n8769 S.n8764 0.025
R44390 S.n7694 S.n7689 0.025
R44391 S.n6596 S.n6591 0.025
R44392 S.n5486 S.n5481 0.025
R44393 S.n4351 S.n4346 0.025
R44394 S.n3215 S.n3210 0.025
R44395 S.n3198 S.n3176 0.025
R44396 S.n4335 S.n4313 0.025
R44397 S.n5470 S.n5448 0.025
R44398 S.n6580 S.n6558 0.025
R44399 S.n7678 S.n7656 0.025
R44400 S.n8753 S.n8731 0.025
R44401 S.n9816 S.n9794 0.025
R44402 S.n10856 S.n10834 0.025
R44403 S.n11884 S.n11862 0.025
R44404 S.n12889 S.n12867 0.025
R44405 S.n13882 S.n13860 0.025
R44406 S.n14852 S.n14830 0.025
R44407 S.n15810 S.n15788 0.025
R44408 S.n16745 S.n16723 0.025
R44409 S.n17668 S.n17646 0.025
R44410 S.n18568 S.n18546 0.025
R44411 S.n19458 S.n19433 0.025
R44412 S.n20330 S.n20305 0.025
R44413 S.n20424 S.n20409 0.025
R44414 S.n2045 S.n2044 0.025
R44415 S.n2073 S.n2072 0.025
R44416 S.n19524 S.n19523 0.025
R44417 S.n18667 S.n18666 0.025
R44418 S.n17799 S.n17798 0.025
R44419 S.n16905 S.n16904 0.025
R44420 S.n16002 S.n16001 0.025
R44421 S.n15073 S.n15072 0.025
R44422 S.n14135 S.n14134 0.025
R44423 S.n13171 S.n13170 0.025
R44424 S.n12198 S.n12197 0.025
R44425 S.n11199 S.n11198 0.025
R44426 S.n10191 S.n10190 0.025
R44427 S.n9157 S.n9156 0.025
R44428 S.n8114 S.n8113 0.025
R44429 S.n7045 S.n7044 0.025
R44430 S.n5967 S.n5966 0.025
R44431 S.n4862 S.n4861 0.025
R44432 S.n3749 S.n3748 0.025
R44433 S.t158 S.n4 0.025
R44434 S.t158 S.n1373 0.025
R44435 S.t158 S.n51 0.025
R44436 S.t158 S.n82 0.025
R44437 S.t158 S.n114 0.025
R44438 S.t158 S.n1001 0.025
R44439 S.t158 S.n1033 0.025
R44440 S.t158 S.n1065 0.025
R44441 S.t158 S.n1097 0.025
R44442 S.t158 S.n1129 0.025
R44443 S.t158 S.n1167 0.025
R44444 S.n20346 S.n20345 0.024
R44445 S.n21979 S.n21978 0.024
R44446 S.n22801 S.n22800 0.024
R44447 S.n1902 S.n1901 0.024
R44448 S.n2012 S.n2011 0.024
R44449 S.n130 S.n129 0.024
R44450 S.n23007 S.n22999 0.023
R44451 S.n19522 S.n19521 0.023
R44452 S.n21151 S.n21149 0.023
R44453 S.n20817 S.n20816 0.023
R44454 S.n20348 S.n20347 0.023
R44455 S.n18665 S.n18664 0.023
R44456 S.n17797 S.n17796 0.023
R44457 S.n16903 S.n16902 0.023
R44458 S.n16000 S.n15999 0.023
R44459 S.n15071 S.n15070 0.023
R44460 S.n14133 S.n14132 0.023
R44461 S.n13169 S.n13168 0.023
R44462 S.n12196 S.n12195 0.023
R44463 S.n11197 S.n11196 0.023
R44464 S.n10189 S.n10188 0.023
R44465 S.n9155 S.n9154 0.023
R44466 S.n8112 S.n8111 0.023
R44467 S.n7043 S.n7042 0.023
R44468 S.n5965 S.n5964 0.023
R44469 S.n4860 S.n4859 0.023
R44470 S.n3747 S.n3746 0.023
R44471 S.n2617 S.n2615 0.023
R44472 S.n1917 S.n1915 0.023
R44473 S.n1914 S.n1913 0.023
R44474 S.n888 S.n885 0.023
R44475 S.n1931 S.n1929 0.023
R44476 S.n396 S.n395 0.023
R44477 S.n836 S.n833 0.023
R44478 S.n2044 S.n2043 0.023
R44479 S.n1359 S.n1357 0.023
R44480 S.t158 S.n1360 0.023
R44481 S.n20437 S.n20436 0.023
R44482 S.n20409 S.n20408 0.023
R44483 S.n20305 S.n20304 0.023
R44484 S.n19433 S.n19432 0.023
R44485 S.n18546 S.n18545 0.023
R44486 S.n17646 S.n17645 0.023
R44487 S.n16723 S.n16722 0.023
R44488 S.n15788 S.n15787 0.023
R44489 S.n14830 S.n14829 0.023
R44490 S.n13860 S.n13859 0.023
R44491 S.n12867 S.n12866 0.023
R44492 S.n11862 S.n11861 0.023
R44493 S.n10834 S.n10833 0.023
R44494 S.n9794 S.n9793 0.023
R44495 S.n8731 S.n8730 0.023
R44496 S.n7656 S.n7655 0.023
R44497 S.n6558 S.n6557 0.023
R44498 S.n5448 S.n5447 0.023
R44499 S.n4313 S.n4312 0.023
R44500 S.n3176 S.n3175 0.023
R44501 S.n1359 S.n1358 0.023
R44502 S.n1360 S.n1359 0.023
R44503 S.n763 S.n758 0.023
R44504 S.n2011 S.n2010 0.023
R44505 S.n861 S.n860 0.023
R44506 S.n2012 S.n2008 0.023
R44507 S.n2045 S.n2041 0.023
R44508 S.n19367 S.n19366 0.023
R44509 S.n393 S.n392 0.023
R44510 S.n397 S.n393 0.023
R44511 S.n364 S.n363 0.023
R44512 S.n17580 S.n17579 0.023
R44513 S.n361 S.n360 0.023
R44514 S.n365 S.n361 0.023
R44515 S.n332 S.n331 0.023
R44516 S.n329 S.n328 0.023
R44517 S.n333 S.n329 0.023
R44518 S.n300 S.n299 0.023
R44519 S.n297 S.n296 0.023
R44520 S.n301 S.n297 0.023
R44521 S.n268 S.n266 0.023
R44522 S.n269 S.n264 0.023
R44523 S.n239 S.n237 0.023
R44524 S.n9728 S.n9727 0.023
R44525 S.n240 S.n235 0.023
R44526 S.n204 S.n203 0.023
R44527 S.n7590 S.n7589 0.023
R44528 S.n201 S.n200 0.023
R44529 S.n205 S.n201 0.023
R44530 S.n172 S.n171 0.023
R44531 S.n5381 S.n5380 0.023
R44532 S.n169 S.n168 0.023
R44533 S.n173 S.n169 0.023
R44534 S.n140 S.n138 0.023
R44535 S.n3111 S.n3110 0.023
R44536 S.n1137 S.n1134 0.023
R44537 S.n141 S.n136 0.023
R44538 S.n22992 S.n22984 0.023
R44539 S.n21977 S.n21976 0.023
R44540 S.n2078 S.n2077 0.023
R44541 S.n17714 S.n17713 0.022
R44542 S.n18614 S.n18613 0.022
R44543 S.n15917 S.n15916 0.022
R44544 S.n16852 S.n16851 0.022
R44545 S.n14050 S.n14049 0.022
R44546 S.n15020 S.n15019 0.022
R44547 S.n12113 S.n12112 0.022
R44548 S.n13118 S.n13117 0.022
R44549 S.n10106 S.n10105 0.022
R44550 S.n11146 S.n11145 0.022
R44551 S.n8029 S.n8028 0.022
R44552 S.n9104 S.n9103 0.022
R44553 S.n5882 S.n5881 0.022
R44554 S.n6992 S.n6991 0.022
R44555 S.n3664 S.n3663 0.022
R44556 S.n4808 S.n4807 0.022
R44557 S.n2564 S.n2563 0.022
R44558 S.n19469 S.n19467 0.022
R44559 S.n18579 S.n18577 0.022
R44560 S.n17679 S.n17677 0.022
R44561 S.n16756 S.n16754 0.022
R44562 S.n15821 S.n15819 0.022
R44563 S.n14863 S.n14861 0.022
R44564 S.n13893 S.n13891 0.022
R44565 S.n12900 S.n12898 0.022
R44566 S.n11895 S.n11893 0.022
R44567 S.n10867 S.n10865 0.022
R44568 S.n9827 S.n9825 0.022
R44569 S.n8764 S.n8762 0.022
R44570 S.n7689 S.n7687 0.022
R44571 S.n6591 S.n6589 0.022
R44572 S.n5481 S.n5479 0.022
R44573 S.n4346 S.n4344 0.022
R44574 S.n3210 S.n3208 0.022
R44575 S.n2072 S.n2070 0.022
R44576 S.n22739 S.n22738 0.022
R44577 S.n2077 S.n2076 0.022
R44578 S.n20323 S.n20320 0.022
R44579 S.n19451 S.n19448 0.022
R44580 S.n18563 S.n18559 0.022
R44581 S.n17663 S.n17659 0.022
R44582 S.n16740 S.n16736 0.022
R44583 S.n15805 S.n15801 0.022
R44584 S.n14847 S.n14843 0.022
R44585 S.n13877 S.n13873 0.022
R44586 S.n12884 S.n12880 0.022
R44587 S.n11879 S.n11875 0.022
R44588 S.n10851 S.n10847 0.022
R44589 S.n9811 S.n9807 0.022
R44590 S.n8748 S.n8744 0.022
R44591 S.n7673 S.n7669 0.022
R44592 S.n6575 S.n6571 0.022
R44593 S.n5465 S.n5461 0.022
R44594 S.n4330 S.n4326 0.022
R44595 S.n3193 S.n3189 0.022
R44596 S.n2025 S.n2021 0.022
R44597 S.n1348 S.n1344 0.022
R44598 S.n20281 S.n20280 0.022
R44599 S.n20352 S.n20351 0.022
R44600 S.n21228 S.n21227 0.022
R44601 S.n18608 S.n18607 0.022
R44602 S.n17708 S.n17707 0.022
R44603 S.n388 S.n387 0.022
R44604 S.n16846 S.n16845 0.022
R44605 S.n15911 S.n15910 0.022
R44606 S.n356 S.n355 0.022
R44607 S.n15014 S.n15013 0.022
R44608 S.n14044 S.n14043 0.022
R44609 S.n324 S.n323 0.022
R44610 S.n13112 S.n13111 0.022
R44611 S.n12107 S.n12106 0.022
R44612 S.n292 S.n291 0.022
R44613 S.n11140 S.n11139 0.022
R44614 S.n10100 S.n10099 0.022
R44615 S.n260 S.n259 0.022
R44616 S.n9098 S.n9097 0.022
R44617 S.n8023 S.n8022 0.022
R44618 S.n231 S.n230 0.022
R44619 S.n6986 S.n6985 0.022
R44620 S.n5876 S.n5875 0.022
R44621 S.n196 S.n195 0.022
R44622 S.n4802 S.n4801 0.022
R44623 S.n3658 S.n3657 0.022
R44624 S.n164 S.n163 0.022
R44625 S.n2558 S.n2557 0.022
R44626 S.n132 S.n131 0.022
R44627 S.n20236 S.n20235 0.022
R44628 S.n19349 S.n19347 0.022
R44629 S.n18481 S.n18480 0.022
R44630 S.n17562 S.n17560 0.022
R44631 S.n16658 S.n16657 0.022
R44632 S.n15704 S.n15702 0.022
R44633 S.n14765 S.n14764 0.022
R44634 S.n13776 S.n13774 0.022
R44635 S.n12802 S.n12801 0.022
R44636 S.n11778 S.n11776 0.022
R44637 S.n10769 S.n10768 0.022
R44638 S.n9710 S.n9708 0.022
R44639 S.n8666 S.n8665 0.022
R44640 S.n7572 S.n7570 0.022
R44641 S.n6493 S.n6492 0.022
R44642 S.n5363 S.n5361 0.022
R44643 S.n4248 S.n4247 0.022
R44644 S.n1952 S.n1951 0.022
R44645 S.n3093 S.n3091 0.022
R44646 S.n925 S.n924 0.022
R44647 S.n21232 S.n21231 0.022
R44648 S.n20356 S.n20355 0.022
R44649 S.n20285 S.n20284 0.022
R44650 S.n22734 S.n22731 0.021
R44651 S.n22307 S.n22306 0.021
R44652 S.n1980 S.n1979 0.021
R44653 S.n3140 S.n3139 0.021
R44654 S.n4278 S.n4277 0.021
R44655 S.n4276 S.n4275 0.021
R44656 S.n5412 S.n5411 0.021
R44657 S.n5410 S.n5409 0.021
R44658 S.n6523 S.n6522 0.021
R44659 S.n6521 S.n6520 0.021
R44660 S.n7621 S.n7620 0.021
R44661 S.n7619 S.n7618 0.021
R44662 S.n8696 S.n8695 0.021
R44663 S.n8694 S.n8693 0.021
R44664 S.n9759 S.n9758 0.021
R44665 S.n9757 S.n9756 0.021
R44666 S.n10799 S.n10798 0.021
R44667 S.n10797 S.n10796 0.021
R44668 S.n11827 S.n11826 0.021
R44669 S.n11825 S.n11824 0.021
R44670 S.n12832 S.n12831 0.021
R44671 S.n12830 S.n12829 0.021
R44672 S.n13825 S.n13824 0.021
R44673 S.n13823 S.n13822 0.021
R44674 S.n14795 S.n14794 0.021
R44675 S.n14793 S.n14792 0.021
R44676 S.n15753 S.n15752 0.021
R44677 S.n15751 S.n15750 0.021
R44678 S.n16688 S.n16687 0.021
R44679 S.n16686 S.n16685 0.021
R44680 S.n17611 S.n17610 0.021
R44681 S.n17609 S.n17608 0.021
R44682 S.n18511 S.n18510 0.021
R44683 S.n18509 S.n18508 0.021
R44684 S.n19398 S.n19397 0.021
R44685 S.n19396 S.n19395 0.021
R44686 S.n20266 S.n20265 0.021
R44687 S.n20264 S.n20263 0.021
R44688 S.n20393 S.n20392 0.021
R44689 S.n21212 S.n21211 0.021
R44690 S.n22733 S.n22732 0.021
R44691 S.n2055 S.n2054 0.021
R44692 S.n3224 S.n3223 0.021
R44693 S.n4362 S.n4361 0.021
R44694 S.n4360 S.n4359 0.021
R44695 S.n5497 S.n5496 0.021
R44696 S.n5495 S.n5494 0.021
R44697 S.n6607 S.n6606 0.021
R44698 S.n6605 S.n6604 0.021
R44699 S.n7705 S.n7704 0.021
R44700 S.n7703 S.n7702 0.021
R44701 S.n8780 S.n8779 0.021
R44702 S.n8778 S.n8777 0.021
R44703 S.n9843 S.n9842 0.021
R44704 S.n9841 S.n9840 0.021
R44705 S.n10883 S.n10882 0.021
R44706 S.n10881 S.n10880 0.021
R44707 S.n11911 S.n11910 0.021
R44708 S.n11909 S.n11908 0.021
R44709 S.n12916 S.n12915 0.021
R44710 S.n12914 S.n12913 0.021
R44711 S.n13909 S.n13908 0.021
R44712 S.n13907 S.n13906 0.021
R44713 S.n14879 S.n14878 0.021
R44714 S.n14877 S.n14876 0.021
R44715 S.n15837 S.n15836 0.021
R44716 S.n15835 S.n15834 0.021
R44717 S.n16772 S.n16771 0.021
R44718 S.n16770 S.n16769 0.021
R44719 S.n17695 S.n17694 0.021
R44720 S.n17693 S.n17692 0.021
R44721 S.n18595 S.n18594 0.021
R44722 S.n19485 S.n19484 0.021
R44723 S.n20230 S.n20229 0.021
R44724 S.n2132 S.n2131 0.021
R44725 S.n3284 S.n3283 0.021
R44726 S.n4423 S.n4422 0.021
R44727 S.n4421 S.n4420 0.021
R44728 S.n5558 S.n5557 0.021
R44729 S.n5556 S.n5555 0.021
R44730 S.n6668 S.n6667 0.021
R44731 S.n6666 S.n6665 0.021
R44732 S.n7766 S.n7765 0.021
R44733 S.n7764 S.n7763 0.021
R44734 S.n8841 S.n8840 0.021
R44735 S.n8839 S.n8838 0.021
R44736 S.n9904 S.n9903 0.021
R44737 S.n9902 S.n9901 0.021
R44738 S.n10944 S.n10943 0.021
R44739 S.n10942 S.n10941 0.021
R44740 S.n11972 S.n11971 0.021
R44741 S.n11970 S.n11969 0.021
R44742 S.n12977 S.n12976 0.021
R44743 S.n12975 S.n12974 0.021
R44744 S.n13970 S.n13969 0.021
R44745 S.n13968 S.n13967 0.021
R44746 S.n14940 S.n14939 0.021
R44747 S.n14938 S.n14937 0.021
R44748 S.n15898 S.n15897 0.021
R44749 S.n15896 S.n15895 0.021
R44750 S.n16833 S.n16832 0.021
R44751 S.n17760 S.n17759 0.021
R44752 S.n18475 S.n18474 0.021
R44753 S.n2191 S.n2190 0.021
R44754 S.n3344 S.n3343 0.021
R44755 S.n4484 S.n4483 0.021
R44756 S.n4482 S.n4481 0.021
R44757 S.n5619 S.n5618 0.021
R44758 S.n5617 S.n5616 0.021
R44759 S.n6729 S.n6728 0.021
R44760 S.n6727 S.n6726 0.021
R44761 S.n7827 S.n7826 0.021
R44762 S.n7825 S.n7824 0.021
R44763 S.n8902 S.n8901 0.021
R44764 S.n8900 S.n8899 0.021
R44765 S.n9965 S.n9964 0.021
R44766 S.n9963 S.n9962 0.021
R44767 S.n11005 S.n11004 0.021
R44768 S.n11003 S.n11002 0.021
R44769 S.n12033 S.n12032 0.021
R44770 S.n12031 S.n12030 0.021
R44771 S.n13038 S.n13037 0.021
R44772 S.n13036 S.n13035 0.021
R44773 S.n14031 S.n14030 0.021
R44774 S.n14029 S.n14028 0.021
R44775 S.n15001 S.n15000 0.021
R44776 S.n15963 S.n15962 0.021
R44777 S.n16652 S.n16651 0.021
R44778 S.n2250 S.n2249 0.021
R44779 S.n3404 S.n3403 0.021
R44780 S.n4545 S.n4544 0.021
R44781 S.n4543 S.n4542 0.021
R44782 S.n5680 S.n5679 0.021
R44783 S.n5678 S.n5677 0.021
R44784 S.n6790 S.n6789 0.021
R44785 S.n6788 S.n6787 0.021
R44786 S.n7888 S.n7887 0.021
R44787 S.n7886 S.n7885 0.021
R44788 S.n8963 S.n8962 0.021
R44789 S.n8961 S.n8960 0.021
R44790 S.n10026 S.n10025 0.021
R44791 S.n10024 S.n10023 0.021
R44792 S.n11066 S.n11065 0.021
R44793 S.n11064 S.n11063 0.021
R44794 S.n12094 S.n12093 0.021
R44795 S.n12092 S.n12091 0.021
R44796 S.n13099 S.n13098 0.021
R44797 S.n14096 S.n14095 0.021
R44798 S.n14759 S.n14758 0.021
R44799 S.n2309 S.n2308 0.021
R44800 S.n3464 S.n3463 0.021
R44801 S.n4606 S.n4605 0.021
R44802 S.n4604 S.n4603 0.021
R44803 S.n5741 S.n5740 0.021
R44804 S.n5739 S.n5738 0.021
R44805 S.n6851 S.n6850 0.021
R44806 S.n6849 S.n6848 0.021
R44807 S.n7949 S.n7948 0.021
R44808 S.n7947 S.n7946 0.021
R44809 S.n9024 S.n9023 0.021
R44810 S.n9022 S.n9021 0.021
R44811 S.n10087 S.n10086 0.021
R44812 S.n10085 S.n10084 0.021
R44813 S.n11127 S.n11126 0.021
R44814 S.n12159 S.n12158 0.021
R44815 S.n12796 S.n12795 0.021
R44816 S.n2368 S.n2367 0.021
R44817 S.n3524 S.n3523 0.021
R44818 S.n4667 S.n4666 0.021
R44819 S.n4665 S.n4664 0.021
R44820 S.n5802 S.n5801 0.021
R44821 S.n5800 S.n5799 0.021
R44822 S.n6912 S.n6911 0.021
R44823 S.n6910 S.n6909 0.021
R44824 S.n8010 S.n8009 0.021
R44825 S.n8008 S.n8007 0.021
R44826 S.n9085 S.n9084 0.021
R44827 S.n10152 S.n10151 0.021
R44828 S.n10763 S.n10762 0.021
R44829 S.n2427 S.n2426 0.021
R44830 S.n3584 S.n3583 0.021
R44831 S.n4728 S.n4727 0.021
R44832 S.n4726 S.n4725 0.021
R44833 S.n5863 S.n5862 0.021
R44834 S.n5861 S.n5860 0.021
R44835 S.n6973 S.n6972 0.021
R44836 S.n8075 S.n8074 0.021
R44837 S.n8660 S.n8659 0.021
R44838 S.n2486 S.n2485 0.021
R44839 S.n3644 S.n3643 0.021
R44840 S.n4789 S.n4788 0.021
R44841 S.n5928 S.n5927 0.021
R44842 S.n6487 S.n6486 0.021
R44843 S.n4242 S.n4241 0.021
R44844 S.n22693 S.n22691 0.021
R44845 S.n21195 S.n21194 0.021
R44846 S.n20376 S.n20375 0.021
R44847 S.n20249 S.n20248 0.021
R44848 S.n19381 S.n19380 0.021
R44849 S.n18494 S.n18493 0.021
R44850 S.n17594 S.n17593 0.021
R44851 S.n16671 S.n16670 0.021
R44852 S.n15736 S.n15735 0.021
R44853 S.n14778 S.n14777 0.021
R44854 S.n13808 S.n13807 0.021
R44855 S.n12815 S.n12814 0.021
R44856 S.n11810 S.n11809 0.021
R44857 S.n10782 S.n10781 0.021
R44858 S.n9742 S.n9741 0.021
R44859 S.n8679 S.n8678 0.021
R44860 S.n7604 S.n7603 0.021
R44861 S.n6506 S.n6505 0.021
R44862 S.n5395 S.n5394 0.021
R44863 S.n4261 S.n4260 0.021
R44864 S.n3125 S.n3124 0.021
R44865 S.n1965 S.n1964 0.021
R44866 S.n22704 S.n22703 0.021
R44867 S.n21252 S.n21251 0.021
R44868 S.n17743 S.n17742 0.021
R44869 S.n16816 S.n16815 0.021
R44870 S.n15881 S.n15880 0.021
R44871 S.n14923 S.n14922 0.021
R44872 S.n13953 S.n13952 0.021
R44873 S.n12960 S.n12959 0.021
R44874 S.n11955 S.n11954 0.021
R44875 S.n10927 S.n10926 0.021
R44876 S.n9887 S.n9886 0.021
R44877 S.n8824 S.n8823 0.021
R44878 S.n7749 S.n7748 0.021
R44879 S.n6651 S.n6650 0.021
R44880 S.n5541 S.n5540 0.021
R44881 S.n4406 S.n4405 0.021
R44882 S.n3269 S.n3268 0.021
R44883 S.n2117 S.n2116 0.021
R44884 S.n19469 S.n19468 0.021
R44885 S.n18579 S.n18578 0.021
R44886 S.n17679 S.n17678 0.021
R44887 S.n16756 S.n16755 0.021
R44888 S.n15821 S.n15820 0.021
R44889 S.n14863 S.n14862 0.021
R44890 S.n13893 S.n13892 0.021
R44891 S.n12900 S.n12899 0.021
R44892 S.n11895 S.n11894 0.021
R44893 S.n10867 S.n10866 0.021
R44894 S.n9827 S.n9826 0.021
R44895 S.n8764 S.n8763 0.021
R44896 S.n7689 S.n7688 0.021
R44897 S.n6591 S.n6590 0.021
R44898 S.n5481 S.n5480 0.021
R44899 S.n4346 S.n4345 0.021
R44900 S.n3210 S.n3209 0.021
R44901 S.n20237 S.n20236 0.021
R44902 S.n20423 S.n20422 0.021
R44903 S.n20329 S.n20328 0.021
R44904 S.n19457 S.n19456 0.021
R44905 S.n2072 S.n2071 0.021
R44906 S.n2103 S.n2102 0.021
R44907 S.n3255 S.n3254 0.021
R44908 S.n4392 S.n4391 0.021
R44909 S.n5527 S.n5526 0.021
R44910 S.n6637 S.n6636 0.021
R44911 S.n7735 S.n7734 0.021
R44912 S.n8810 S.n8809 0.021
R44913 S.n9873 S.n9872 0.021
R44914 S.n10913 S.n10912 0.021
R44915 S.n11941 S.n11940 0.021
R44916 S.n12946 S.n12945 0.021
R44917 S.n13939 S.n13938 0.021
R44918 S.n14909 S.n14908 0.021
R44919 S.n15867 S.n15866 0.021
R44920 S.n16802 S.n16801 0.021
R44921 S.n17729 S.n17728 0.021
R44922 S.n18629 S.n18628 0.021
R44923 S.n19351 S.n19349 0.021
R44924 S.n18482 S.n18481 0.021
R44925 S.n15946 S.n15945 0.021
R44926 S.n14984 S.n14983 0.021
R44927 S.n14014 S.n14013 0.021
R44928 S.n13021 S.n13020 0.021
R44929 S.n12016 S.n12015 0.021
R44930 S.n10988 S.n10987 0.021
R44931 S.n9948 S.n9947 0.021
R44932 S.n8885 S.n8884 0.021
R44933 S.n7810 S.n7809 0.021
R44934 S.n6712 S.n6711 0.021
R44935 S.n5602 S.n5601 0.021
R44936 S.n4467 S.n4466 0.021
R44937 S.n3329 S.n3328 0.021
R44938 S.n2176 S.n2175 0.021
R44939 S.n2162 S.n2161 0.021
R44940 S.n3315 S.n3314 0.021
R44941 S.n4453 S.n4452 0.021
R44942 S.n5588 S.n5587 0.021
R44943 S.n6698 S.n6697 0.021
R44944 S.n7796 S.n7795 0.021
R44945 S.n8871 S.n8870 0.021
R44946 S.n9934 S.n9933 0.021
R44947 S.n10974 S.n10973 0.021
R44948 S.n12002 S.n12001 0.021
R44949 S.n13007 S.n13006 0.021
R44950 S.n14000 S.n13999 0.021
R44951 S.n14970 S.n14969 0.021
R44952 S.n15932 S.n15931 0.021
R44953 S.n16867 S.n16866 0.021
R44954 S.n17564 S.n17562 0.021
R44955 S.n16659 S.n16658 0.021
R44956 S.n14079 S.n14078 0.021
R44957 S.n13082 S.n13081 0.021
R44958 S.n12077 S.n12076 0.021
R44959 S.n11049 S.n11048 0.021
R44960 S.n10009 S.n10008 0.021
R44961 S.n8946 S.n8945 0.021
R44962 S.n7871 S.n7870 0.021
R44963 S.n6773 S.n6772 0.021
R44964 S.n5663 S.n5662 0.021
R44965 S.n4528 S.n4527 0.021
R44966 S.n3389 S.n3388 0.021
R44967 S.n2235 S.n2234 0.021
R44968 S.n2221 S.n2220 0.021
R44969 S.n3375 S.n3374 0.021
R44970 S.n4514 S.n4513 0.021
R44971 S.n5649 S.n5648 0.021
R44972 S.n6759 S.n6758 0.021
R44973 S.n7857 S.n7856 0.021
R44974 S.n8932 S.n8931 0.021
R44975 S.n9995 S.n9994 0.021
R44976 S.n11035 S.n11034 0.021
R44977 S.n12063 S.n12062 0.021
R44978 S.n13068 S.n13067 0.021
R44979 S.n14065 S.n14064 0.021
R44980 S.n15035 S.n15034 0.021
R44981 S.n15706 S.n15704 0.021
R44982 S.n14766 S.n14765 0.021
R44983 S.n12142 S.n12141 0.021
R44984 S.n11110 S.n11109 0.021
R44985 S.n10070 S.n10069 0.021
R44986 S.n9007 S.n9006 0.021
R44987 S.n7932 S.n7931 0.021
R44988 S.n6834 S.n6833 0.021
R44989 S.n5724 S.n5723 0.021
R44990 S.n4589 S.n4588 0.021
R44991 S.n3449 S.n3448 0.021
R44992 S.n2294 S.n2293 0.021
R44993 S.n2280 S.n2279 0.021
R44994 S.n3435 S.n3434 0.021
R44995 S.n4575 S.n4574 0.021
R44996 S.n5710 S.n5709 0.021
R44997 S.n6820 S.n6819 0.021
R44998 S.n7918 S.n7917 0.021
R44999 S.n8993 S.n8992 0.021
R45000 S.n10056 S.n10055 0.021
R45001 S.n11096 S.n11095 0.021
R45002 S.n12128 S.n12127 0.021
R45003 S.n13133 S.n13132 0.021
R45004 S.n13778 S.n13776 0.021
R45005 S.n12803 S.n12802 0.021
R45006 S.n10135 S.n10134 0.021
R45007 S.n9068 S.n9067 0.021
R45008 S.n7993 S.n7992 0.021
R45009 S.n6895 S.n6894 0.021
R45010 S.n5785 S.n5784 0.021
R45011 S.n4650 S.n4649 0.021
R45012 S.n3509 S.n3508 0.021
R45013 S.n2353 S.n2352 0.021
R45014 S.n2339 S.n2338 0.021
R45015 S.n3495 S.n3494 0.021
R45016 S.n4636 S.n4635 0.021
R45017 S.n5771 S.n5770 0.021
R45018 S.n6881 S.n6880 0.021
R45019 S.n7979 S.n7978 0.021
R45020 S.n9054 S.n9053 0.021
R45021 S.n10121 S.n10120 0.021
R45022 S.n11161 S.n11160 0.021
R45023 S.n11780 S.n11778 0.021
R45024 S.n10770 S.n10769 0.021
R45025 S.n8058 S.n8057 0.021
R45026 S.n6956 S.n6955 0.021
R45027 S.n5846 S.n5845 0.021
R45028 S.n4711 S.n4710 0.021
R45029 S.n3569 S.n3568 0.021
R45030 S.n2412 S.n2411 0.021
R45031 S.n2398 S.n2397 0.021
R45032 S.n3555 S.n3554 0.021
R45033 S.n4697 S.n4696 0.021
R45034 S.n5832 S.n5831 0.021
R45035 S.n6942 S.n6941 0.021
R45036 S.n8044 S.n8043 0.021
R45037 S.n9119 S.n9118 0.021
R45038 S.n9712 S.n9710 0.021
R45039 S.n8667 S.n8666 0.021
R45040 S.n5911 S.n5910 0.021
R45041 S.n4772 S.n4771 0.021
R45042 S.n3629 S.n3628 0.021
R45043 S.n2471 S.n2470 0.021
R45044 S.n2457 S.n2456 0.021
R45045 S.n3615 S.n3614 0.021
R45046 S.n4758 S.n4757 0.021
R45047 S.n5897 S.n5896 0.021
R45048 S.n7007 S.n7006 0.021
R45049 S.n7574 S.n7572 0.021
R45050 S.n6494 S.n6493 0.021
R45051 S.n3693 S.n3692 0.021
R45052 S.n2530 S.n2529 0.021
R45053 S.n2516 S.n2515 0.021
R45054 S.n3679 S.n3678 0.021
R45055 S.n4823 S.n4822 0.021
R45056 S.n5365 S.n5363 0.021
R45057 S.n4249 S.n4248 0.021
R45058 S.n1953 S.n1952 0.021
R45059 S.n2579 S.n2578 0.021
R45060 S.n3095 S.n3093 0.021
R45061 S.n926 S.n925 0.021
R45062 S.n911 S.n905 0.021
R45063 S.n389 S.n382 0.021
R45064 S.n357 S.n350 0.021
R45065 S.n325 S.n318 0.021
R45066 S.n293 S.n286 0.021
R45067 S.n261 S.n254 0.021
R45068 S.n232 S.n225 0.021
R45069 S.n197 S.n190 0.021
R45070 S.n165 S.n158 0.021
R45071 S.n133 S.n126 0.021
R45072 S.n887 S.n886 0.02
R45073 S.n22991 S.n22990 0.02
R45074 S.n23006 S.n23000 0.02
R45075 S.n1355 S.n1354 0.02
R45076 S.n846 S.n845 0.02
R45077 S.n7 S.n6 0.02
R45078 S.n54 S.n53 0.02
R45079 S.n87 S.n86 0.02
R45080 S.n118 S.n117 0.02
R45081 S.n1005 S.n1004 0.02
R45082 S.n1038 S.n1037 0.02
R45083 S.n1069 S.n1068 0.02
R45084 S.n1101 S.n1100 0.02
R45085 S.n937 S.n936 0.02
R45086 S.n22755 S.n22754 0.02
R45087 S.n20397 S.n20396 0.02
R45088 S.n21216 S.n21215 0.02
R45089 S.n22740 S.n22737 0.02
R45090 S.n18599 S.n18598 0.02
R45091 S.n19489 S.n19488 0.02
R45092 S.n20237 S.n20233 0.02
R45093 S.n20282 S.n20279 0.02
R45094 S.n20353 S.n20350 0.02
R45095 S.n21229 S.n21226 0.02
R45096 S.n19351 S.n19350 0.02
R45097 S.n18611 S.n18610 0.02
R45098 S.n17711 S.n17710 0.02
R45099 S.n16837 S.n16836 0.02
R45100 S.n17764 S.n17763 0.02
R45101 S.n18482 S.n18478 0.02
R45102 S.n17564 S.n17563 0.02
R45103 S.n16849 S.n16848 0.02
R45104 S.n15914 S.n15913 0.02
R45105 S.n15005 S.n15004 0.02
R45106 S.n15967 S.n15966 0.02
R45107 S.n16659 S.n16655 0.02
R45108 S.n15706 S.n15705 0.02
R45109 S.n15017 S.n15016 0.02
R45110 S.n14047 S.n14046 0.02
R45111 S.n13103 S.n13102 0.02
R45112 S.n14100 S.n14099 0.02
R45113 S.n14766 S.n14762 0.02
R45114 S.n13778 S.n13777 0.02
R45115 S.n13115 S.n13114 0.02
R45116 S.n12110 S.n12109 0.02
R45117 S.n11131 S.n11130 0.02
R45118 S.n12163 S.n12162 0.02
R45119 S.n12803 S.n12799 0.02
R45120 S.n11780 S.n11779 0.02
R45121 S.n11143 S.n11142 0.02
R45122 S.n10103 S.n10102 0.02
R45123 S.n9089 S.n9088 0.02
R45124 S.n10156 S.n10155 0.02
R45125 S.n10770 S.n10766 0.02
R45126 S.n9712 S.n9711 0.02
R45127 S.n9101 S.n9100 0.02
R45128 S.n8026 S.n8025 0.02
R45129 S.n6977 S.n6976 0.02
R45130 S.n8079 S.n8078 0.02
R45131 S.n8667 S.n8663 0.02
R45132 S.n7574 S.n7573 0.02
R45133 S.n6989 S.n6988 0.02
R45134 S.n5879 S.n5878 0.02
R45135 S.n4793 S.n4792 0.02
R45136 S.n5932 S.n5931 0.02
R45137 S.n6494 S.n6490 0.02
R45138 S.n5365 S.n5364 0.02
R45139 S.n4805 S.n4804 0.02
R45140 S.n3661 S.n3660 0.02
R45141 S.n2549 S.n2548 0.02
R45142 S.n3713 S.n3712 0.02
R45143 S.n4249 S.n4245 0.02
R45144 S.n1953 S.n1949 0.02
R45145 S.n3095 S.n3094 0.02
R45146 S.n2561 S.n2560 0.02
R45147 S.n926 S.n922 0.02
R45148 S.n1364 S.n1363 0.02
R45149 S.n20440 S.n20439 0.019
R45150 S.n21153 S.n21152 0.019
R45151 S.t158 S.n1313 0.019
R45152 S.n1322 S.n1321 0.019
R45153 S.n1836 S.n1835 0.019
R45154 S.n18567 S.n18566 0.019
R45155 S.n17667 S.n17666 0.019
R45156 S.n16744 S.n16743 0.019
R45157 S.n15809 S.n15808 0.019
R45158 S.n14851 S.n14850 0.019
R45159 S.n13881 S.n13880 0.019
R45160 S.n12888 S.n12887 0.019
R45161 S.n11883 S.n11882 0.019
R45162 S.n10855 S.n10854 0.019
R45163 S.n9815 S.n9814 0.019
R45164 S.n8752 S.n8751 0.019
R45165 S.n7677 S.n7676 0.019
R45166 S.n6579 S.n6578 0.019
R45167 S.n5469 S.n5468 0.019
R45168 S.n4334 S.n4333 0.019
R45169 S.n3197 S.n3196 0.019
R45170 S.n2029 S.n2028 0.019
R45171 S.n20391 S.n20390 0.019
R45172 S.n21210 S.n21209 0.019
R45173 S.n18593 S.n18592 0.019
R45174 S.n19483 S.n19482 0.019
R45175 S.n16831 S.n16830 0.019
R45176 S.n17758 S.n17757 0.019
R45177 S.n14999 S.n14998 0.019
R45178 S.n15961 S.n15960 0.019
R45179 S.n13097 S.n13096 0.019
R45180 S.n14094 S.n14093 0.019
R45181 S.n11125 S.n11124 0.019
R45182 S.n12157 S.n12156 0.019
R45183 S.n9083 S.n9082 0.019
R45184 S.n10150 S.n10149 0.019
R45185 S.n6971 S.n6970 0.019
R45186 S.n8073 S.n8072 0.019
R45187 S.n4787 S.n4786 0.019
R45188 S.n5926 S.n5925 0.019
R45189 S.n2545 S.n2544 0.019
R45190 S.n3708 S.n3707 0.019
R45191 S.n968 S.n965 0.018
R45192 S.n426 S.n422 0.018
R45193 S.n1908 S.n1906 0.018
R45194 S.n1454 S.n1452 0.018
R45195 S.n2609 S.n2606 0.018
R45196 S.n2648 S.n2646 0.018
R45197 S.n3740 S.n3737 0.018
R45198 S.n3793 S.n3791 0.018
R45199 S.n4853 S.n4850 0.018
R45200 S.n4923 S.n4921 0.018
R45201 S.n5958 S.n5955 0.018
R45202 S.n6041 S.n6039 0.018
R45203 S.n7036 S.n7033 0.018
R45204 S.n7136 S.n7134 0.018
R45205 S.n8105 S.n8102 0.018
R45206 S.n8218 S.n8216 0.018
R45207 S.n9148 S.n9145 0.018
R45208 S.n9278 S.n9276 0.018
R45209 S.n10182 S.n10179 0.018
R45210 S.n10325 S.n10323 0.018
R45211 S.n11190 S.n11187 0.018
R45212 S.n11350 S.n11348 0.018
R45213 S.n12189 S.n12186 0.018
R45214 S.n12362 S.n12360 0.018
R45215 S.n13162 S.n13159 0.018
R45216 S.n13352 S.n13350 0.018
R45217 S.n14126 S.n14123 0.018
R45218 S.n14329 S.n14327 0.018
R45219 S.n15064 S.n15061 0.018
R45220 S.n15284 S.n15282 0.018
R45221 S.n15993 S.n15990 0.018
R45222 S.n16226 S.n16224 0.018
R45223 S.n16896 S.n16893 0.018
R45224 S.n17146 S.n17144 0.018
R45225 S.n17790 S.n17787 0.018
R45226 S.n18053 S.n18051 0.018
R45227 S.n18658 S.n18655 0.018
R45228 S.n18938 S.n18936 0.018
R45229 S.n19515 S.n19512 0.018
R45230 S.n19808 S.n19806 0.018
R45231 S.n21165 S.n21162 0.018
R45232 S.n20446 S.n20444 0.018
R45233 S.n21183 S.n21180 0.018
R45234 S.n21290 S.n21288 0.018
R45235 S.n22781 S.n22778 0.018
R45236 S.n22281 S.n22276 0.018
R45237 S.n22796 S.n22794 0.018
R45238 S.n21629 S.n21628 0.018
R45239 S.n20806 S.n20805 0.018
R45240 S.n1313 S.n1312 0.018
R45241 S.n20408 S.n20407 0.018
R45242 S.n20413 S.n20412 0.018
R45243 S.n20304 S.n20303 0.018
R45244 S.n20309 S.n20308 0.018
R45245 S.n19432 S.n19431 0.018
R45246 S.n19437 S.n19436 0.018
R45247 S.n18545 S.n18544 0.018
R45248 S.n18550 S.n18549 0.018
R45249 S.n17645 S.n17644 0.018
R45250 S.n17650 S.n17649 0.018
R45251 S.n16722 S.n16721 0.018
R45252 S.n16727 S.n16726 0.018
R45253 S.n15787 S.n15786 0.018
R45254 S.n15792 S.n15791 0.018
R45255 S.n14829 S.n14828 0.018
R45256 S.n14834 S.n14833 0.018
R45257 S.n13859 S.n13858 0.018
R45258 S.n13864 S.n13863 0.018
R45259 S.n12866 S.n12865 0.018
R45260 S.n12871 S.n12870 0.018
R45261 S.n11861 S.n11860 0.018
R45262 S.n11866 S.n11865 0.018
R45263 S.n10833 S.n10832 0.018
R45264 S.n10838 S.n10837 0.018
R45265 S.n9793 S.n9792 0.018
R45266 S.n9798 S.n9797 0.018
R45267 S.n8730 S.n8729 0.018
R45268 S.n8735 S.n8734 0.018
R45269 S.n7655 S.n7654 0.018
R45270 S.n7660 S.n7659 0.018
R45271 S.n6557 S.n6556 0.018
R45272 S.n6562 S.n6561 0.018
R45273 S.n5447 S.n5446 0.018
R45274 S.n5452 S.n5451 0.018
R45275 S.n4312 S.n4311 0.018
R45276 S.n4317 S.n4316 0.018
R45277 S.n3175 S.n3174 0.018
R45278 S.n3180 S.n3179 0.018
R45279 S.n2043 S.n2042 0.018
R45280 S.n2040 S.n2039 0.018
R45281 S S.n1441 0.018
R45282 S.n1317 S.n1316 0.018
R45283 S.n386 S.n385 0.018
R45284 S.n354 S.n353 0.018
R45285 S.n322 S.n321 0.018
R45286 S.n290 S.n289 0.018
R45287 S.n258 S.n257 0.018
R45288 S.n229 S.n228 0.018
R45289 S.n194 S.n193 0.018
R45290 S.n162 S.n161 0.018
R45291 S.n21626 S.n21625 0.017
R45292 S.n20803 S.n20802 0.017
R45293 S.n913 S.n912 0.017
R45294 S.n391 S.n390 0.017
R45295 S.n359 S.n358 0.017
R45296 S.n327 S.n326 0.017
R45297 S.n295 S.n294 0.017
R45298 S.n263 S.n262 0.017
R45299 S.n234 S.n233 0.017
R45300 S.n199 S.n198 0.017
R45301 S.n167 S.n166 0.017
R45302 S.n135 S.n134 0.017
R45303 S.n22300 S.n22299 0.017
R45304 S.n22322 S.n22321 0.017
R45305 S.n20818 S.n20814 0.017
R45306 S.n382 S.n381 0.017
R45307 S.n350 S.n349 0.017
R45308 S.n318 S.n317 0.017
R45309 S.n286 S.n285 0.017
R45310 S.n254 S.n253 0.017
R45311 S.n225 S.n224 0.017
R45312 S.n190 S.n189 0.017
R45313 S.n158 S.n157 0.017
R45314 S.n1139 S.n1138 0.017
R45315 S.n2978 S.n2973 0.016
R45316 S.n4105 S.n4100 0.016
R45317 S.n5217 S.n5212 0.016
R45318 S.n6317 S.n6312 0.016
R45319 S.n7394 S.n7389 0.016
R45320 S.n8458 S.n8453 0.016
R45321 S.n9500 S.n9495 0.016
R45322 S.n10529 S.n10524 0.016
R45323 S.n11536 S.n11531 0.016
R45324 S.n12530 S.n12525 0.016
R45325 S.n13502 S.n13497 0.016
R45326 S.n14461 S.n14456 0.016
R45327 S.n15398 S.n15393 0.016
R45328 S.n16322 S.n16317 0.016
R45329 S.n17224 S.n17219 0.016
R45330 S.n18113 S.n18108 0.016
R45331 S.n18978 S.n18973 0.016
R45332 S.n19830 S.n19825 0.016
R45333 S.n2079 S.n2078 0.016
R45334 S.n1799 S.n1795 0.016
R45335 S.n19370 S.n19362 0.016
R45336 S.n17583 S.n17575 0.016
R45337 S.n15725 S.n15717 0.016
R45338 S.n13797 S.n13789 0.016
R45339 S.n11799 S.n11791 0.016
R45340 S.n9731 S.n9723 0.016
R45341 S.n7593 S.n7585 0.016
R45342 S.n5384 S.n5376 0.016
R45343 S.n3114 S.n3106 0.016
R45344 S.n19467 S.n19466 0.016
R45345 S.n18577 S.n18576 0.016
R45346 S.n17677 S.n17676 0.016
R45347 S.n16754 S.n16753 0.016
R45348 S.n15819 S.n15818 0.016
R45349 S.n14861 S.n14860 0.016
R45350 S.n13891 S.n13890 0.016
R45351 S.n12898 S.n12897 0.016
R45352 S.n11893 S.n11892 0.016
R45353 S.n10865 S.n10864 0.016
R45354 S.n9825 S.n9824 0.016
R45355 S.n8762 S.n8761 0.016
R45356 S.n7687 S.n7686 0.016
R45357 S.n6589 S.n6588 0.016
R45358 S.n5479 S.n5478 0.016
R45359 S.n4344 S.n4343 0.016
R45360 S.n3208 S.n3207 0.016
R45361 S.n2070 S.n2069 0.016
R45362 S.n21984 S.n21983 0.015
R45363 S.n21950 S.n21949 0.015
R45364 S.n21628 S.n21627 0.015
R45365 S.n20805 S.n20804 0.015
R45366 S.n21172 S.n21170 0.015
R45367 S.t41 S.n22834 0.015
R45368 S.t41 S.n22825 0.015
R45369 S.n22731 S.n22730 0.015
R45370 S.t41 S.n22810 0.015
R45371 S.n17713 S.n17712 0.015
R45372 S.n18613 S.n18612 0.015
R45373 S.n20324 S.n20318 0.015
R45374 S.n20324 S.n20323 0.015
R45375 S.n20323 S.n20322 0.015
R45376 S.n19452 S.n19446 0.015
R45377 S.n19452 S.n19451 0.015
R45378 S.n19451 S.n19450 0.015
R45379 S.n18565 S.n18564 0.015
R45380 S.n18564 S.n18563 0.015
R45381 S.n18563 S.n18562 0.015
R45382 S.n17665 S.n17664 0.015
R45383 S.n17664 S.n17663 0.015
R45384 S.n17663 S.n17662 0.015
R45385 S.n16742 S.n16741 0.015
R45386 S.n16741 S.n16740 0.015
R45387 S.n16740 S.n16739 0.015
R45388 S.n15807 S.n15806 0.015
R45389 S.n15806 S.n15805 0.015
R45390 S.n15805 S.n15804 0.015
R45391 S.n14849 S.n14848 0.015
R45392 S.n14848 S.n14847 0.015
R45393 S.n14847 S.n14846 0.015
R45394 S.n13879 S.n13878 0.015
R45395 S.n13878 S.n13877 0.015
R45396 S.n13877 S.n13876 0.015
R45397 S.n12886 S.n12885 0.015
R45398 S.n12885 S.n12884 0.015
R45399 S.n12884 S.n12883 0.015
R45400 S.n11881 S.n11880 0.015
R45401 S.n11880 S.n11879 0.015
R45402 S.n11879 S.n11878 0.015
R45403 S.n10853 S.n10852 0.015
R45404 S.n10852 S.n10851 0.015
R45405 S.n10851 S.n10850 0.015
R45406 S.n9813 S.n9812 0.015
R45407 S.n9812 S.n9811 0.015
R45408 S.n9811 S.n9810 0.015
R45409 S.n8750 S.n8749 0.015
R45410 S.n8749 S.n8748 0.015
R45411 S.n8748 S.n8747 0.015
R45412 S.n7675 S.n7674 0.015
R45413 S.n7674 S.n7673 0.015
R45414 S.n7673 S.n7672 0.015
R45415 S.n6577 S.n6576 0.015
R45416 S.n6576 S.n6575 0.015
R45417 S.n6575 S.n6574 0.015
R45418 S.n5467 S.n5466 0.015
R45419 S.n5466 S.n5465 0.015
R45420 S.n5465 S.n5464 0.015
R45421 S.n4332 S.n4331 0.015
R45422 S.n4331 S.n4330 0.015
R45423 S.n4330 S.n4329 0.015
R45424 S.n3195 S.n3194 0.015
R45425 S.n3194 S.n3193 0.015
R45426 S.n3193 S.n3192 0.015
R45427 S.n2027 S.n2026 0.015
R45428 S.n2026 S.n2025 0.015
R45429 S.n2025 S.n2024 0.015
R45430 S.n1349 S.n1348 0.015
R45431 S.n1348 S.n1347 0.015
R45432 S.n21231 S.n21230 0.015
R45433 S.n20355 S.n20354 0.015
R45434 S.n20284 S.n20283 0.015
R45435 S.n863 S.n862 0.015
R45436 S.n15916 S.n15915 0.015
R45437 S.n16851 S.n16850 0.015
R45438 S.n14049 S.n14048 0.015
R45439 S.n15019 S.n15018 0.015
R45440 S.n12112 S.n12111 0.015
R45441 S.n13117 S.n13116 0.015
R45442 S.n10105 S.n10104 0.015
R45443 S.n11145 S.n11144 0.015
R45444 S.n8028 S.n8027 0.015
R45445 S.n9103 S.n9102 0.015
R45446 S.n5881 S.n5880 0.015
R45447 S.n6991 S.n6990 0.015
R45448 S.n3663 S.n3662 0.015
R45449 S.n4807 S.n4806 0.015
R45450 S.n2563 S.n2562 0.015
R45451 S.n2079 S.n2074 0.015
R45452 S.n21198 S.n21197 0.015
R45453 S.n20379 S.n20378 0.015
R45454 S.n20252 S.n20251 0.015
R45455 S.n19384 S.n19383 0.015
R45456 S.n18497 S.n18496 0.015
R45457 S.n17597 S.n17596 0.015
R45458 S.n16674 S.n16673 0.015
R45459 S.n15739 S.n15738 0.015
R45460 S.n14781 S.n14780 0.015
R45461 S.n13811 S.n13810 0.015
R45462 S.n12818 S.n12817 0.015
R45463 S.n11813 S.n11812 0.015
R45464 S.n10785 S.n10784 0.015
R45465 S.n9745 S.n9744 0.015
R45466 S.n8682 S.n8681 0.015
R45467 S.n7607 S.n7606 0.015
R45468 S.n6509 S.n6508 0.015
R45469 S.n5398 S.n5397 0.015
R45470 S.n4264 S.n4263 0.015
R45471 S.n3128 S.n3127 0.015
R45472 S.n1968 S.n1967 0.015
R45473 S.n17746 S.n17745 0.015
R45474 S.n16819 S.n16818 0.015
R45475 S.n15884 S.n15883 0.015
R45476 S.n14926 S.n14925 0.015
R45477 S.n13956 S.n13955 0.015
R45478 S.n12963 S.n12962 0.015
R45479 S.n11958 S.n11957 0.015
R45480 S.n10930 S.n10929 0.015
R45481 S.n9890 S.n9889 0.015
R45482 S.n8827 S.n8826 0.015
R45483 S.n7752 S.n7751 0.015
R45484 S.n6654 S.n6653 0.015
R45485 S.n5544 S.n5543 0.015
R45486 S.n4409 S.n4408 0.015
R45487 S.n3272 S.n3271 0.015
R45488 S.n2120 S.n2119 0.015
R45489 S.n18624 S.n18623 0.015
R45490 S.n17724 S.n17723 0.015
R45491 S.n16797 S.n16796 0.015
R45492 S.n15862 S.n15861 0.015
R45493 S.n14904 S.n14903 0.015
R45494 S.n13934 S.n13933 0.015
R45495 S.n12941 S.n12940 0.015
R45496 S.n11936 S.n11935 0.015
R45497 S.n10908 S.n10907 0.015
R45498 S.n9868 S.n9867 0.015
R45499 S.n8805 S.n8804 0.015
R45500 S.n7730 S.n7729 0.015
R45501 S.n6632 S.n6631 0.015
R45502 S.n5522 S.n5521 0.015
R45503 S.n4387 S.n4386 0.015
R45504 S.n3250 S.n3249 0.015
R45505 S.n2099 S.n2098 0.015
R45506 S.n15949 S.n15948 0.015
R45507 S.n14987 S.n14986 0.015
R45508 S.n14017 S.n14016 0.015
R45509 S.n13024 S.n13023 0.015
R45510 S.n12019 S.n12018 0.015
R45511 S.n10991 S.n10990 0.015
R45512 S.n9951 S.n9950 0.015
R45513 S.n8888 S.n8887 0.015
R45514 S.n7813 S.n7812 0.015
R45515 S.n6715 S.n6714 0.015
R45516 S.n5605 S.n5604 0.015
R45517 S.n4470 S.n4469 0.015
R45518 S.n3332 S.n3331 0.015
R45519 S.n2179 S.n2178 0.015
R45520 S.n16862 S.n16861 0.015
R45521 S.n15927 S.n15926 0.015
R45522 S.n14965 S.n14964 0.015
R45523 S.n13995 S.n13994 0.015
R45524 S.n13002 S.n13001 0.015
R45525 S.n11997 S.n11996 0.015
R45526 S.n10969 S.n10968 0.015
R45527 S.n9929 S.n9928 0.015
R45528 S.n8866 S.n8865 0.015
R45529 S.n7791 S.n7790 0.015
R45530 S.n6693 S.n6692 0.015
R45531 S.n5583 S.n5582 0.015
R45532 S.n4448 S.n4447 0.015
R45533 S.n3310 S.n3309 0.015
R45534 S.n2157 S.n2156 0.015
R45535 S.n14082 S.n14081 0.015
R45536 S.n13085 S.n13084 0.015
R45537 S.n12080 S.n12079 0.015
R45538 S.n11052 S.n11051 0.015
R45539 S.n10012 S.n10011 0.015
R45540 S.n8949 S.n8948 0.015
R45541 S.n7874 S.n7873 0.015
R45542 S.n6776 S.n6775 0.015
R45543 S.n5666 S.n5665 0.015
R45544 S.n4531 S.n4530 0.015
R45545 S.n3392 S.n3391 0.015
R45546 S.n2238 S.n2237 0.015
R45547 S.n15030 S.n15029 0.015
R45548 S.n14060 S.n14059 0.015
R45549 S.n13063 S.n13062 0.015
R45550 S.n12058 S.n12057 0.015
R45551 S.n11030 S.n11029 0.015
R45552 S.n9990 S.n9989 0.015
R45553 S.n8927 S.n8926 0.015
R45554 S.n7852 S.n7851 0.015
R45555 S.n6754 S.n6753 0.015
R45556 S.n5644 S.n5643 0.015
R45557 S.n4509 S.n4508 0.015
R45558 S.n3370 S.n3369 0.015
R45559 S.n2216 S.n2215 0.015
R45560 S.n12145 S.n12144 0.015
R45561 S.n11113 S.n11112 0.015
R45562 S.n10073 S.n10072 0.015
R45563 S.n9010 S.n9009 0.015
R45564 S.n7935 S.n7934 0.015
R45565 S.n6837 S.n6836 0.015
R45566 S.n5727 S.n5726 0.015
R45567 S.n4592 S.n4591 0.015
R45568 S.n3452 S.n3451 0.015
R45569 S.n2297 S.n2296 0.015
R45570 S.n13128 S.n13127 0.015
R45571 S.n12123 S.n12122 0.015
R45572 S.n11091 S.n11090 0.015
R45573 S.n10051 S.n10050 0.015
R45574 S.n8988 S.n8987 0.015
R45575 S.n7913 S.n7912 0.015
R45576 S.n6815 S.n6814 0.015
R45577 S.n5705 S.n5704 0.015
R45578 S.n4570 S.n4569 0.015
R45579 S.n3430 S.n3429 0.015
R45580 S.n2275 S.n2274 0.015
R45581 S.n10138 S.n10137 0.015
R45582 S.n9071 S.n9070 0.015
R45583 S.n7996 S.n7995 0.015
R45584 S.n6898 S.n6897 0.015
R45585 S.n5788 S.n5787 0.015
R45586 S.n4653 S.n4652 0.015
R45587 S.n3512 S.n3511 0.015
R45588 S.n2356 S.n2355 0.015
R45589 S.n11156 S.n11155 0.015
R45590 S.n10116 S.n10115 0.015
R45591 S.n9049 S.n9048 0.015
R45592 S.n7974 S.n7973 0.015
R45593 S.n6876 S.n6875 0.015
R45594 S.n5766 S.n5765 0.015
R45595 S.n4631 S.n4630 0.015
R45596 S.n3490 S.n3489 0.015
R45597 S.n2334 S.n2333 0.015
R45598 S.n8061 S.n8060 0.015
R45599 S.n6959 S.n6958 0.015
R45600 S.n5849 S.n5848 0.015
R45601 S.n4714 S.n4713 0.015
R45602 S.n3572 S.n3571 0.015
R45603 S.n2415 S.n2414 0.015
R45604 S.n9114 S.n9113 0.015
R45605 S.n8039 S.n8038 0.015
R45606 S.n6937 S.n6936 0.015
R45607 S.n5827 S.n5826 0.015
R45608 S.n4692 S.n4691 0.015
R45609 S.n3550 S.n3549 0.015
R45610 S.n2393 S.n2392 0.015
R45611 S.n5914 S.n5913 0.015
R45612 S.n4775 S.n4774 0.015
R45613 S.n3632 S.n3631 0.015
R45614 S.n2474 S.n2473 0.015
R45615 S.n7002 S.n7001 0.015
R45616 S.n5892 S.n5891 0.015
R45617 S.n4753 S.n4752 0.015
R45618 S.n3610 S.n3609 0.015
R45619 S.n2452 S.n2451 0.015
R45620 S.n3696 S.n3695 0.015
R45621 S.n2533 S.n2532 0.015
R45622 S.n4818 S.n4817 0.015
R45623 S.n3674 S.n3673 0.015
R45624 S.n2511 S.n2510 0.015
R45625 S.n2574 S.n2573 0.015
R45626 S.n1352 S.n1351 0.014
R45627 S.n1137 S.n1136 0.014
R45628 S.n1972 S.n1971 0.014
R45629 S.n2124 S.n2123 0.014
R45630 S.n3258 S.n3257 0.014
R45631 S.n4395 S.n4394 0.014
R45632 S.n5530 S.n5529 0.014
R45633 S.n6640 S.n6639 0.014
R45634 S.n7738 S.n7737 0.014
R45635 S.n8813 S.n8812 0.014
R45636 S.n9876 S.n9875 0.014
R45637 S.n10916 S.n10915 0.014
R45638 S.n11944 S.n11943 0.014
R45639 S.n12949 S.n12948 0.014
R45640 S.n13942 S.n13941 0.014
R45641 S.n14912 S.n14911 0.014
R45642 S.n15870 S.n15869 0.014
R45643 S.n16805 S.n16804 0.014
R45644 S.n17732 S.n17731 0.014
R45645 S.n18632 S.n18631 0.014
R45646 S.n2183 S.n2182 0.014
R45647 S.n3318 S.n3317 0.014
R45648 S.n4456 S.n4455 0.014
R45649 S.n5591 S.n5590 0.014
R45650 S.n6701 S.n6700 0.014
R45651 S.n7799 S.n7798 0.014
R45652 S.n8874 S.n8873 0.014
R45653 S.n9937 S.n9936 0.014
R45654 S.n10977 S.n10976 0.014
R45655 S.n12005 S.n12004 0.014
R45656 S.n13010 S.n13009 0.014
R45657 S.n14003 S.n14002 0.014
R45658 S.n14973 S.n14972 0.014
R45659 S.n15935 S.n15934 0.014
R45660 S.n16870 S.n16869 0.014
R45661 S.n2242 S.n2241 0.014
R45662 S.n3378 S.n3377 0.014
R45663 S.n4517 S.n4516 0.014
R45664 S.n5652 S.n5651 0.014
R45665 S.n6762 S.n6761 0.014
R45666 S.n7860 S.n7859 0.014
R45667 S.n8935 S.n8934 0.014
R45668 S.n9998 S.n9997 0.014
R45669 S.n11038 S.n11037 0.014
R45670 S.n12066 S.n12065 0.014
R45671 S.n13071 S.n13070 0.014
R45672 S.n14068 S.n14067 0.014
R45673 S.n15038 S.n15037 0.014
R45674 S.n2301 S.n2300 0.014
R45675 S.n3438 S.n3437 0.014
R45676 S.n4578 S.n4577 0.014
R45677 S.n5713 S.n5712 0.014
R45678 S.n6823 S.n6822 0.014
R45679 S.n7921 S.n7920 0.014
R45680 S.n8996 S.n8995 0.014
R45681 S.n10059 S.n10058 0.014
R45682 S.n11099 S.n11098 0.014
R45683 S.n12131 S.n12130 0.014
R45684 S.n13136 S.n13135 0.014
R45685 S.n2360 S.n2359 0.014
R45686 S.n3498 S.n3497 0.014
R45687 S.n4639 S.n4638 0.014
R45688 S.n5774 S.n5773 0.014
R45689 S.n6884 S.n6883 0.014
R45690 S.n7982 S.n7981 0.014
R45691 S.n9057 S.n9056 0.014
R45692 S.n10124 S.n10123 0.014
R45693 S.n11164 S.n11163 0.014
R45694 S.n2419 S.n2418 0.014
R45695 S.n3558 S.n3557 0.014
R45696 S.n4700 S.n4699 0.014
R45697 S.n5835 S.n5834 0.014
R45698 S.n6945 S.n6944 0.014
R45699 S.n8047 S.n8046 0.014
R45700 S.n9122 S.n9121 0.014
R45701 S.n2478 S.n2477 0.014
R45702 S.n3618 S.n3617 0.014
R45703 S.n4761 S.n4760 0.014
R45704 S.n5900 S.n5899 0.014
R45705 S.n7010 S.n7009 0.014
R45706 S.n2537 S.n2536 0.014
R45707 S.n3682 S.n3681 0.014
R45708 S.n4826 S.n4825 0.014
R45709 S.n2582 S.n2581 0.014
R45710 S.n21995 S.n21986 0.014
R45711 S.n21962 S.n21952 0.014
R45712 S.n1775 S.n1774 0.014
R45713 S.n2074 S.n2073 0.014
R45714 S.n21202 S.n21201 0.013
R45715 S.n20383 S.n20382 0.013
R45716 S.n20256 S.n20255 0.013
R45717 S.n19388 S.n19387 0.013
R45718 S.n18501 S.n18500 0.013
R45719 S.n17601 S.n17600 0.013
R45720 S.n16678 S.n16677 0.013
R45721 S.n15743 S.n15742 0.013
R45722 S.n14785 S.n14784 0.013
R45723 S.n13815 S.n13814 0.013
R45724 S.n12822 S.n12821 0.013
R45725 S.n11817 S.n11816 0.013
R45726 S.n10789 S.n10788 0.013
R45727 S.n9749 S.n9748 0.013
R45728 S.n8686 S.n8685 0.013
R45729 S.n7611 S.n7610 0.013
R45730 S.n6513 S.n6512 0.013
R45731 S.n5402 S.n5401 0.013
R45732 S.n4268 S.n4267 0.013
R45733 S.n3132 S.n3131 0.013
R45734 S.n17750 S.n17749 0.013
R45735 S.n16823 S.n16822 0.013
R45736 S.n15888 S.n15887 0.013
R45737 S.n14930 S.n14929 0.013
R45738 S.n13960 S.n13959 0.013
R45739 S.n12967 S.n12966 0.013
R45740 S.n11962 S.n11961 0.013
R45741 S.n10934 S.n10933 0.013
R45742 S.n9894 S.n9893 0.013
R45743 S.n8831 S.n8830 0.013
R45744 S.n7756 S.n7755 0.013
R45745 S.n6658 S.n6657 0.013
R45746 S.n5548 S.n5547 0.013
R45747 S.n4413 S.n4412 0.013
R45748 S.n3276 S.n3275 0.013
R45749 S.n2106 S.n2105 0.013
R45750 S.n15953 S.n15952 0.013
R45751 S.n14991 S.n14990 0.013
R45752 S.n14021 S.n14020 0.013
R45753 S.n13028 S.n13027 0.013
R45754 S.n12023 S.n12022 0.013
R45755 S.n10995 S.n10994 0.013
R45756 S.n9955 S.n9954 0.013
R45757 S.n8892 S.n8891 0.013
R45758 S.n7817 S.n7816 0.013
R45759 S.n6719 S.n6718 0.013
R45760 S.n5609 S.n5608 0.013
R45761 S.n4474 S.n4473 0.013
R45762 S.n3336 S.n3335 0.013
R45763 S.n2165 S.n2164 0.013
R45764 S.n14086 S.n14085 0.013
R45765 S.n13089 S.n13088 0.013
R45766 S.n12084 S.n12083 0.013
R45767 S.n11056 S.n11055 0.013
R45768 S.n10016 S.n10015 0.013
R45769 S.n8953 S.n8952 0.013
R45770 S.n7878 S.n7877 0.013
R45771 S.n6780 S.n6779 0.013
R45772 S.n5670 S.n5669 0.013
R45773 S.n4535 S.n4534 0.013
R45774 S.n3396 S.n3395 0.013
R45775 S.n2224 S.n2223 0.013
R45776 S.n12149 S.n12148 0.013
R45777 S.n11117 S.n11116 0.013
R45778 S.n10077 S.n10076 0.013
R45779 S.n9014 S.n9013 0.013
R45780 S.n7939 S.n7938 0.013
R45781 S.n6841 S.n6840 0.013
R45782 S.n5731 S.n5730 0.013
R45783 S.n4596 S.n4595 0.013
R45784 S.n3456 S.n3455 0.013
R45785 S.n2283 S.n2282 0.013
R45786 S.n10142 S.n10141 0.013
R45787 S.n9075 S.n9074 0.013
R45788 S.n8000 S.n7999 0.013
R45789 S.n6902 S.n6901 0.013
R45790 S.n5792 S.n5791 0.013
R45791 S.n4657 S.n4656 0.013
R45792 S.n3516 S.n3515 0.013
R45793 S.n2342 S.n2341 0.013
R45794 S.n8065 S.n8064 0.013
R45795 S.n6963 S.n6962 0.013
R45796 S.n5853 S.n5852 0.013
R45797 S.n4718 S.n4717 0.013
R45798 S.n3576 S.n3575 0.013
R45799 S.n2401 S.n2400 0.013
R45800 S.n5918 S.n5917 0.013
R45801 S.n4779 S.n4778 0.013
R45802 S.n3636 S.n3635 0.013
R45803 S.n2460 S.n2459 0.013
R45804 S.n3700 S.n3699 0.013
R45805 S.n2519 S.n2518 0.013
R45806 S.n20421 S.n20420 0.013
R45807 S.n21170 S.n21154 0.013
R45808 S.n1931 S.n1930 0.013
R45809 S.n905 S.n904 0.013
R45810 S.n718 S.n717 0.013
R45811 S.n683 S.n682 0.013
R45812 S.n648 S.n647 0.013
R45813 S.n613 S.n612 0.013
R45814 S.n578 S.n577 0.013
R45815 S.n543 S.n542 0.013
R45816 S.n508 S.n507 0.013
R45817 S.n473 S.n472 0.013
R45818 S.n126 S.n125 0.013
R45819 S.t158 S.n1377 0.012
R45820 S.t158 S.n0 0.012
R45821 S.t158 S.n47 0.012
R45822 S.t158 S.n78 0.012
R45823 S.t158 S.n110 0.012
R45824 S.t158 S.n997 0.012
R45825 S.t158 S.n1029 0.012
R45826 S.t158 S.n1061 0.012
R45827 S.t158 S.n1093 0.012
R45828 S.t158 S.n1125 0.012
R45829 S.t158 S.n1163 0.012
R45830 S.n21199 S.n21198 0.012
R45831 S.n20380 S.n20379 0.012
R45832 S.n20253 S.n20252 0.012
R45833 S.n19385 S.n19384 0.012
R45834 S.n18498 S.n18497 0.012
R45835 S.n17598 S.n17597 0.012
R45836 S.n16675 S.n16674 0.012
R45837 S.n15740 S.n15739 0.012
R45838 S.n14782 S.n14781 0.012
R45839 S.n13812 S.n13811 0.012
R45840 S.n12819 S.n12818 0.012
R45841 S.n11814 S.n11813 0.012
R45842 S.n10786 S.n10785 0.012
R45843 S.n9746 S.n9745 0.012
R45844 S.n8683 S.n8682 0.012
R45845 S.n7608 S.n7607 0.012
R45846 S.n6510 S.n6509 0.012
R45847 S.n5399 S.n5398 0.012
R45848 S.n4265 S.n4264 0.012
R45849 S.n3129 S.n3128 0.012
R45850 S.n1969 S.n1968 0.012
R45851 S.n909 S.n908 0.012
R45852 S.n17747 S.n17746 0.012
R45853 S.n16820 S.n16819 0.012
R45854 S.n15885 S.n15884 0.012
R45855 S.n14927 S.n14926 0.012
R45856 S.n13957 S.n13956 0.012
R45857 S.n12964 S.n12963 0.012
R45858 S.n11959 S.n11958 0.012
R45859 S.n10931 S.n10930 0.012
R45860 S.n9891 S.n9890 0.012
R45861 S.n8828 S.n8827 0.012
R45862 S.n7753 S.n7752 0.012
R45863 S.n6655 S.n6654 0.012
R45864 S.n5545 S.n5544 0.012
R45865 S.n4410 S.n4409 0.012
R45866 S.n3273 S.n3272 0.012
R45867 S.n2121 S.n2120 0.012
R45868 S.n18625 S.n18624 0.012
R45869 S.n17725 S.n17724 0.012
R45870 S.n16798 S.n16797 0.012
R45871 S.n15863 S.n15862 0.012
R45872 S.n14905 S.n14904 0.012
R45873 S.n13935 S.n13934 0.012
R45874 S.n12942 S.n12941 0.012
R45875 S.n11937 S.n11936 0.012
R45876 S.n10909 S.n10908 0.012
R45877 S.n9869 S.n9868 0.012
R45878 S.n8806 S.n8805 0.012
R45879 S.n7731 S.n7730 0.012
R45880 S.n6633 S.n6632 0.012
R45881 S.n5523 S.n5522 0.012
R45882 S.n4388 S.n4387 0.012
R45883 S.n3251 S.n3250 0.012
R45884 S.n2067 S.n2066 0.012
R45885 S.n19472 S.n19471 0.012
R45886 S.n18582 S.n18581 0.012
R45887 S.n17682 S.n17681 0.012
R45888 S.n16759 S.n16758 0.012
R45889 S.n15824 S.n15823 0.012
R45890 S.n14866 S.n14865 0.012
R45891 S.n13896 S.n13895 0.012
R45892 S.n12903 S.n12902 0.012
R45893 S.n11898 S.n11897 0.012
R45894 S.n10870 S.n10869 0.012
R45895 S.n9830 S.n9829 0.012
R45896 S.n8767 S.n8766 0.012
R45897 S.n7692 S.n7691 0.012
R45898 S.n6594 S.n6593 0.012
R45899 S.n5484 S.n5483 0.012
R45900 S.n4349 S.n4348 0.012
R45901 S.n3213 S.n3212 0.012
R45902 S.n2100 S.n2099 0.012
R45903 S.n387 S.n386 0.012
R45904 S.n15950 S.n15949 0.012
R45905 S.n14988 S.n14987 0.012
R45906 S.n14018 S.n14017 0.012
R45907 S.n13025 S.n13024 0.012
R45908 S.n12020 S.n12019 0.012
R45909 S.n10992 S.n10991 0.012
R45910 S.n9952 S.n9951 0.012
R45911 S.n8889 S.n8888 0.012
R45912 S.n7814 S.n7813 0.012
R45913 S.n6716 S.n6715 0.012
R45914 S.n5606 S.n5605 0.012
R45915 S.n4471 S.n4470 0.012
R45916 S.n3333 S.n3332 0.012
R45917 S.n2180 S.n2179 0.012
R45918 S.n16863 S.n16862 0.012
R45919 S.n15928 S.n15927 0.012
R45920 S.n14966 S.n14965 0.012
R45921 S.n13996 S.n13995 0.012
R45922 S.n13003 S.n13002 0.012
R45923 S.n11998 S.n11997 0.012
R45924 S.n10970 S.n10969 0.012
R45925 S.n9930 S.n9929 0.012
R45926 S.n8867 S.n8866 0.012
R45927 S.n7792 S.n7791 0.012
R45928 S.n6694 S.n6693 0.012
R45929 S.n5584 S.n5583 0.012
R45930 S.n4449 S.n4448 0.012
R45931 S.n3311 S.n3310 0.012
R45932 S.n2158 S.n2157 0.012
R45933 S.n355 S.n354 0.012
R45934 S.n14083 S.n14082 0.012
R45935 S.n13086 S.n13085 0.012
R45936 S.n12081 S.n12080 0.012
R45937 S.n11053 S.n11052 0.012
R45938 S.n10013 S.n10012 0.012
R45939 S.n8950 S.n8949 0.012
R45940 S.n7875 S.n7874 0.012
R45941 S.n6777 S.n6776 0.012
R45942 S.n5667 S.n5666 0.012
R45943 S.n4532 S.n4531 0.012
R45944 S.n3393 S.n3392 0.012
R45945 S.n2239 S.n2238 0.012
R45946 S.n15031 S.n15030 0.012
R45947 S.n14061 S.n14060 0.012
R45948 S.n13064 S.n13063 0.012
R45949 S.n12059 S.n12058 0.012
R45950 S.n11031 S.n11030 0.012
R45951 S.n9991 S.n9990 0.012
R45952 S.n8928 S.n8927 0.012
R45953 S.n7853 S.n7852 0.012
R45954 S.n6755 S.n6754 0.012
R45955 S.n5645 S.n5644 0.012
R45956 S.n4510 S.n4509 0.012
R45957 S.n3371 S.n3370 0.012
R45958 S.n2217 S.n2216 0.012
R45959 S.n323 S.n322 0.012
R45960 S.n12146 S.n12145 0.012
R45961 S.n11114 S.n11113 0.012
R45962 S.n10074 S.n10073 0.012
R45963 S.n9011 S.n9010 0.012
R45964 S.n7936 S.n7935 0.012
R45965 S.n6838 S.n6837 0.012
R45966 S.n5728 S.n5727 0.012
R45967 S.n4593 S.n4592 0.012
R45968 S.n3453 S.n3452 0.012
R45969 S.n2298 S.n2297 0.012
R45970 S.n13129 S.n13128 0.012
R45971 S.n12124 S.n12123 0.012
R45972 S.n11092 S.n11091 0.012
R45973 S.n10052 S.n10051 0.012
R45974 S.n8989 S.n8988 0.012
R45975 S.n7914 S.n7913 0.012
R45976 S.n6816 S.n6815 0.012
R45977 S.n5706 S.n5705 0.012
R45978 S.n4571 S.n4570 0.012
R45979 S.n3431 S.n3430 0.012
R45980 S.n2276 S.n2275 0.012
R45981 S.n291 S.n290 0.012
R45982 S.n10139 S.n10138 0.012
R45983 S.n9072 S.n9071 0.012
R45984 S.n7997 S.n7996 0.012
R45985 S.n6899 S.n6898 0.012
R45986 S.n5789 S.n5788 0.012
R45987 S.n4654 S.n4653 0.012
R45988 S.n3513 S.n3512 0.012
R45989 S.n2357 S.n2356 0.012
R45990 S.n11157 S.n11156 0.012
R45991 S.n10117 S.n10116 0.012
R45992 S.n9050 S.n9049 0.012
R45993 S.n7975 S.n7974 0.012
R45994 S.n6877 S.n6876 0.012
R45995 S.n5767 S.n5766 0.012
R45996 S.n4632 S.n4631 0.012
R45997 S.n3491 S.n3490 0.012
R45998 S.n2335 S.n2334 0.012
R45999 S.n259 S.n258 0.012
R46000 S.n8062 S.n8061 0.012
R46001 S.n6960 S.n6959 0.012
R46002 S.n5850 S.n5849 0.012
R46003 S.n4715 S.n4714 0.012
R46004 S.n3573 S.n3572 0.012
R46005 S.n2416 S.n2415 0.012
R46006 S.n9115 S.n9114 0.012
R46007 S.n8040 S.n8039 0.012
R46008 S.n6938 S.n6937 0.012
R46009 S.n5828 S.n5827 0.012
R46010 S.n4693 S.n4692 0.012
R46011 S.n3551 S.n3550 0.012
R46012 S.n2394 S.n2393 0.012
R46013 S.n230 S.n229 0.012
R46014 S.n5915 S.n5914 0.012
R46015 S.n4776 S.n4775 0.012
R46016 S.n3633 S.n3632 0.012
R46017 S.n2475 S.n2474 0.012
R46018 S.n7003 S.n7002 0.012
R46019 S.n5893 S.n5892 0.012
R46020 S.n4754 S.n4753 0.012
R46021 S.n3611 S.n3610 0.012
R46022 S.n2453 S.n2452 0.012
R46023 S.n195 S.n194 0.012
R46024 S.n3697 S.n3696 0.012
R46025 S.n2534 S.n2533 0.012
R46026 S.n4819 S.n4818 0.012
R46027 S.n3675 S.n3674 0.012
R46028 S.n2512 S.n2511 0.012
R46029 S.n163 S.n162 0.012
R46030 S.n2575 S.n2574 0.012
R46031 S.n22988 S.n22987 0.012
R46032 S.n23004 S.n23003 0.012
R46033 S.n889 S.n888 0.011
R46034 S.n914 S.n902 0.011
R46035 S.n1140 S.n1139 0.011
R46036 S.n22328 S.n22325 0.011
R46037 S.n21154 S.n21153 0.011
R46038 S.n20326 S.n20316 0.011
R46039 S.n19454 S.n19444 0.011
R46040 S.n1141 S.n1140 0.01
R46041 S.n21638 S.n21626 0.01
R46042 S.n20818 S.n20803 0.01
R46043 S.n734 S.n733 0.01
R46044 S.n699 S.n698 0.01
R46045 S.n664 S.n663 0.01
R46046 S.n629 S.n628 0.01
R46047 S.n594 S.n593 0.01
R46048 S.n559 S.n558 0.01
R46049 S.n524 S.n523 0.01
R46050 S.n489 S.n488 0.01
R46051 S.n20219 S.n20218 0.01
R46052 S.n21172 S.n20348 0.01
R46053 S.n20344 S.n19522 0.01
R46054 S.n19504 S.n18665 0.01
R46055 S.n18647 S.n17797 0.01
R46056 S.n17779 S.n16903 0.01
R46057 S.n16885 S.n16000 0.01
R46058 S.n15982 S.n15071 0.01
R46059 S.n15053 S.n14133 0.01
R46060 S.n14115 S.n13169 0.01
R46061 S.n13151 S.n12196 0.01
R46062 S.n12178 S.n11197 0.01
R46063 S.n11179 S.n10189 0.01
R46064 S.n10171 S.n9155 0.01
R46065 S.n9137 S.n8112 0.01
R46066 S.n8094 S.n7043 0.01
R46067 S.n7025 S.n5965 0.01
R46068 S.n5947 S.n4860 0.01
R46069 S.n4841 S.n3747 0.01
R46070 S.n3728 S.n2617 0.01
R46071 S.n2597 S.n1914 0.01
R46072 S.n2597 S.n1917 0.01
R46073 S.n806 S.n803 0.01
R46074 S.n914 S.n913 0.01
R46075 S.n838 S.n836 0.01
R46076 S.n1823 S.n1815 0.01
R46077 S.n2986 S.n2978 0.01
R46078 S.n4113 S.n4105 0.01
R46079 S.n5225 S.n5217 0.01
R46080 S.n6325 S.n6317 0.01
R46081 S.n7402 S.n7394 0.01
R46082 S.n8466 S.n8458 0.01
R46083 S.n9508 S.n9500 0.01
R46084 S.n10537 S.n10529 0.01
R46085 S.n11544 S.n11536 0.01
R46086 S.n12538 S.n12530 0.01
R46087 S.n13510 S.n13502 0.01
R46088 S.n14469 S.n14461 0.01
R46089 S.n15406 S.n15398 0.01
R46090 S.n16330 S.n16322 0.01
R46091 S.n17232 S.n17224 0.01
R46092 S.n18121 S.n18113 0.01
R46093 S.n18987 S.n18978 0.01
R46094 S.n19839 S.n19830 0.01
R46095 S.n767 S.n763 0.01
R46096 S.n20472 S.n20468 0.01
R46097 S.n19861 S.n19857 0.01
R46098 S.n19007 S.n19003 0.01
R46099 S.n18141 S.n18137 0.01
R46100 S.n17252 S.n17248 0.01
R46101 S.n16350 S.n16346 0.01
R46102 S.n15426 S.n15422 0.01
R46103 S.n14489 S.n14485 0.01
R46104 S.n13530 S.n13526 0.01
R46105 S.n12558 S.n12554 0.01
R46106 S.n11564 S.n11560 0.01
R46107 S.n10557 S.n10553 0.01
R46108 S.n9528 S.n9524 0.01
R46109 S.n8486 S.n8482 0.01
R46110 S.n7422 S.n7418 0.01
R46111 S.n6345 S.n6341 0.01
R46112 S.n5245 S.n5241 0.01
R46113 S.n4132 S.n4129 0.01
R46114 S.n3006 S.n3002 0.01
R46115 S.n1845 S.n1836 0.01
R46116 S.n786 S.n783 0.01
R46117 S.n406 S.n397 0.01
R46118 S.n406 S.n391 0.01
R46119 S.n374 S.n365 0.01
R46120 S.n374 S.n359 0.01
R46121 S.n342 S.n333 0.01
R46122 S.n342 S.n327 0.01
R46123 S.n310 S.n301 0.01
R46124 S.n310 S.n295 0.01
R46125 S.n278 S.n269 0.01
R46126 S.n278 S.n263 0.01
R46127 S.n249 S.n240 0.01
R46128 S.n249 S.n234 0.01
R46129 S.n214 S.n205 0.01
R46130 S.n214 S.n199 0.01
R46131 S.n182 S.n173 0.01
R46132 S.n182 S.n167 0.01
R46133 S.n150 S.n141 0.01
R46134 S.n150 S.n135 0.01
R46135 S.n21980 S.n21977 0.01
R46136 S.n22307 S.n22300 0.01
R46137 S.n22328 S.n22322 0.01
R46138 S.n1798 S.n1796 0.01
R46139 S.n20451 S.n20440 0.01
R46140 S.n18943 S.n18931 0.01
R46141 S.n17151 S.n17139 0.01
R46142 S.n15289 S.n15277 0.01
R46143 S.n13357 S.n13345 0.01
R46144 S.n11355 S.n11343 0.01
R46145 S.n9283 S.n9271 0.01
R46146 S.n7141 S.n7129 0.01
R46147 S.n4928 S.n4916 0.01
R46148 S.n2653 S.n2641 0.01
R46149 S.n21980 S.n21190 0.009
R46150 S.n22791 S.n21981 0.009
R46151 S.n1136 S.n1135 0.009
R46152 S.n22694 S.n22693 0.009
R46153 S.n22713 S.n22704 0.009
R46154 S.n21261 S.n21252 0.009
R46155 S.n20424 S.n20423 0.009
R46156 S.n20329 S.n20327 0.009
R46157 S.n20330 S.n20329 0.009
R46158 S.n19457 S.n19455 0.009
R46159 S.n19458 S.n19457 0.009
R46160 S.n717 S.n716 0.009
R46161 S.n682 S.n681 0.009
R46162 S.n647 S.n646 0.009
R46163 S.n612 S.n611 0.009
R46164 S.n577 S.n576 0.009
R46165 S.n542 S.n541 0.009
R46166 S.n507 S.n506 0.009
R46167 S.n472 S.n471 0.009
R46168 S.n912 S.n911 0.008
R46169 S.n390 S.n389 0.008
R46170 S.n358 S.n357 0.008
R46171 S.n326 S.n325 0.008
R46172 S.n294 S.n293 0.008
R46173 S.n262 S.n261 0.008
R46174 S.n233 S.n232 0.008
R46175 S.n198 S.n197 0.008
R46176 S.n166 S.n165 0.008
R46177 S.n134 S.n133 0.008
R46178 S.n22299 S.n22298 0.008
R46179 S.n22321 S.n22320 0.008
R46180 S.n22991 S.n22989 0.008
R46181 S.n23006 S.n23005 0.008
R46182 S.n21200 S.n21199 0.008
R46183 S.n20381 S.n20380 0.008
R46184 S.n20254 S.n20253 0.008
R46185 S.n19386 S.n19385 0.008
R46186 S.n18499 S.n18498 0.008
R46187 S.n17599 S.n17598 0.008
R46188 S.n16676 S.n16675 0.008
R46189 S.n15741 S.n15740 0.008
R46190 S.n14783 S.n14782 0.008
R46191 S.n13813 S.n13812 0.008
R46192 S.n12820 S.n12819 0.008
R46193 S.n11815 S.n11814 0.008
R46194 S.n10787 S.n10786 0.008
R46195 S.n9747 S.n9746 0.008
R46196 S.n8684 S.n8683 0.008
R46197 S.n7609 S.n7608 0.008
R46198 S.n6511 S.n6510 0.008
R46199 S.n5400 S.n5399 0.008
R46200 S.n4266 S.n4265 0.008
R46201 S.n3130 S.n3129 0.008
R46202 S.n1970 S.n1969 0.008
R46203 S.n17748 S.n17747 0.008
R46204 S.n16821 S.n16820 0.008
R46205 S.n15886 S.n15885 0.008
R46206 S.n14928 S.n14927 0.008
R46207 S.n13958 S.n13957 0.008
R46208 S.n12965 S.n12964 0.008
R46209 S.n11960 S.n11959 0.008
R46210 S.n10932 S.n10931 0.008
R46211 S.n9892 S.n9891 0.008
R46212 S.n8829 S.n8828 0.008
R46213 S.n7754 S.n7753 0.008
R46214 S.n6656 S.n6655 0.008
R46215 S.n5546 S.n5545 0.008
R46216 S.n4411 S.n4410 0.008
R46217 S.n3274 S.n3273 0.008
R46218 S.n2122 S.n2121 0.008
R46219 S.n18626 S.n18625 0.008
R46220 S.n17726 S.n17725 0.008
R46221 S.n16799 S.n16798 0.008
R46222 S.n15864 S.n15863 0.008
R46223 S.n14906 S.n14905 0.008
R46224 S.n13936 S.n13935 0.008
R46225 S.n12943 S.n12942 0.008
R46226 S.n11938 S.n11937 0.008
R46227 S.n10910 S.n10909 0.008
R46228 S.n9870 S.n9869 0.008
R46229 S.n8807 S.n8806 0.008
R46230 S.n7732 S.n7731 0.008
R46231 S.n6634 S.n6633 0.008
R46232 S.n5524 S.n5523 0.008
R46233 S.n4389 S.n4388 0.008
R46234 S.n3252 S.n3251 0.008
R46235 S.n2101 S.n2100 0.008
R46236 S.n15951 S.n15950 0.008
R46237 S.n14989 S.n14988 0.008
R46238 S.n14019 S.n14018 0.008
R46239 S.n13026 S.n13025 0.008
R46240 S.n12021 S.n12020 0.008
R46241 S.n10993 S.n10992 0.008
R46242 S.n9953 S.n9952 0.008
R46243 S.n8890 S.n8889 0.008
R46244 S.n7815 S.n7814 0.008
R46245 S.n6717 S.n6716 0.008
R46246 S.n5607 S.n5606 0.008
R46247 S.n4472 S.n4471 0.008
R46248 S.n3334 S.n3333 0.008
R46249 S.n2181 S.n2180 0.008
R46250 S.n16864 S.n16863 0.008
R46251 S.n15929 S.n15928 0.008
R46252 S.n14967 S.n14966 0.008
R46253 S.n13997 S.n13996 0.008
R46254 S.n13004 S.n13003 0.008
R46255 S.n11999 S.n11998 0.008
R46256 S.n10971 S.n10970 0.008
R46257 S.n9931 S.n9930 0.008
R46258 S.n8868 S.n8867 0.008
R46259 S.n7793 S.n7792 0.008
R46260 S.n6695 S.n6694 0.008
R46261 S.n5585 S.n5584 0.008
R46262 S.n4450 S.n4449 0.008
R46263 S.n3312 S.n3311 0.008
R46264 S.n2159 S.n2158 0.008
R46265 S.n14084 S.n14083 0.008
R46266 S.n13087 S.n13086 0.008
R46267 S.n12082 S.n12081 0.008
R46268 S.n11054 S.n11053 0.008
R46269 S.n10014 S.n10013 0.008
R46270 S.n8951 S.n8950 0.008
R46271 S.n7876 S.n7875 0.008
R46272 S.n6778 S.n6777 0.008
R46273 S.n5668 S.n5667 0.008
R46274 S.n4533 S.n4532 0.008
R46275 S.n3394 S.n3393 0.008
R46276 S.n2240 S.n2239 0.008
R46277 S.n15032 S.n15031 0.008
R46278 S.n14062 S.n14061 0.008
R46279 S.n13065 S.n13064 0.008
R46280 S.n12060 S.n12059 0.008
R46281 S.n11032 S.n11031 0.008
R46282 S.n9992 S.n9991 0.008
R46283 S.n8929 S.n8928 0.008
R46284 S.n7854 S.n7853 0.008
R46285 S.n6756 S.n6755 0.008
R46286 S.n5646 S.n5645 0.008
R46287 S.n4511 S.n4510 0.008
R46288 S.n3372 S.n3371 0.008
R46289 S.n2218 S.n2217 0.008
R46290 S.n12147 S.n12146 0.008
R46291 S.n11115 S.n11114 0.008
R46292 S.n10075 S.n10074 0.008
R46293 S.n9012 S.n9011 0.008
R46294 S.n7937 S.n7936 0.008
R46295 S.n6839 S.n6838 0.008
R46296 S.n5729 S.n5728 0.008
R46297 S.n4594 S.n4593 0.008
R46298 S.n3454 S.n3453 0.008
R46299 S.n2299 S.n2298 0.008
R46300 S.n13130 S.n13129 0.008
R46301 S.n12125 S.n12124 0.008
R46302 S.n11093 S.n11092 0.008
R46303 S.n10053 S.n10052 0.008
R46304 S.n8990 S.n8989 0.008
R46305 S.n7915 S.n7914 0.008
R46306 S.n6817 S.n6816 0.008
R46307 S.n5707 S.n5706 0.008
R46308 S.n4572 S.n4571 0.008
R46309 S.n3432 S.n3431 0.008
R46310 S.n2277 S.n2276 0.008
R46311 S.n10140 S.n10139 0.008
R46312 S.n9073 S.n9072 0.008
R46313 S.n7998 S.n7997 0.008
R46314 S.n6900 S.n6899 0.008
R46315 S.n5790 S.n5789 0.008
R46316 S.n4655 S.n4654 0.008
R46317 S.n3514 S.n3513 0.008
R46318 S.n2358 S.n2357 0.008
R46319 S.n11158 S.n11157 0.008
R46320 S.n10118 S.n10117 0.008
R46321 S.n9051 S.n9050 0.008
R46322 S.n7976 S.n7975 0.008
R46323 S.n6878 S.n6877 0.008
R46324 S.n5768 S.n5767 0.008
R46325 S.n4633 S.n4632 0.008
R46326 S.n3492 S.n3491 0.008
R46327 S.n2336 S.n2335 0.008
R46328 S.n8063 S.n8062 0.008
R46329 S.n6961 S.n6960 0.008
R46330 S.n5851 S.n5850 0.008
R46331 S.n4716 S.n4715 0.008
R46332 S.n3574 S.n3573 0.008
R46333 S.n2417 S.n2416 0.008
R46334 S.n9116 S.n9115 0.008
R46335 S.n8041 S.n8040 0.008
R46336 S.n6939 S.n6938 0.008
R46337 S.n5829 S.n5828 0.008
R46338 S.n4694 S.n4693 0.008
R46339 S.n3552 S.n3551 0.008
R46340 S.n2395 S.n2394 0.008
R46341 S.n5916 S.n5915 0.008
R46342 S.n4777 S.n4776 0.008
R46343 S.n3634 S.n3633 0.008
R46344 S.n2476 S.n2475 0.008
R46345 S.n7004 S.n7003 0.008
R46346 S.n5894 S.n5893 0.008
R46347 S.n4755 S.n4754 0.008
R46348 S.n3612 S.n3611 0.008
R46349 S.n2454 S.n2453 0.008
R46350 S.n3698 S.n3697 0.008
R46351 S.n2535 S.n2534 0.008
R46352 S.n4820 S.n4819 0.008
R46353 S.n3676 S.n3675 0.008
R46354 S.n2513 S.n2512 0.008
R46355 S.n2576 S.n2575 0.008
R46356 S.n20818 S.n20817 0.008
R46357 S.n1984 S.n1983 0.008
R46358 S.n1864 S.n1863 0.008
R46359 S.n3145 S.n3144 0.008
R46360 S.n3024 S.n3023 0.008
R46361 S.n4282 S.n4281 0.008
R46362 S.n4150 S.n4149 0.008
R46363 S.n5416 S.n5415 0.008
R46364 S.n5263 S.n5262 0.008
R46365 S.n6527 S.n6526 0.008
R46366 S.n6363 S.n6362 0.008
R46367 S.n7625 S.n7624 0.008
R46368 S.n7440 S.n7439 0.008
R46369 S.n8700 S.n8699 0.008
R46370 S.n8504 S.n8503 0.008
R46371 S.n9763 S.n9762 0.008
R46372 S.n9546 S.n9545 0.008
R46373 S.n10803 S.n10802 0.008
R46374 S.n10575 S.n10574 0.008
R46375 S.n11831 S.n11830 0.008
R46376 S.n11582 S.n11581 0.008
R46377 S.n12836 S.n12835 0.008
R46378 S.n12576 S.n12575 0.008
R46379 S.n13829 S.n13828 0.008
R46380 S.n13548 S.n13547 0.008
R46381 S.n14799 S.n14798 0.008
R46382 S.n14507 S.n14506 0.008
R46383 S.n15757 S.n15756 0.008
R46384 S.n15444 S.n15443 0.008
R46385 S.n16692 S.n16691 0.008
R46386 S.n16368 S.n16367 0.008
R46387 S.n17615 S.n17614 0.008
R46388 S.n17270 S.n17269 0.008
R46389 S.n18515 S.n18514 0.008
R46390 S.n18159 S.n18158 0.008
R46391 S.n19402 S.n19401 0.008
R46392 S.n19025 S.n19024 0.008
R46393 S.n20270 S.n20269 0.008
R46394 S.n19879 S.n19878 0.008
R46395 S.n20490 S.n20489 0.008
R46396 S.n21313 S.n21312 0.008
R46397 S.n974 S.n950 0.008
R46398 S.n806 S.n805 0.008
R46399 S.n2053 S.n2052 0.008
R46400 S.n1784 S.n1783 0.008
R46401 S.n3229 S.n3228 0.008
R46402 S.n2960 S.n2959 0.008
R46403 S.n4366 S.n4365 0.008
R46404 S.n4087 S.n4086 0.008
R46405 S.n5501 S.n5500 0.008
R46406 S.n5199 S.n5198 0.008
R46407 S.n6611 S.n6610 0.008
R46408 S.n6299 S.n6298 0.008
R46409 S.n7709 S.n7708 0.008
R46410 S.n7376 S.n7375 0.008
R46411 S.n8784 S.n8783 0.008
R46412 S.n8440 S.n8439 0.008
R46413 S.n9847 S.n9846 0.008
R46414 S.n9482 S.n9481 0.008
R46415 S.n10887 S.n10886 0.008
R46416 S.n10511 S.n10510 0.008
R46417 S.n11915 S.n11914 0.008
R46418 S.n11518 S.n11517 0.008
R46419 S.n12920 S.n12919 0.008
R46420 S.n12512 S.n12511 0.008
R46421 S.n13913 S.n13912 0.008
R46422 S.n13484 S.n13483 0.008
R46423 S.n14883 S.n14882 0.008
R46424 S.n14443 S.n14442 0.008
R46425 S.n15841 S.n15840 0.008
R46426 S.n15380 S.n15379 0.008
R46427 S.n16776 S.n16775 0.008
R46428 S.n16304 S.n16303 0.008
R46429 S.n17699 S.n17698 0.008
R46430 S.n17206 S.n17205 0.008
R46431 S.n18095 S.n18094 0.008
R46432 S.n18960 S.n18959 0.008
R46433 S.n1823 S.n1810 0.008
R46434 S.n2986 S.n2972 0.008
R46435 S.n4113 S.n4099 0.008
R46436 S.n5225 S.n5211 0.008
R46437 S.n6325 S.n6311 0.008
R46438 S.n7402 S.n7388 0.008
R46439 S.n8466 S.n8452 0.008
R46440 S.n9508 S.n9494 0.008
R46441 S.n10537 S.n10523 0.008
R46442 S.n11544 S.n11530 0.008
R46443 S.n12538 S.n12524 0.008
R46444 S.n13510 S.n13496 0.008
R46445 S.n14469 S.n14455 0.008
R46446 S.n15406 S.n15392 0.008
R46447 S.n16330 S.n16316 0.008
R46448 S.n17232 S.n17218 0.008
R46449 S.n18121 S.n18107 0.008
R46450 S.n18987 S.n18972 0.008
R46451 S.n19839 S.n19824 0.008
R46452 S.n1336 S.n1335 0.008
R46453 S.n767 S.n766 0.008
R46454 S.n20472 S.n20471 0.008
R46455 S.n19861 S.n19860 0.008
R46456 S.n19007 S.n19006 0.008
R46457 S.n18141 S.n18140 0.008
R46458 S.n17252 S.n17251 0.008
R46459 S.n16350 S.n16349 0.008
R46460 S.n15426 S.n15425 0.008
R46461 S.n14489 S.n14488 0.008
R46462 S.n13530 S.n13529 0.008
R46463 S.n12558 S.n12557 0.008
R46464 S.n11564 S.n11563 0.008
R46465 S.n10557 S.n10556 0.008
R46466 S.n9528 S.n9527 0.008
R46467 S.n8486 S.n8485 0.008
R46468 S.n7422 S.n7421 0.008
R46469 S.n6345 S.n6344 0.008
R46470 S.n5245 S.n5244 0.008
R46471 S.n4132 S.n4131 0.008
R46472 S.n3006 S.n3005 0.008
R46473 S.n1845 S.n1834 0.008
R46474 S.n1993 S.n1992 0.008
R46475 S.n3154 S.n3153 0.008
R46476 S.n4291 S.n4290 0.008
R46477 S.n5425 S.n5424 0.008
R46478 S.n6536 S.n6535 0.008
R46479 S.n7634 S.n7633 0.008
R46480 S.n8709 S.n8708 0.008
R46481 S.n9772 S.n9771 0.008
R46482 S.n10812 S.n10811 0.008
R46483 S.n11840 S.n11839 0.008
R46484 S.n12845 S.n12844 0.008
R46485 S.n13838 S.n13837 0.008
R46486 S.n14808 S.n14807 0.008
R46487 S.n15766 S.n15765 0.008
R46488 S.n16701 S.n16700 0.008
R46489 S.n17624 S.n17623 0.008
R46490 S.n18524 S.n18523 0.008
R46491 S.n19411 S.n19410 0.008
R46492 S.n848 S.n847 0.008
R46493 S.n862 S.n858 0.008
R46494 S.n862 S.n861 0.008
R46495 S.n786 S.n785 0.008
R46496 S.n19369 S.n19367 0.008
R46497 S.n16785 S.n16784 0.008
R46498 S.n15850 S.n15849 0.008
R46499 S.n14892 S.n14891 0.008
R46500 S.n13922 S.n13921 0.008
R46501 S.n12929 S.n12928 0.008
R46502 S.n11924 S.n11923 0.008
R46503 S.n10896 S.n10895 0.008
R46504 S.n9856 S.n9855 0.008
R46505 S.n8793 S.n8792 0.008
R46506 S.n7718 S.n7717 0.008
R46507 S.n6620 S.n6619 0.008
R46508 S.n5510 S.n5509 0.008
R46509 S.n4375 S.n4374 0.008
R46510 S.n3238 S.n3237 0.008
R46511 S.n2088 S.n2087 0.008
R46512 S.n8 S.n5 0.008
R46513 S.n2136 S.n2135 0.008
R46514 S.n1756 S.n1755 0.008
R46515 S.n3289 S.n3288 0.008
R46516 S.n2924 S.n2923 0.008
R46517 S.n4427 S.n4426 0.008
R46518 S.n4051 S.n4050 0.008
R46519 S.n5562 S.n5561 0.008
R46520 S.n5163 S.n5162 0.008
R46521 S.n6672 S.n6671 0.008
R46522 S.n6263 S.n6262 0.008
R46523 S.n7770 S.n7769 0.008
R46524 S.n7340 S.n7339 0.008
R46525 S.n8845 S.n8844 0.008
R46526 S.n8404 S.n8403 0.008
R46527 S.n9908 S.n9907 0.008
R46528 S.n9446 S.n9445 0.008
R46529 S.n10948 S.n10947 0.008
R46530 S.n10475 S.n10474 0.008
R46531 S.n11976 S.n11975 0.008
R46532 S.n11482 S.n11481 0.008
R46533 S.n12981 S.n12980 0.008
R46534 S.n12476 S.n12475 0.008
R46535 S.n13974 S.n13973 0.008
R46536 S.n13448 S.n13447 0.008
R46537 S.n14944 S.n14943 0.008
R46538 S.n14407 S.n14406 0.008
R46539 S.n15902 S.n15901 0.008
R46540 S.n15344 S.n15343 0.008
R46541 S.n16268 S.n16267 0.008
R46542 S.n17168 S.n17167 0.008
R46543 S.n17582 S.n17580 0.008
R46544 S.n14953 S.n14952 0.008
R46545 S.n13983 S.n13982 0.008
R46546 S.n12990 S.n12989 0.008
R46547 S.n11985 S.n11984 0.008
R46548 S.n10957 S.n10956 0.008
R46549 S.n9917 S.n9916 0.008
R46550 S.n8854 S.n8853 0.008
R46551 S.n7779 S.n7778 0.008
R46552 S.n6681 S.n6680 0.008
R46553 S.n5571 S.n5570 0.008
R46554 S.n4436 S.n4435 0.008
R46555 S.n3298 S.n3297 0.008
R46556 S.n2146 S.n2145 0.008
R46557 S.n55 S.n52 0.008
R46558 S.n2195 S.n2194 0.008
R46559 S.n1719 S.n1718 0.008
R46560 S.n3349 S.n3348 0.008
R46561 S.n2888 S.n2887 0.008
R46562 S.n4488 S.n4487 0.008
R46563 S.n4015 S.n4014 0.008
R46564 S.n5623 S.n5622 0.008
R46565 S.n5127 S.n5126 0.008
R46566 S.n6733 S.n6732 0.008
R46567 S.n6227 S.n6226 0.008
R46568 S.n7831 S.n7830 0.008
R46569 S.n7304 S.n7303 0.008
R46570 S.n8906 S.n8905 0.008
R46571 S.n8368 S.n8367 0.008
R46572 S.n9969 S.n9968 0.008
R46573 S.n9410 S.n9409 0.008
R46574 S.n11009 S.n11008 0.008
R46575 S.n10439 S.n10438 0.008
R46576 S.n12037 S.n12036 0.008
R46577 S.n11446 S.n11445 0.008
R46578 S.n13042 S.n13041 0.008
R46579 S.n12440 S.n12439 0.008
R46580 S.n14035 S.n14034 0.008
R46581 S.n13412 S.n13411 0.008
R46582 S.n14371 S.n14370 0.008
R46583 S.n15306 S.n15305 0.008
R46584 S.n15724 S.n15720 0.008
R46585 S.n13051 S.n13050 0.008
R46586 S.n12046 S.n12045 0.008
R46587 S.n11018 S.n11017 0.008
R46588 S.n9978 S.n9977 0.008
R46589 S.n8915 S.n8914 0.008
R46590 S.n7840 S.n7839 0.008
R46591 S.n6742 S.n6741 0.008
R46592 S.n5632 S.n5631 0.008
R46593 S.n4497 S.n4496 0.008
R46594 S.n3358 S.n3357 0.008
R46595 S.n2205 S.n2204 0.008
R46596 S.n85 S.n84 0.008
R46597 S.n2254 S.n2253 0.008
R46598 S.n1682 S.n1681 0.008
R46599 S.n3409 S.n3408 0.008
R46600 S.n2852 S.n2851 0.008
R46601 S.n4549 S.n4548 0.008
R46602 S.n3979 S.n3978 0.008
R46603 S.n5684 S.n5683 0.008
R46604 S.n5091 S.n5090 0.008
R46605 S.n6794 S.n6793 0.008
R46606 S.n6191 S.n6190 0.008
R46607 S.n7892 S.n7891 0.008
R46608 S.n7268 S.n7267 0.008
R46609 S.n8967 S.n8966 0.008
R46610 S.n8332 S.n8331 0.008
R46611 S.n10030 S.n10029 0.008
R46612 S.n9374 S.n9373 0.008
R46613 S.n11070 S.n11069 0.008
R46614 S.n10403 S.n10402 0.008
R46615 S.n12098 S.n12097 0.008
R46616 S.n11410 S.n11409 0.008
R46617 S.n12404 S.n12403 0.008
R46618 S.n13374 S.n13373 0.008
R46619 S.n13796 S.n13792 0.008
R46620 S.n11079 S.n11078 0.008
R46621 S.n10039 S.n10038 0.008
R46622 S.n8976 S.n8975 0.008
R46623 S.n7901 S.n7900 0.008
R46624 S.n6803 S.n6802 0.008
R46625 S.n5693 S.n5692 0.008
R46626 S.n4558 S.n4557 0.008
R46627 S.n3418 S.n3417 0.008
R46628 S.n2264 S.n2263 0.008
R46629 S.n119 S.n116 0.008
R46630 S.n2313 S.n2312 0.008
R46631 S.n1645 S.n1644 0.008
R46632 S.n3469 S.n3468 0.008
R46633 S.n2816 S.n2815 0.008
R46634 S.n4610 S.n4609 0.008
R46635 S.n3943 S.n3942 0.008
R46636 S.n5745 S.n5744 0.008
R46637 S.n5055 S.n5054 0.008
R46638 S.n6855 S.n6854 0.008
R46639 S.n6155 S.n6154 0.008
R46640 S.n7953 S.n7952 0.008
R46641 S.n7232 S.n7231 0.008
R46642 S.n9028 S.n9027 0.008
R46643 S.n8296 S.n8295 0.008
R46644 S.n10091 S.n10090 0.008
R46645 S.n9338 S.n9337 0.008
R46646 S.n10367 S.n10366 0.008
R46647 S.n11372 S.n11371 0.008
R46648 S.n11798 S.n11794 0.008
R46649 S.n9037 S.n9036 0.008
R46650 S.n7962 S.n7961 0.008
R46651 S.n6864 S.n6863 0.008
R46652 S.n5754 S.n5753 0.008
R46653 S.n4619 S.n4618 0.008
R46654 S.n3478 S.n3477 0.008
R46655 S.n2323 S.n2322 0.008
R46656 S.n1006 S.n1003 0.008
R46657 S.n2372 S.n2371 0.008
R46658 S.n1608 S.n1607 0.008
R46659 S.n3529 S.n3528 0.008
R46660 S.n2780 S.n2779 0.008
R46661 S.n4671 S.n4670 0.008
R46662 S.n3907 S.n3906 0.008
R46663 S.n5806 S.n5805 0.008
R46664 S.n5019 S.n5018 0.008
R46665 S.n6916 S.n6915 0.008
R46666 S.n6119 S.n6118 0.008
R46667 S.n8014 S.n8013 0.008
R46668 S.n7196 S.n7195 0.008
R46669 S.n8260 S.n8259 0.008
R46670 S.n9300 S.n9299 0.008
R46671 S.n9730 S.n9728 0.008
R46672 S.n6925 S.n6924 0.008
R46673 S.n5815 S.n5814 0.008
R46674 S.n4680 S.n4679 0.008
R46675 S.n3538 S.n3537 0.008
R46676 S.n2382 S.n2381 0.008
R46677 S.n1036 S.n1035 0.008
R46678 S.n2431 S.n2430 0.008
R46679 S.n1571 S.n1570 0.008
R46680 S.n3589 S.n3588 0.008
R46681 S.n2744 S.n2743 0.008
R46682 S.n4732 S.n4731 0.008
R46683 S.n3871 S.n3870 0.008
R46684 S.n5867 S.n5866 0.008
R46685 S.n4983 S.n4982 0.008
R46686 S.n6083 S.n6082 0.008
R46687 S.n7158 S.n7157 0.008
R46688 S.n7592 S.n7590 0.008
R46689 S.n4741 S.n4740 0.008
R46690 S.n3598 S.n3597 0.008
R46691 S.n2441 S.n2440 0.008
R46692 S.n1070 S.n1067 0.008
R46693 S.n2490 S.n2489 0.008
R46694 S.n1534 S.n1533 0.008
R46695 S.n3649 S.n3648 0.008
R46696 S.n2708 S.n2707 0.008
R46697 S.n3835 S.n3834 0.008
R46698 S.n4945 S.n4944 0.008
R46699 S.n5383 S.n5381 0.008
R46700 S.n2500 S.n2499 0.008
R46701 S.n1102 S.n1099 0.008
R46702 S.n1497 S.n1496 0.008
R46703 S.n2670 S.n2669 0.008
R46704 S.n3113 S.n3111 0.008
R46705 S.n1132 S.n1131 0.008
R46706 S.n941 S.n940 0.008
R46707 S.n22753 S.n22752 0.008
R46708 S.t158 S.n1305 0.007
R46709 S.t158 S.n1298 0.007
R46710 S.t158 S.n1286 0.007
R46711 S.t158 S.n1274 0.007
R46712 S.t158 S.n1261 0.007
R46713 S.t158 S.n1248 0.007
R46714 S.t158 S.n1235 0.007
R46715 S.t158 S.n1222 0.007
R46716 S.t158 S.n1209 0.007
R46717 S.t158 S.n1196 0.007
R46718 S.n21625 S.n21624 0.007
R46719 S.n20802 S.n20801 0.007
R46720 S.n20326 S.n20325 0.007
R46721 S.n19454 S.n19453 0.007
R46722 S.n1351 S.n1350 0.007
R46723 S.n929 S.n928 0.007
R46724 S.t41 S.n22959 0.006
R46725 S.t41 S.n22954 0.006
R46726 S.t41 S.n22947 0.006
R46727 S.t41 S.n22940 0.006
R46728 S.t41 S.n22933 0.006
R46729 S.t41 S.n22926 0.006
R46730 S.t41 S.n22919 0.006
R46731 S.t41 S.n22912 0.006
R46732 S.t41 S.n22905 0.006
R46733 S.t41 S.n22898 0.006
R46734 S.t41 S.n22891 0.006
R46735 S.t41 S.n22884 0.006
R46736 S.t41 S.n22877 0.006
R46737 S.t41 S.n22870 0.006
R46738 S.t41 S.n22863 0.006
R46739 S.t41 S.n22856 0.006
R46740 S.t41 S.n22849 0.006
R46741 S.t41 S.n22842 0.006
R46742 S.n131 S.n130 0.006
R46743 S.n848 S.n846 0.006
R46744 S.n8 S.n7 0.006
R46745 S.n55 S.n54 0.006
R46746 S.n119 S.n118 0.006
R46747 S.n1006 S.n1005 0.006
R46748 S.n1070 S.n1069 0.006
R46749 S.n1102 S.n1101 0.006
R46750 S.n22754 S.n22753 0.006
R46751 S.n888 S.n887 0.006
R46752 S.n22992 S.n22991 0.006
R46753 S.n23007 S.n23006 0.006
R46754 S.n914 S.n892 0.006
R46755 S.n838 S.n825 0.006
R46756 S.n2068 S.n2067 0.005
R46757 S.n19473 S.n19472 0.005
R46758 S.n18583 S.n18582 0.005
R46759 S.n17683 S.n17682 0.005
R46760 S.n16760 S.n16759 0.005
R46761 S.n15825 S.n15824 0.005
R46762 S.n14867 S.n14866 0.005
R46763 S.n13897 S.n13896 0.005
R46764 S.n12904 S.n12903 0.005
R46765 S.n11899 S.n11898 0.005
R46766 S.n10871 S.n10870 0.005
R46767 S.n9831 S.n9830 0.005
R46768 S.n8768 S.n8767 0.005
R46769 S.n7693 S.n7692 0.005
R46770 S.n6595 S.n6594 0.005
R46771 S.n5485 S.n5484 0.005
R46772 S.n4350 S.n4349 0.005
R46773 S.n3214 S.n3213 0.005
R46774 S.n904 S.n903 0.005
R46775 S.t158 S.n1310 0.005
R46776 S.n19364 S.n19363 0.005
R46777 S.n17577 S.n17576 0.005
R46778 S.n15719 S.n15718 0.005
R46779 S.n13791 S.n13790 0.005
R46780 S.n11793 S.n11792 0.005
R46781 S.n9725 S.n9724 0.005
R46782 S.n7587 S.n7586 0.005
R46783 S.n5378 S.n5377 0.005
R46784 S.n3108 S.n3107 0.005
R46785 S.n22989 S.n22985 0.005
R46786 S.n23005 S.n23001 0.005
R46787 S.t158 S.n1353 0.005
R46788 S.n20181 S.n20180 0.004
R46789 S.n21129 S.n21128 0.004
R46790 S.n22635 S.n22634 0.004
R46791 S.n22006 S.n22005 0.004
R46792 S.n21612 S.n21611 0.004
R46793 S.n21938 S.n21937 0.004
R46794 S.n20789 S.n20788 0.004
R46795 S.n21146 S.n21145 0.004
R46796 S.n22654 S.n22653 0.004
R46797 S.n21993 S.n21992 0.004
R46798 S.n21636 S.n21635 0.004
R46799 S.n21959 S.n21958 0.004
R46800 S.n20813 S.n20812 0.004
R46801 S.n20341 S.n20340 0.004
R46802 S.n19311 S.n19310 0.004
R46803 S.n19529 S.n19528 0.004
R46804 S.n22619 S.n22618 0.004
R46805 S.n22021 S.n22020 0.004
R46806 S.n21596 S.n21595 0.004
R46807 S.n21923 S.n21922 0.004
R46808 S.n20773 S.n20772 0.004
R46809 S.n21113 S.n21112 0.004
R46810 S.n20162 S.n20161 0.004
R46811 S.n19501 S.n19500 0.004
R46812 S.n18429 S.n18428 0.004
R46813 S.n18672 S.n18671 0.004
R46814 S.n22603 S.n22602 0.004
R46815 S.n22036 S.n22035 0.004
R46816 S.n21580 S.n21579 0.004
R46817 S.n21908 S.n21907 0.004
R46818 S.n20757 S.n20756 0.004
R46819 S.n21098 S.n21097 0.004
R46820 S.n20146 S.n20145 0.004
R46821 S.n19544 S.n19543 0.004
R46822 S.n19292 S.n19291 0.004
R46823 S.n18644 S.n18643 0.004
R46824 S.n17524 S.n17523 0.004
R46825 S.n17804 S.n17803 0.004
R46826 S.n22587 S.n22586 0.004
R46827 S.n22051 S.n22050 0.004
R46828 S.n21564 S.n21563 0.004
R46829 S.n21893 S.n21892 0.004
R46830 S.n20741 S.n20740 0.004
R46831 S.n21083 S.n21082 0.004
R46832 S.n20130 S.n20129 0.004
R46833 S.n19559 S.n19558 0.004
R46834 S.n19276 S.n19275 0.004
R46835 S.n18687 S.n18686 0.004
R46836 S.n18410 S.n18409 0.004
R46837 S.n17776 S.n17775 0.004
R46838 S.n16606 S.n16605 0.004
R46839 S.n16910 S.n16909 0.004
R46840 S.n22571 S.n22570 0.004
R46841 S.n22066 S.n22065 0.004
R46842 S.n21548 S.n21547 0.004
R46843 S.n21878 S.n21877 0.004
R46844 S.n20725 S.n20724 0.004
R46845 S.n21068 S.n21067 0.004
R46846 S.n20114 S.n20113 0.004
R46847 S.n19574 S.n19573 0.004
R46848 S.n19260 S.n19259 0.004
R46849 S.n18702 S.n18701 0.004
R46850 S.n18394 S.n18393 0.004
R46851 S.n17819 S.n17818 0.004
R46852 S.n17505 S.n17504 0.004
R46853 S.n16882 S.n16881 0.004
R46854 S.n15666 S.n15665 0.004
R46855 S.n16007 S.n16006 0.004
R46856 S.n22555 S.n22554 0.004
R46857 S.n22081 S.n22080 0.004
R46858 S.n21532 S.n21531 0.004
R46859 S.n21863 S.n21862 0.004
R46860 S.n20709 S.n20708 0.004
R46861 S.n21053 S.n21052 0.004
R46862 S.n20098 S.n20097 0.004
R46863 S.n19589 S.n19588 0.004
R46864 S.n19244 S.n19243 0.004
R46865 S.n18717 S.n18716 0.004
R46866 S.n18378 S.n18377 0.004
R46867 S.n17834 S.n17833 0.004
R46868 S.n17489 S.n17488 0.004
R46869 S.n16925 S.n16924 0.004
R46870 S.n16587 S.n16586 0.004
R46871 S.n15979 S.n15978 0.004
R46872 S.n14713 S.n14712 0.004
R46873 S.n15078 S.n15077 0.004
R46874 S.n22539 S.n22538 0.004
R46875 S.n22096 S.n22095 0.004
R46876 S.n21516 S.n21515 0.004
R46877 S.n21848 S.n21847 0.004
R46878 S.n20693 S.n20692 0.004
R46879 S.n21038 S.n21037 0.004
R46880 S.n20082 S.n20081 0.004
R46881 S.n19604 S.n19603 0.004
R46882 S.n19228 S.n19227 0.004
R46883 S.n18732 S.n18731 0.004
R46884 S.n18362 S.n18361 0.004
R46885 S.n17849 S.n17848 0.004
R46886 S.n17473 S.n17472 0.004
R46887 S.n16940 S.n16939 0.004
R46888 S.n16571 S.n16570 0.004
R46889 S.n16022 S.n16021 0.004
R46890 S.n15647 S.n15646 0.004
R46891 S.n15050 S.n15049 0.004
R46892 S.n13738 S.n13737 0.004
R46893 S.n14140 S.n14139 0.004
R46894 S.n22523 S.n22522 0.004
R46895 S.n22111 S.n22110 0.004
R46896 S.n21500 S.n21499 0.004
R46897 S.n21833 S.n21832 0.004
R46898 S.n20677 S.n20676 0.004
R46899 S.n21023 S.n21022 0.004
R46900 S.n20066 S.n20065 0.004
R46901 S.n19619 S.n19618 0.004
R46902 S.n19212 S.n19211 0.004
R46903 S.n18747 S.n18746 0.004
R46904 S.n18346 S.n18345 0.004
R46905 S.n17864 S.n17863 0.004
R46906 S.n17457 S.n17456 0.004
R46907 S.n16955 S.n16954 0.004
R46908 S.n16555 S.n16554 0.004
R46909 S.n16037 S.n16036 0.004
R46910 S.n15631 S.n15630 0.004
R46911 S.n15093 S.n15092 0.004
R46912 S.n14694 S.n14693 0.004
R46913 S.n14112 S.n14111 0.004
R46914 S.n12750 S.n12749 0.004
R46915 S.n13176 S.n13175 0.004
R46916 S.n22507 S.n22506 0.004
R46917 S.n22126 S.n22125 0.004
R46918 S.n21484 S.n21483 0.004
R46919 S.n21818 S.n21817 0.004
R46920 S.n20661 S.n20660 0.004
R46921 S.n21008 S.n21007 0.004
R46922 S.n20050 S.n20049 0.004
R46923 S.n19634 S.n19633 0.004
R46924 S.n19196 S.n19195 0.004
R46925 S.n18762 S.n18761 0.004
R46926 S.n18330 S.n18329 0.004
R46927 S.n17879 S.n17878 0.004
R46928 S.n17441 S.n17440 0.004
R46929 S.n16970 S.n16969 0.004
R46930 S.n16539 S.n16538 0.004
R46931 S.n16052 S.n16051 0.004
R46932 S.n15615 S.n15614 0.004
R46933 S.n15108 S.n15107 0.004
R46934 S.n14678 S.n14677 0.004
R46935 S.n14155 S.n14154 0.004
R46936 S.n13719 S.n13718 0.004
R46937 S.n13148 S.n13147 0.004
R46938 S.n11740 S.n11739 0.004
R46939 S.n12203 S.n12202 0.004
R46940 S.n22491 S.n22490 0.004
R46941 S.n22141 S.n22140 0.004
R46942 S.n21468 S.n21467 0.004
R46943 S.n21803 S.n21802 0.004
R46944 S.n20645 S.n20644 0.004
R46945 S.n20993 S.n20992 0.004
R46946 S.n20034 S.n20033 0.004
R46947 S.n19649 S.n19648 0.004
R46948 S.n19180 S.n19179 0.004
R46949 S.n18777 S.n18776 0.004
R46950 S.n18314 S.n18313 0.004
R46951 S.n17894 S.n17893 0.004
R46952 S.n17425 S.n17424 0.004
R46953 S.n16985 S.n16984 0.004
R46954 S.n16523 S.n16522 0.004
R46955 S.n16067 S.n16066 0.004
R46956 S.n15599 S.n15598 0.004
R46957 S.n15123 S.n15122 0.004
R46958 S.n14662 S.n14661 0.004
R46959 S.n14170 S.n14169 0.004
R46960 S.n13703 S.n13702 0.004
R46961 S.n13191 S.n13190 0.004
R46962 S.n12731 S.n12730 0.004
R46963 S.n12175 S.n12174 0.004
R46964 S.n10717 S.n10716 0.004
R46965 S.n11204 S.n11203 0.004
R46966 S.n22475 S.n22474 0.004
R46967 S.n22156 S.n22155 0.004
R46968 S.n21452 S.n21451 0.004
R46969 S.n21788 S.n21787 0.004
R46970 S.n20629 S.n20628 0.004
R46971 S.n20978 S.n20977 0.004
R46972 S.n20018 S.n20017 0.004
R46973 S.n19664 S.n19663 0.004
R46974 S.n19164 S.n19163 0.004
R46975 S.n18792 S.n18791 0.004
R46976 S.n18298 S.n18297 0.004
R46977 S.n17909 S.n17908 0.004
R46978 S.n17409 S.n17408 0.004
R46979 S.n17000 S.n16999 0.004
R46980 S.n16507 S.n16506 0.004
R46981 S.n16082 S.n16081 0.004
R46982 S.n15583 S.n15582 0.004
R46983 S.n15138 S.n15137 0.004
R46984 S.n14646 S.n14645 0.004
R46985 S.n14185 S.n14184 0.004
R46986 S.n13687 S.n13686 0.004
R46987 S.n13206 S.n13205 0.004
R46988 S.n12715 S.n12714 0.004
R46989 S.n12218 S.n12217 0.004
R46990 S.n11721 S.n11720 0.004
R46991 S.n11176 S.n11175 0.004
R46992 S.n9672 S.n9671 0.004
R46993 S.n10196 S.n10195 0.004
R46994 S.n22459 S.n22458 0.004
R46995 S.n22171 S.n22170 0.004
R46996 S.n21436 S.n21435 0.004
R46997 S.n21773 S.n21772 0.004
R46998 S.n20613 S.n20612 0.004
R46999 S.n20963 S.n20962 0.004
R47000 S.n20002 S.n20001 0.004
R47001 S.n19679 S.n19678 0.004
R47002 S.n19148 S.n19147 0.004
R47003 S.n18807 S.n18806 0.004
R47004 S.n18282 S.n18281 0.004
R47005 S.n17924 S.n17923 0.004
R47006 S.n17393 S.n17392 0.004
R47007 S.n17015 S.n17014 0.004
R47008 S.n16491 S.n16490 0.004
R47009 S.n16097 S.n16096 0.004
R47010 S.n15567 S.n15566 0.004
R47011 S.n15153 S.n15152 0.004
R47012 S.n14630 S.n14629 0.004
R47013 S.n14200 S.n14199 0.004
R47014 S.n13671 S.n13670 0.004
R47015 S.n13221 S.n13220 0.004
R47016 S.n12699 S.n12698 0.004
R47017 S.n12233 S.n12232 0.004
R47018 S.n11705 S.n11704 0.004
R47019 S.n11219 S.n11218 0.004
R47020 S.n10698 S.n10697 0.004
R47021 S.n10168 S.n10167 0.004
R47022 S.n8614 S.n8613 0.004
R47023 S.n9162 S.n9161 0.004
R47024 S.n22443 S.n22442 0.004
R47025 S.n22186 S.n22185 0.004
R47026 S.n21420 S.n21419 0.004
R47027 S.n21758 S.n21757 0.004
R47028 S.n20597 S.n20596 0.004
R47029 S.n20948 S.n20947 0.004
R47030 S.n19986 S.n19985 0.004
R47031 S.n19694 S.n19693 0.004
R47032 S.n19132 S.n19131 0.004
R47033 S.n18822 S.n18821 0.004
R47034 S.n18266 S.n18265 0.004
R47035 S.n17939 S.n17938 0.004
R47036 S.n17377 S.n17376 0.004
R47037 S.n17030 S.n17029 0.004
R47038 S.n16475 S.n16474 0.004
R47039 S.n16112 S.n16111 0.004
R47040 S.n15551 S.n15550 0.004
R47041 S.n15168 S.n15167 0.004
R47042 S.n14614 S.n14613 0.004
R47043 S.n14215 S.n14214 0.004
R47044 S.n13655 S.n13654 0.004
R47045 S.n13236 S.n13235 0.004
R47046 S.n12683 S.n12682 0.004
R47047 S.n12248 S.n12247 0.004
R47048 S.n11689 S.n11688 0.004
R47049 S.n11234 S.n11233 0.004
R47050 S.n10682 S.n10681 0.004
R47051 S.n10211 S.n10210 0.004
R47052 S.n9653 S.n9652 0.004
R47053 S.n9134 S.n9133 0.004
R47054 S.n7534 S.n7533 0.004
R47055 S.n8119 S.n8118 0.004
R47056 S.n22427 S.n22426 0.004
R47057 S.n22201 S.n22200 0.004
R47058 S.n21404 S.n21403 0.004
R47059 S.n21743 S.n21742 0.004
R47060 S.n20581 S.n20580 0.004
R47061 S.n20933 S.n20932 0.004
R47062 S.n19970 S.n19969 0.004
R47063 S.n19709 S.n19708 0.004
R47064 S.n19116 S.n19115 0.004
R47065 S.n18837 S.n18836 0.004
R47066 S.n18250 S.n18249 0.004
R47067 S.n17954 S.n17953 0.004
R47068 S.n17361 S.n17360 0.004
R47069 S.n17045 S.n17044 0.004
R47070 S.n16459 S.n16458 0.004
R47071 S.n16127 S.n16126 0.004
R47072 S.n15535 S.n15534 0.004
R47073 S.n15183 S.n15182 0.004
R47074 S.n14598 S.n14597 0.004
R47075 S.n14230 S.n14229 0.004
R47076 S.n13639 S.n13638 0.004
R47077 S.n13251 S.n13250 0.004
R47078 S.n12667 S.n12666 0.004
R47079 S.n12263 S.n12262 0.004
R47080 S.n11673 S.n11672 0.004
R47081 S.n11249 S.n11248 0.004
R47082 S.n10666 S.n10665 0.004
R47083 S.n10226 S.n10225 0.004
R47084 S.n9637 S.n9636 0.004
R47085 S.n9177 S.n9176 0.004
R47086 S.n8595 S.n8594 0.004
R47087 S.n8091 S.n8090 0.004
R47088 S.n6441 S.n6440 0.004
R47089 S.n7050 S.n7049 0.004
R47090 S.n22411 S.n22410 0.004
R47091 S.n22216 S.n22215 0.004
R47092 S.n21388 S.n21387 0.004
R47093 S.n21728 S.n21727 0.004
R47094 S.n20565 S.n20564 0.004
R47095 S.n20918 S.n20917 0.004
R47096 S.n19954 S.n19953 0.004
R47097 S.n19724 S.n19723 0.004
R47098 S.n19100 S.n19099 0.004
R47099 S.n18852 S.n18851 0.004
R47100 S.n18234 S.n18233 0.004
R47101 S.n17969 S.n17968 0.004
R47102 S.n17345 S.n17344 0.004
R47103 S.n17060 S.n17059 0.004
R47104 S.n16443 S.n16442 0.004
R47105 S.n16142 S.n16141 0.004
R47106 S.n15519 S.n15518 0.004
R47107 S.n15198 S.n15197 0.004
R47108 S.n14582 S.n14581 0.004
R47109 S.n14245 S.n14244 0.004
R47110 S.n13623 S.n13622 0.004
R47111 S.n13266 S.n13265 0.004
R47112 S.n12651 S.n12650 0.004
R47113 S.n12278 S.n12277 0.004
R47114 S.n11657 S.n11656 0.004
R47115 S.n11264 S.n11263 0.004
R47116 S.n10650 S.n10649 0.004
R47117 S.n10241 S.n10240 0.004
R47118 S.n9621 S.n9620 0.004
R47119 S.n9192 S.n9191 0.004
R47120 S.n8579 S.n8578 0.004
R47121 S.n8134 S.n8133 0.004
R47122 S.n7515 S.n7514 0.004
R47123 S.n7022 S.n7021 0.004
R47124 S.n5325 S.n5324 0.004
R47125 S.n5972 S.n5971 0.004
R47126 S.n22395 S.n22394 0.004
R47127 S.n22231 S.n22230 0.004
R47128 S.n21372 S.n21371 0.004
R47129 S.n21713 S.n21712 0.004
R47130 S.n20549 S.n20548 0.004
R47131 S.n20903 S.n20902 0.004
R47132 S.n19938 S.n19937 0.004
R47133 S.n19739 S.n19738 0.004
R47134 S.n19084 S.n19083 0.004
R47135 S.n18867 S.n18866 0.004
R47136 S.n18218 S.n18217 0.004
R47137 S.n17984 S.n17983 0.004
R47138 S.n17329 S.n17328 0.004
R47139 S.n17075 S.n17074 0.004
R47140 S.n16427 S.n16426 0.004
R47141 S.n16157 S.n16156 0.004
R47142 S.n15503 S.n15502 0.004
R47143 S.n15213 S.n15212 0.004
R47144 S.n14566 S.n14565 0.004
R47145 S.n14260 S.n14259 0.004
R47146 S.n13607 S.n13606 0.004
R47147 S.n13281 S.n13280 0.004
R47148 S.n12635 S.n12634 0.004
R47149 S.n12293 S.n12292 0.004
R47150 S.n11641 S.n11640 0.004
R47151 S.n11279 S.n11278 0.004
R47152 S.n10634 S.n10633 0.004
R47153 S.n10256 S.n10255 0.004
R47154 S.n9605 S.n9604 0.004
R47155 S.n9207 S.n9206 0.004
R47156 S.n8563 S.n8562 0.004
R47157 S.n8149 S.n8148 0.004
R47158 S.n7499 S.n7498 0.004
R47159 S.n7065 S.n7064 0.004
R47160 S.n6422 S.n6421 0.004
R47161 S.n5944 S.n5943 0.004
R47162 S.n4196 S.n4195 0.004
R47163 S.n4867 S.n4866 0.004
R47164 S.n22379 S.n22378 0.004
R47165 S.n22246 S.n22245 0.004
R47166 S.n21356 S.n21355 0.004
R47167 S.n21698 S.n21697 0.004
R47168 S.n20533 S.n20532 0.004
R47169 S.n20888 S.n20887 0.004
R47170 S.n19922 S.n19921 0.004
R47171 S.n19754 S.n19753 0.004
R47172 S.n19068 S.n19067 0.004
R47173 S.n18882 S.n18881 0.004
R47174 S.n18202 S.n18201 0.004
R47175 S.n17999 S.n17998 0.004
R47176 S.n17313 S.n17312 0.004
R47177 S.n17090 S.n17089 0.004
R47178 S.n16411 S.n16410 0.004
R47179 S.n16172 S.n16171 0.004
R47180 S.n15487 S.n15486 0.004
R47181 S.n15228 S.n15227 0.004
R47182 S.n14550 S.n14549 0.004
R47183 S.n14275 S.n14274 0.004
R47184 S.n13591 S.n13590 0.004
R47185 S.n13296 S.n13295 0.004
R47186 S.n12619 S.n12618 0.004
R47187 S.n12308 S.n12307 0.004
R47188 S.n11625 S.n11624 0.004
R47189 S.n11294 S.n11293 0.004
R47190 S.n10618 S.n10617 0.004
R47191 S.n10271 S.n10270 0.004
R47192 S.n9589 S.n9588 0.004
R47193 S.n9225 S.n9224 0.004
R47194 S.n8547 S.n8546 0.004
R47195 S.n8164 S.n8163 0.004
R47196 S.n7483 S.n7482 0.004
R47197 S.n7080 S.n7079 0.004
R47198 S.n6406 S.n6405 0.004
R47199 S.n5987 S.n5986 0.004
R47200 S.n5306 S.n5305 0.004
R47201 S.n4838 S.n4837 0.004
R47202 S.n3055 S.n3054 0.004
R47203 S.n3754 S.n3753 0.004
R47204 S.n22269 S.n22268 0.004
R47205 S.n22261 S.n22260 0.004
R47206 S.n21675 S.n21674 0.004
R47207 S.n21667 S.n21666 0.004
R47208 S.n20518 S.n20517 0.004
R47209 S.n20872 S.n20871 0.004
R47210 S.n19907 S.n19906 0.004
R47211 S.n19769 S.n19768 0.004
R47212 S.n19053 S.n19052 0.004
R47213 S.n18897 S.n18896 0.004
R47214 S.n18187 S.n18186 0.004
R47215 S.n18014 S.n18013 0.004
R47216 S.n17298 S.n17297 0.004
R47217 S.n17105 S.n17104 0.004
R47218 S.n16396 S.n16395 0.004
R47219 S.n16187 S.n16186 0.004
R47220 S.n15472 S.n15471 0.004
R47221 S.n15243 S.n15242 0.004
R47222 S.n14535 S.n14534 0.004
R47223 S.n14290 S.n14289 0.004
R47224 S.n13576 S.n13575 0.004
R47225 S.n13311 S.n13310 0.004
R47226 S.n12604 S.n12603 0.004
R47227 S.n12323 S.n12322 0.004
R47228 S.n11610 S.n11609 0.004
R47229 S.n11309 S.n11308 0.004
R47230 S.n10603 S.n10602 0.004
R47231 S.n10286 S.n10285 0.004
R47232 S.n9574 S.n9573 0.004
R47233 S.n9237 S.n9236 0.004
R47234 S.n8532 S.n8531 0.004
R47235 S.n8179 S.n8178 0.004
R47236 S.n7468 S.n7467 0.004
R47237 S.n7095 S.n7094 0.004
R47238 S.n6391 S.n6390 0.004
R47239 S.n6002 S.n6001 0.004
R47240 S.n5291 S.n5290 0.004
R47241 S.n4882 S.n4881 0.004
R47242 S.n4178 S.n4177 0.004
R47243 S.n3725 S.n3724 0.004
R47244 S.n1897 S.n1896 0.004
R47245 S.n2623 S.n2622 0.004
R47246 S.n22362 S.n22361 0.004
R47247 S.n22686 S.n22685 0.004
R47248 S.n21280 S.n21279 0.004
R47249 S.n21272 S.n21271 0.004
R47250 S.n20503 S.n20502 0.004
R47251 S.n20856 S.n20855 0.004
R47252 S.n19892 S.n19891 0.004
R47253 S.n19785 S.n19784 0.004
R47254 S.n19038 S.n19037 0.004
R47255 S.n18913 S.n18912 0.004
R47256 S.n18172 S.n18171 0.004
R47257 S.n18030 S.n18029 0.004
R47258 S.n17283 S.n17282 0.004
R47259 S.n17121 S.n17120 0.004
R47260 S.n16381 S.n16380 0.004
R47261 S.n16203 S.n16202 0.004
R47262 S.n15457 S.n15456 0.004
R47263 S.n15259 S.n15258 0.004
R47264 S.n14520 S.n14519 0.004
R47265 S.n14306 S.n14305 0.004
R47266 S.n13561 S.n13560 0.004
R47267 S.n13327 S.n13326 0.004
R47268 S.n12589 S.n12588 0.004
R47269 S.n12339 S.n12338 0.004
R47270 S.n11595 S.n11594 0.004
R47271 S.n11325 S.n11324 0.004
R47272 S.n10588 S.n10587 0.004
R47273 S.n10302 S.n10301 0.004
R47274 S.n9559 S.n9558 0.004
R47275 S.n9253 S.n9252 0.004
R47276 S.n8517 S.n8516 0.004
R47277 S.n8195 S.n8194 0.004
R47278 S.n7453 S.n7452 0.004
R47279 S.n7111 S.n7110 0.004
R47280 S.n6376 S.n6375 0.004
R47281 S.n6018 S.n6017 0.004
R47282 S.n5276 S.n5275 0.004
R47283 S.n4898 S.n4897 0.004
R47284 S.n4163 S.n4162 0.004
R47285 S.n3770 S.n3769 0.004
R47286 S.n3037 S.n3036 0.004
R47287 S.n2594 S.n2593 0.004
R47288 S.n899 S.n898 0.004
R47289 S.n1975 S.n1974 0.004
R47290 S.n22726 S.n22725 0.004
R47291 S.n21306 S.n21305 0.004
R47292 S.n21205 S.n21204 0.004
R47293 S.n20483 S.n20482 0.004
R47294 S.n20386 S.n20385 0.004
R47295 S.n19872 S.n19871 0.004
R47296 S.n20259 S.n20258 0.004
R47297 S.n19018 S.n19017 0.004
R47298 S.n19391 S.n19390 0.004
R47299 S.n18152 S.n18151 0.004
R47300 S.n18504 S.n18503 0.004
R47301 S.n17263 S.n17262 0.004
R47302 S.n17604 S.n17603 0.004
R47303 S.n16361 S.n16360 0.004
R47304 S.n16681 S.n16680 0.004
R47305 S.n15437 S.n15436 0.004
R47306 S.n15746 S.n15745 0.004
R47307 S.n14500 S.n14499 0.004
R47308 S.n14788 S.n14787 0.004
R47309 S.n13541 S.n13540 0.004
R47310 S.n13818 S.n13817 0.004
R47311 S.n12569 S.n12568 0.004
R47312 S.n12825 S.n12824 0.004
R47313 S.n11575 S.n11574 0.004
R47314 S.n11820 S.n11819 0.004
R47315 S.n10568 S.n10567 0.004
R47316 S.n10792 S.n10791 0.004
R47317 S.n9539 S.n9538 0.004
R47318 S.n9752 S.n9751 0.004
R47319 S.n8497 S.n8496 0.004
R47320 S.n8689 S.n8688 0.004
R47321 S.n7433 S.n7432 0.004
R47322 S.n7614 S.n7613 0.004
R47323 S.n6356 S.n6355 0.004
R47324 S.n6516 S.n6515 0.004
R47325 S.n5256 S.n5255 0.004
R47326 S.n5405 S.n5404 0.004
R47327 S.n4143 S.n4142 0.004
R47328 S.n4271 S.n4270 0.004
R47329 S.n3017 S.n3016 0.004
R47330 S.n3135 S.n3134 0.004
R47331 S.n1856 S.n1855 0.004
R47332 S.n883 S.n882 0.004
R47333 S.n801 S.n800 0.004
R47334 S.n954 S.n953 0.004
R47335 S.n22349 S.n22348 0.004
R47336 S.n22711 S.n22710 0.004
R47337 S.n21343 S.n21342 0.004
R47338 S.n21259 S.n21258 0.004
R47339 S.n20833 S.n20832 0.004
R47340 S.n20843 S.n20842 0.004
R47341 S.n20198 S.n20197 0.004
R47342 S.n20208 S.n20207 0.004
R47343 S.n19328 S.n19327 0.004
R47344 S.n19338 S.n19337 0.004
R47345 S.n18446 S.n18445 0.004
R47346 S.n18456 S.n18455 0.004
R47347 S.n17541 S.n17540 0.004
R47348 S.n17551 S.n17550 0.004
R47349 S.n16623 S.n16622 0.004
R47350 S.n16633 S.n16632 0.004
R47351 S.n15683 S.n15682 0.004
R47352 S.n15693 S.n15692 0.004
R47353 S.n14730 S.n14729 0.004
R47354 S.n14740 S.n14739 0.004
R47355 S.n13755 S.n13754 0.004
R47356 S.n13765 S.n13764 0.004
R47357 S.n12767 S.n12766 0.004
R47358 S.n12777 S.n12776 0.004
R47359 S.n11757 S.n11756 0.004
R47360 S.n11767 S.n11766 0.004
R47361 S.n10734 S.n10733 0.004
R47362 S.n10744 S.n10743 0.004
R47363 S.n9689 S.n9688 0.004
R47364 S.n9699 S.n9698 0.004
R47365 S.n8631 S.n8630 0.004
R47366 S.n8641 S.n8640 0.004
R47367 S.n7551 S.n7550 0.004
R47368 S.n7561 S.n7560 0.004
R47369 S.n6458 S.n6457 0.004
R47370 S.n6468 S.n6467 0.004
R47371 S.n5342 S.n5341 0.004
R47372 S.n5352 S.n5351 0.004
R47373 S.n4213 S.n4212 0.004
R47374 S.n4223 S.n4222 0.004
R47375 S.n3072 S.n3071 0.004
R47376 S.n3082 S.n3081 0.004
R47377 S.n1880 S.n1879 0.004
R47378 S.n1925 S.n1924 0.004
R47379 S.n404 S.n403 0.004
R47380 S.n2127 S.n2126 0.004
R47381 S.n18469 S.n18468 0.004
R47382 S.n17161 S.n17160 0.004
R47383 S.n17753 S.n17752 0.004
R47384 S.n16261 S.n16260 0.004
R47385 S.n16826 S.n16825 0.004
R47386 S.n15337 S.n15336 0.004
R47387 S.n15891 S.n15890 0.004
R47388 S.n14400 S.n14399 0.004
R47389 S.n14933 S.n14932 0.004
R47390 S.n13441 S.n13440 0.004
R47391 S.n13963 S.n13962 0.004
R47392 S.n12469 S.n12468 0.004
R47393 S.n12970 S.n12969 0.004
R47394 S.n11475 S.n11474 0.004
R47395 S.n11965 S.n11964 0.004
R47396 S.n10468 S.n10467 0.004
R47397 S.n10937 S.n10936 0.004
R47398 S.n9439 S.n9438 0.004
R47399 S.n9897 S.n9896 0.004
R47400 S.n8397 S.n8396 0.004
R47401 S.n8834 S.n8833 0.004
R47402 S.n7333 S.n7332 0.004
R47403 S.n7759 S.n7758 0.004
R47404 S.n6256 S.n6255 0.004
R47405 S.n6661 S.n6660 0.004
R47406 S.n5156 S.n5155 0.004
R47407 S.n5551 S.n5550 0.004
R47408 S.n4044 S.n4043 0.004
R47409 S.n4416 S.n4415 0.004
R47410 S.n2917 S.n2916 0.004
R47411 S.n3279 S.n3278 0.004
R47412 S.n1748 S.n1747 0.004
R47413 S.n22 S.n21 0.004
R47414 S.n19361 S.n19360 0.004
R47415 S.n18075 S.n18074 0.004
R47416 S.n18622 S.n18621 0.004
R47417 S.n17186 S.n17185 0.004
R47418 S.n17722 S.n17721 0.004
R47419 S.n16284 S.n16283 0.004
R47420 S.n16795 S.n16794 0.004
R47421 S.n15360 S.n15359 0.004
R47422 S.n15860 S.n15859 0.004
R47423 S.n14423 S.n14422 0.004
R47424 S.n14902 S.n14901 0.004
R47425 S.n13464 S.n13463 0.004
R47426 S.n13932 S.n13931 0.004
R47427 S.n12492 S.n12491 0.004
R47428 S.n12939 S.n12938 0.004
R47429 S.n11498 S.n11497 0.004
R47430 S.n11934 S.n11933 0.004
R47431 S.n10491 S.n10490 0.004
R47432 S.n10906 S.n10905 0.004
R47433 S.n9462 S.n9461 0.004
R47434 S.n9866 S.n9865 0.004
R47435 S.n8420 S.n8419 0.004
R47436 S.n8803 S.n8802 0.004
R47437 S.n7356 S.n7355 0.004
R47438 S.n7728 S.n7727 0.004
R47439 S.n6279 S.n6278 0.004
R47440 S.n6630 S.n6629 0.004
R47441 S.n5179 S.n5178 0.004
R47442 S.n5520 S.n5519 0.004
R47443 S.n4067 S.n4066 0.004
R47444 S.n4385 S.n4384 0.004
R47445 S.n2940 S.n2939 0.004
R47446 S.n3248 S.n3247 0.004
R47447 S.n1772 S.n1771 0.004
R47448 S.n1794 S.n1793 0.004
R47449 S.n2064 S.n2063 0.004
R47450 S.n821 S.n820 0.004
R47451 S.n832 S.n831 0.004
R47452 S.n3219 S.n3218 0.004
R47453 S.n4355 S.n4354 0.004
R47454 S.n5490 S.n5489 0.004
R47455 S.n6600 S.n6599 0.004
R47456 S.n7698 S.n7697 0.004
R47457 S.n8773 S.n8772 0.004
R47458 S.n9836 S.n9835 0.004
R47459 S.n10876 S.n10875 0.004
R47460 S.n11904 S.n11903 0.004
R47461 S.n12909 S.n12908 0.004
R47462 S.n13902 S.n13901 0.004
R47463 S.n14872 S.n14871 0.004
R47464 S.n15830 S.n15829 0.004
R47465 S.n16765 S.n16764 0.004
R47466 S.n17688 S.n17687 0.004
R47467 S.n18588 S.n18587 0.004
R47468 S.n19478 S.n19477 0.004
R47469 S.n20224 S.n20223 0.004
R47470 S.n18953 S.n18952 0.004
R47471 S.n18088 S.n18087 0.004
R47472 S.n17199 S.n17198 0.004
R47473 S.n16297 S.n16296 0.004
R47474 S.n15373 S.n15372 0.004
R47475 S.n14436 S.n14435 0.004
R47476 S.n13477 S.n13476 0.004
R47477 S.n12505 S.n12504 0.004
R47478 S.n11511 S.n11510 0.004
R47479 S.n10504 S.n10503 0.004
R47480 S.n9475 S.n9474 0.004
R47481 S.n8433 S.n8432 0.004
R47482 S.n7369 S.n7368 0.004
R47483 S.n6292 S.n6291 0.004
R47484 S.n5192 S.n5191 0.004
R47485 S.n4080 S.n4079 0.004
R47486 S.n2953 S.n2952 0.004
R47487 S.n2036 S.n2035 0.004
R47488 S.n757 S.n756 0.004
R47489 S.n1334 S.n1333 0.004
R47490 S.n20416 S.n20415 0.004
R47491 S.n19833 S.n19832 0.004
R47492 S.n20312 S.n20311 0.004
R47493 S.n18981 S.n18980 0.004
R47494 S.n19440 S.n19439 0.004
R47495 S.n18116 S.n18115 0.004
R47496 S.n18553 S.n18552 0.004
R47497 S.n17227 S.n17226 0.004
R47498 S.n17653 S.n17652 0.004
R47499 S.n16325 S.n16324 0.004
R47500 S.n16730 S.n16729 0.004
R47501 S.n15401 S.n15400 0.004
R47502 S.n15795 S.n15794 0.004
R47503 S.n14464 S.n14463 0.004
R47504 S.n14837 S.n14836 0.004
R47505 S.n13505 S.n13504 0.004
R47506 S.n13867 S.n13866 0.004
R47507 S.n12533 S.n12532 0.004
R47508 S.n12874 S.n12873 0.004
R47509 S.n11539 S.n11538 0.004
R47510 S.n11869 S.n11868 0.004
R47511 S.n10532 S.n10531 0.004
R47512 S.n10841 S.n10840 0.004
R47513 S.n9503 S.n9502 0.004
R47514 S.n9801 S.n9800 0.004
R47515 S.n8461 S.n8460 0.004
R47516 S.n8738 S.n8737 0.004
R47517 S.n7397 S.n7396 0.004
R47518 S.n7663 S.n7662 0.004
R47519 S.n6320 S.n6319 0.004
R47520 S.n6565 S.n6564 0.004
R47521 S.n5220 S.n5219 0.004
R47522 S.n5455 S.n5454 0.004
R47523 S.n4108 S.n4107 0.004
R47524 S.n4320 S.n4319 0.004
R47525 S.n2981 S.n2980 0.004
R47526 S.n3183 S.n3182 0.004
R47527 S.n1818 S.n1817 0.004
R47528 S.n2003 S.n2002 0.004
R47529 S.n781 S.n780 0.004
R47530 S.n1839 S.n1838 0.004
R47531 S.n3164 S.n3163 0.004
R47532 S.n3001 S.n3000 0.004
R47533 S.n4301 S.n4300 0.004
R47534 S.n4128 S.n4127 0.004
R47535 S.n5435 S.n5434 0.004
R47536 S.n5240 S.n5239 0.004
R47537 S.n6546 S.n6545 0.004
R47538 S.n6340 S.n6339 0.004
R47539 S.n7644 S.n7643 0.004
R47540 S.n7417 S.n7416 0.004
R47541 S.n8719 S.n8718 0.004
R47542 S.n8481 S.n8480 0.004
R47543 S.n9782 S.n9781 0.004
R47544 S.n9523 S.n9522 0.004
R47545 S.n10822 S.n10821 0.004
R47546 S.n10552 S.n10551 0.004
R47547 S.n11850 S.n11849 0.004
R47548 S.n11559 S.n11558 0.004
R47549 S.n12855 S.n12854 0.004
R47550 S.n12553 S.n12552 0.004
R47551 S.n13848 S.n13847 0.004
R47552 S.n13525 S.n13524 0.004
R47553 S.n14818 S.n14817 0.004
R47554 S.n14484 S.n14483 0.004
R47555 S.n15776 S.n15775 0.004
R47556 S.n15421 S.n15420 0.004
R47557 S.n16711 S.n16710 0.004
R47558 S.n16345 S.n16344 0.004
R47559 S.n17634 S.n17633 0.004
R47560 S.n17247 S.n17246 0.004
R47561 S.n18534 S.n18533 0.004
R47562 S.n18136 S.n18135 0.004
R47563 S.n19421 S.n19420 0.004
R47564 S.n19002 S.n19001 0.004
R47565 S.n20293 S.n20292 0.004
R47566 S.n19856 S.n19855 0.004
R47567 S.n20364 S.n20363 0.004
R47568 S.n20467 S.n20466 0.004
R47569 S.n21240 S.n21239 0.004
R47570 S.n856 S.n855 0.004
R47571 S.n2097 S.n2096 0.004
R47572 S.n741 S.n740 0.004
R47573 S.n724 S.n723 0.004
R47574 S.n372 S.n371 0.004
R47575 S.n2186 S.n2185 0.004
R47576 S.n16646 S.n16645 0.004
R47577 S.n15299 S.n15298 0.004
R47578 S.n15956 S.n15955 0.004
R47579 S.n14364 S.n14363 0.004
R47580 S.n14994 S.n14993 0.004
R47581 S.n13405 S.n13404 0.004
R47582 S.n14024 S.n14023 0.004
R47583 S.n12433 S.n12432 0.004
R47584 S.n13031 S.n13030 0.004
R47585 S.n11439 S.n11438 0.004
R47586 S.n12026 S.n12025 0.004
R47587 S.n10432 S.n10431 0.004
R47588 S.n10998 S.n10997 0.004
R47589 S.n9403 S.n9402 0.004
R47590 S.n9958 S.n9957 0.004
R47591 S.n8361 S.n8360 0.004
R47592 S.n8895 S.n8894 0.004
R47593 S.n7297 S.n7296 0.004
R47594 S.n7820 S.n7819 0.004
R47595 S.n6220 S.n6219 0.004
R47596 S.n6722 S.n6721 0.004
R47597 S.n5120 S.n5119 0.004
R47598 S.n5612 S.n5611 0.004
R47599 S.n4008 S.n4007 0.004
R47600 S.n4477 S.n4476 0.004
R47601 S.n2881 S.n2880 0.004
R47602 S.n3339 S.n3338 0.004
R47603 S.n1711 S.n1710 0.004
R47604 S.n69 S.n68 0.004
R47605 S.n17574 S.n17573 0.004
R47606 S.n16248 S.n16247 0.004
R47607 S.n16860 S.n16859 0.004
R47608 S.n15324 S.n15323 0.004
R47609 S.n15925 S.n15924 0.004
R47610 S.n14387 S.n14386 0.004
R47611 S.n14963 S.n14962 0.004
R47612 S.n13428 S.n13427 0.004
R47613 S.n13993 S.n13992 0.004
R47614 S.n12456 S.n12455 0.004
R47615 S.n13000 S.n12999 0.004
R47616 S.n11462 S.n11461 0.004
R47617 S.n11995 S.n11994 0.004
R47618 S.n10455 S.n10454 0.004
R47619 S.n10967 S.n10966 0.004
R47620 S.n9426 S.n9425 0.004
R47621 S.n9927 S.n9926 0.004
R47622 S.n8384 S.n8383 0.004
R47623 S.n8864 S.n8863 0.004
R47624 S.n7320 S.n7319 0.004
R47625 S.n7789 S.n7788 0.004
R47626 S.n6243 S.n6242 0.004
R47627 S.n6691 S.n6690 0.004
R47628 S.n5143 S.n5142 0.004
R47629 S.n5581 S.n5580 0.004
R47630 S.n4031 S.n4030 0.004
R47631 S.n4446 S.n4445 0.004
R47632 S.n2904 S.n2903 0.004
R47633 S.n3308 S.n3307 0.004
R47634 S.n1735 S.n1734 0.004
R47635 S.n2155 S.n2154 0.004
R47636 S.n706 S.n705 0.004
R47637 S.n689 S.n688 0.004
R47638 S.n340 S.n339 0.004
R47639 S.n2245 S.n2244 0.004
R47640 S.n14753 S.n14752 0.004
R47641 S.n13367 S.n13366 0.004
R47642 S.n14089 S.n14088 0.004
R47643 S.n12397 S.n12396 0.004
R47644 S.n13092 S.n13091 0.004
R47645 S.n11403 S.n11402 0.004
R47646 S.n12087 S.n12086 0.004
R47647 S.n10396 S.n10395 0.004
R47648 S.n11059 S.n11058 0.004
R47649 S.n9367 S.n9366 0.004
R47650 S.n10019 S.n10018 0.004
R47651 S.n8325 S.n8324 0.004
R47652 S.n8956 S.n8955 0.004
R47653 S.n7261 S.n7260 0.004
R47654 S.n7881 S.n7880 0.004
R47655 S.n6184 S.n6183 0.004
R47656 S.n6783 S.n6782 0.004
R47657 S.n5084 S.n5083 0.004
R47658 S.n5673 S.n5672 0.004
R47659 S.n3972 S.n3971 0.004
R47660 S.n4538 S.n4537 0.004
R47661 S.n2845 S.n2844 0.004
R47662 S.n3399 S.n3398 0.004
R47663 S.n1674 S.n1673 0.004
R47664 S.n101 S.n100 0.004
R47665 S.n15716 S.n15715 0.004
R47666 S.n14351 S.n14350 0.004
R47667 S.n15028 S.n15027 0.004
R47668 S.n13392 S.n13391 0.004
R47669 S.n14058 S.n14057 0.004
R47670 S.n12420 S.n12419 0.004
R47671 S.n13061 S.n13060 0.004
R47672 S.n11426 S.n11425 0.004
R47673 S.n12056 S.n12055 0.004
R47674 S.n10419 S.n10418 0.004
R47675 S.n11028 S.n11027 0.004
R47676 S.n9390 S.n9389 0.004
R47677 S.n9988 S.n9987 0.004
R47678 S.n8348 S.n8347 0.004
R47679 S.n8925 S.n8924 0.004
R47680 S.n7284 S.n7283 0.004
R47681 S.n7850 S.n7849 0.004
R47682 S.n6207 S.n6206 0.004
R47683 S.n6752 S.n6751 0.004
R47684 S.n5107 S.n5106 0.004
R47685 S.n5642 S.n5641 0.004
R47686 S.n3995 S.n3994 0.004
R47687 S.n4507 S.n4506 0.004
R47688 S.n2868 S.n2867 0.004
R47689 S.n3368 S.n3367 0.004
R47690 S.n1698 S.n1697 0.004
R47691 S.n2214 S.n2213 0.004
R47692 S.n671 S.n670 0.004
R47693 S.n654 S.n653 0.004
R47694 S.n308 S.n307 0.004
R47695 S.n2304 S.n2303 0.004
R47696 S.n12790 S.n12789 0.004
R47697 S.n11365 S.n11364 0.004
R47698 S.n12152 S.n12151 0.004
R47699 S.n10360 S.n10359 0.004
R47700 S.n11120 S.n11119 0.004
R47701 S.n9331 S.n9330 0.004
R47702 S.n10080 S.n10079 0.004
R47703 S.n8289 S.n8288 0.004
R47704 S.n9017 S.n9016 0.004
R47705 S.n7225 S.n7224 0.004
R47706 S.n7942 S.n7941 0.004
R47707 S.n6148 S.n6147 0.004
R47708 S.n6844 S.n6843 0.004
R47709 S.n5048 S.n5047 0.004
R47710 S.n5734 S.n5733 0.004
R47711 S.n3936 S.n3935 0.004
R47712 S.n4599 S.n4598 0.004
R47713 S.n2809 S.n2808 0.004
R47714 S.n3459 S.n3458 0.004
R47715 S.n1637 S.n1636 0.004
R47716 S.n988 S.n987 0.004
R47717 S.n13788 S.n13787 0.004
R47718 S.n12384 S.n12383 0.004
R47719 S.n13126 S.n13125 0.004
R47720 S.n11390 S.n11389 0.004
R47721 S.n12121 S.n12120 0.004
R47722 S.n10383 S.n10382 0.004
R47723 S.n11089 S.n11088 0.004
R47724 S.n9354 S.n9353 0.004
R47725 S.n10049 S.n10048 0.004
R47726 S.n8312 S.n8311 0.004
R47727 S.n8986 S.n8985 0.004
R47728 S.n7248 S.n7247 0.004
R47729 S.n7911 S.n7910 0.004
R47730 S.n6171 S.n6170 0.004
R47731 S.n6813 S.n6812 0.004
R47732 S.n5071 S.n5070 0.004
R47733 S.n5703 S.n5702 0.004
R47734 S.n3959 S.n3958 0.004
R47735 S.n4568 S.n4567 0.004
R47736 S.n2832 S.n2831 0.004
R47737 S.n3428 S.n3427 0.004
R47738 S.n1661 S.n1660 0.004
R47739 S.n2273 S.n2272 0.004
R47740 S.n636 S.n635 0.004
R47741 S.n619 S.n618 0.004
R47742 S.n276 S.n275 0.004
R47743 S.n2363 S.n2362 0.004
R47744 S.n10757 S.n10756 0.004
R47745 S.n9293 S.n9292 0.004
R47746 S.n10145 S.n10144 0.004
R47747 S.n8253 S.n8252 0.004
R47748 S.n9078 S.n9077 0.004
R47749 S.n7189 S.n7188 0.004
R47750 S.n8003 S.n8002 0.004
R47751 S.n6112 S.n6111 0.004
R47752 S.n6905 S.n6904 0.004
R47753 S.n5012 S.n5011 0.004
R47754 S.n5795 S.n5794 0.004
R47755 S.n3900 S.n3899 0.004
R47756 S.n4660 S.n4659 0.004
R47757 S.n2773 S.n2772 0.004
R47758 S.n3519 S.n3518 0.004
R47759 S.n1600 S.n1599 0.004
R47760 S.n1020 S.n1019 0.004
R47761 S.n11790 S.n11789 0.004
R47762 S.n10347 S.n10346 0.004
R47763 S.n11154 S.n11153 0.004
R47764 S.n9318 S.n9317 0.004
R47765 S.n10114 S.n10113 0.004
R47766 S.n8276 S.n8275 0.004
R47767 S.n9047 S.n9046 0.004
R47768 S.n7212 S.n7211 0.004
R47769 S.n7972 S.n7971 0.004
R47770 S.n6135 S.n6134 0.004
R47771 S.n6874 S.n6873 0.004
R47772 S.n5035 S.n5034 0.004
R47773 S.n5764 S.n5763 0.004
R47774 S.n3923 S.n3922 0.004
R47775 S.n4629 S.n4628 0.004
R47776 S.n2796 S.n2795 0.004
R47777 S.n3488 S.n3487 0.004
R47778 S.n1624 S.n1623 0.004
R47779 S.n2332 S.n2331 0.004
R47780 S.n601 S.n600 0.004
R47781 S.n584 S.n583 0.004
R47782 S.n247 S.n246 0.004
R47783 S.n2422 S.n2421 0.004
R47784 S.n8654 S.n8653 0.004
R47785 S.n7151 S.n7150 0.004
R47786 S.n8068 S.n8067 0.004
R47787 S.n6076 S.n6075 0.004
R47788 S.n6966 S.n6965 0.004
R47789 S.n4976 S.n4975 0.004
R47790 S.n5856 S.n5855 0.004
R47791 S.n3864 S.n3863 0.004
R47792 S.n4721 S.n4720 0.004
R47793 S.n2737 S.n2736 0.004
R47794 S.n3579 S.n3578 0.004
R47795 S.n1563 S.n1562 0.004
R47796 S.n1052 S.n1051 0.004
R47797 S.n9722 S.n9721 0.004
R47798 S.n8240 S.n8239 0.004
R47799 S.n9112 S.n9111 0.004
R47800 S.n7176 S.n7175 0.004
R47801 S.n8037 S.n8036 0.004
R47802 S.n6099 S.n6098 0.004
R47803 S.n6935 S.n6934 0.004
R47804 S.n4999 S.n4998 0.004
R47805 S.n5825 S.n5824 0.004
R47806 S.n3887 S.n3886 0.004
R47807 S.n4690 S.n4689 0.004
R47808 S.n2760 S.n2759 0.004
R47809 S.n3548 S.n3547 0.004
R47810 S.n1587 S.n1586 0.004
R47811 S.n2391 S.n2390 0.004
R47812 S.n566 S.n565 0.004
R47813 S.n549 S.n548 0.004
R47814 S.n212 S.n211 0.004
R47815 S.n2481 S.n2480 0.004
R47816 S.n6481 S.n6480 0.004
R47817 S.n4938 S.n4937 0.004
R47818 S.n5921 S.n5920 0.004
R47819 S.n3828 S.n3827 0.004
R47820 S.n4782 S.n4781 0.004
R47821 S.n2701 S.n2700 0.004
R47822 S.n3639 S.n3638 0.004
R47823 S.n1526 S.n1525 0.004
R47824 S.n1084 S.n1083 0.004
R47825 S.n7584 S.n7583 0.004
R47826 S.n6063 S.n6062 0.004
R47827 S.n7000 S.n6999 0.004
R47828 S.n4963 S.n4962 0.004
R47829 S.n5890 S.n5889 0.004
R47830 S.n3851 S.n3850 0.004
R47831 S.n4751 S.n4750 0.004
R47832 S.n2724 S.n2723 0.004
R47833 S.n3608 S.n3607 0.004
R47834 S.n1550 S.n1549 0.004
R47835 S.n2450 S.n2449 0.004
R47836 S.n531 S.n530 0.004
R47837 S.n514 S.n513 0.004
R47838 S.n180 S.n179 0.004
R47839 S.n2540 S.n2539 0.004
R47840 S.n4236 S.n4235 0.004
R47841 S.n2663 S.n2662 0.004
R47842 S.n3703 S.n3702 0.004
R47843 S.n1489 S.n1488 0.004
R47844 S.n1116 S.n1115 0.004
R47845 S.n5375 S.n5374 0.004
R47846 S.n3815 S.n3814 0.004
R47847 S.n4816 S.n4815 0.004
R47848 S.n2688 S.n2687 0.004
R47849 S.n3672 S.n3671 0.004
R47850 S.n1513 S.n1512 0.004
R47851 S.n2509 S.n2508 0.004
R47852 S.n496 S.n495 0.004
R47853 S.n479 S.n478 0.004
R47854 S.n148 S.n147 0.004
R47855 S.n1942 S.n1941 0.004
R47856 S.n1154 S.n1153 0.004
R47857 S.n3105 S.n3104 0.004
R47858 S.n1476 S.n1475 0.004
R47859 S.n2572 S.n2571 0.004
R47860 S.n461 S.n460 0.004
R47861 S.n445 S.n444 0.004
R47862 S.n935 S.n934 0.004
R47863 S.n1429 S.n1428 0.004
R47864 S.n21975 S.n21974 0.004
R47865 S.n22763 S.n22762 0.004
R47866 S.n21326 S.n21325 0.004
R47867 S.n22303 S.n22302 0.004
R47868 S.n22331 S.n22330 0.004
R47869 S.n22316 S.n22315 0.004
R47870 S.t158 S.n1317 0.004
R47871 S.n24 S.n23 0.004
R47872 S.n406 S.n405 0.004
R47873 S.n71 S.n70 0.004
R47874 S.n374 S.n373 0.004
R47875 S.n103 S.n102 0.004
R47876 S.n342 S.n341 0.004
R47877 S.n990 S.n989 0.004
R47878 S.n310 S.n309 0.004
R47879 S.n1022 S.n1021 0.004
R47880 S.n278 S.n277 0.004
R47881 S.n1054 S.n1053 0.004
R47882 S.n249 S.n248 0.004
R47883 S.n1086 S.n1085 0.004
R47884 S.n214 S.n213 0.004
R47885 S.n1118 S.n1117 0.004
R47886 S.n182 S.n181 0.004
R47887 S.n1156 S.n1155 0.004
R47888 S.n150 S.n149 0.004
R47889 S.t158 S.n1365 0.004
R47890 S.n19814 S.n19813 0.004
R47891 S.n432 S.n431 0.004
R47892 S.n21151 S.n21150 0.004
R47893 S.n20320 S.n20319 0.004
R47894 S.n19448 S.n19447 0.004
R47895 S.n18559 S.n18558 0.004
R47896 S.n17659 S.n17658 0.004
R47897 S.n16736 S.n16735 0.004
R47898 S.n15801 S.n15800 0.004
R47899 S.n14843 S.n14842 0.004
R47900 S.n13873 S.n13872 0.004
R47901 S.n12880 S.n12879 0.004
R47902 S.n11875 S.n11874 0.004
R47903 S.n10847 S.n10846 0.004
R47904 S.n9807 S.n9806 0.004
R47905 S.n8744 S.n8743 0.004
R47906 S.n7669 S.n7668 0.004
R47907 S.n6571 S.n6570 0.004
R47908 S.n5461 S.n5460 0.004
R47909 S.n4326 S.n4325 0.004
R47910 S.n3189 S.n3188 0.004
R47911 S.n2021 S.n2020 0.004
R47912 S.n1344 S.n1343 0.004
R47913 S.n22288 S.n22287 0.004
R47914 S.n19814 S.n19812 0.004
R47915 S.n786 S.n774 0.004
R47916 S.n1845 S.n1844 0.004
R47917 S.n3006 S.n2994 0.004
R47918 S.n4132 S.n4121 0.004
R47919 S.n5245 S.n5233 0.004
R47920 S.n6345 S.n6333 0.004
R47921 S.n7422 S.n7410 0.004
R47922 S.n8486 S.n8474 0.004
R47923 S.n9528 S.n9516 0.004
R47924 S.n10557 S.n10545 0.004
R47925 S.n11564 S.n11552 0.004
R47926 S.n12558 S.n12546 0.004
R47927 S.n13530 S.n13518 0.004
R47928 S.n14489 S.n14477 0.004
R47929 S.n15426 S.n15414 0.004
R47930 S.n16350 S.n16338 0.004
R47931 S.n17252 S.n17240 0.004
R47932 S.n18141 S.n18129 0.004
R47933 S.n19007 S.n18995 0.004
R47934 S.n19861 S.n19849 0.004
R47935 S.n20472 S.n20460 0.004
R47936 S.n21296 S.n21294 0.004
R47937 S.n18943 S.n18942 0.004
R47938 S.n743 S.n734 0.004
R47939 S.n18059 S.n18057 0.004
R47940 S.n17151 S.n17150 0.004
R47941 S.n708 S.n699 0.004
R47942 S.n16232 S.n16230 0.004
R47943 S.n15289 S.n15288 0.004
R47944 S.n673 S.n664 0.004
R47945 S.n14335 S.n14333 0.004
R47946 S.n13357 S.n13356 0.004
R47947 S.n638 S.n629 0.004
R47948 S.n12368 S.n12366 0.004
R47949 S.n11355 S.n11354 0.004
R47950 S.n603 S.n594 0.004
R47951 S.n10331 S.n10329 0.004
R47952 S.n9283 S.n9282 0.004
R47953 S.n568 S.n559 0.004
R47954 S.n8224 S.n8222 0.004
R47955 S.n7141 S.n7140 0.004
R47956 S.n533 S.n524 0.004
R47957 S.n6047 S.n6045 0.004
R47958 S.n4928 S.n4927 0.004
R47959 S.n498 S.n489 0.004
R47960 S.n3799 S.n3797 0.004
R47961 S.n1460 S.n1458 0.004
R47962 S.n2653 S.n2652 0.004
R47963 S.n432 S.n430 0.004
R47964 S.n22765 S.n22756 0.004
R47965 S.n21172 S.n21171 0.004
R47966 S.n2066 S.n2065 0.004
R47967 S.n19471 S.n19470 0.004
R47968 S.n18581 S.n18580 0.004
R47969 S.n17681 S.n17680 0.004
R47970 S.n16758 S.n16757 0.004
R47971 S.n15823 S.n15822 0.004
R47972 S.n14865 S.n14864 0.004
R47973 S.n13895 S.n13894 0.004
R47974 S.n12902 S.n12901 0.004
R47975 S.n11897 S.n11896 0.004
R47976 S.n10869 S.n10868 0.004
R47977 S.n9829 S.n9828 0.004
R47978 S.n8766 S.n8765 0.004
R47979 S.n7691 S.n7690 0.004
R47980 S.n6593 S.n6592 0.004
R47981 S.n5483 S.n5482 0.004
R47982 S.n4348 S.n4347 0.004
R47983 S.n3212 S.n3211 0.004
R47984 S.n20451 S.n20437 0.004
R47985 S.n18567 S.n18565 0.004
R47986 S.n17667 S.n17665 0.004
R47987 S.n16744 S.n16742 0.004
R47988 S.n15809 S.n15807 0.004
R47989 S.n14851 S.n14849 0.004
R47990 S.n13881 S.n13879 0.004
R47991 S.n12888 S.n12886 0.004
R47992 S.n11883 S.n11881 0.004
R47993 S.n10855 S.n10853 0.004
R47994 S.n9815 S.n9813 0.004
R47995 S.n8752 S.n8750 0.004
R47996 S.n7677 S.n7675 0.004
R47997 S.n6579 S.n6577 0.004
R47998 S.n5469 S.n5467 0.004
R47999 S.n4334 S.n4332 0.004
R48000 S.n3197 S.n3195 0.004
R48001 S.n2029 S.n2027 0.004
R48002 S.n1799 S.n1798 0.004
R48003 S.n19370 S.n19369 0.004
R48004 S.n18943 S.n18930 0.004
R48005 S.n17583 S.n17582 0.004
R48006 S.n17151 S.n17138 0.004
R48007 S.n15725 S.n15724 0.004
R48008 S.n15289 S.n15276 0.004
R48009 S.n13797 S.n13796 0.004
R48010 S.n13357 S.n13344 0.004
R48011 S.n11799 S.n11798 0.004
R48012 S.n11355 S.n11342 0.004
R48013 S.n9731 S.n9730 0.004
R48014 S.n9283 S.n9270 0.004
R48015 S.n7593 S.n7592 0.004
R48016 S.n7141 S.n7128 0.004
R48017 S.n5384 S.n5383 0.004
R48018 S.n4928 S.n4915 0.004
R48019 S.n3114 S.n3113 0.004
R48020 S.n2653 S.n2640 0.004
R48021 S.n463 S.n455 0.004
R48022 S.t41 S.n22953 0.004
R48023 S.t41 S.n22961 0.004
R48024 S.t41 S.n22946 0.004
R48025 S.t41 S.n22939 0.004
R48026 S.t41 S.n22932 0.004
R48027 S.t41 S.n22925 0.004
R48028 S.t41 S.n22918 0.004
R48029 S.t41 S.n22911 0.004
R48030 S.t41 S.n22904 0.004
R48031 S.t41 S.n22897 0.004
R48032 S.t41 S.n22890 0.004
R48033 S.t41 S.n22883 0.004
R48034 S.t41 S.n22876 0.004
R48035 S.t41 S.n22869 0.004
R48036 S.t41 S.n22862 0.004
R48037 S.t41 S.n22855 0.004
R48038 S.t41 S.n22848 0.004
R48039 S.t41 S.n22841 0.004
R48040 S.t41 S.n22832 0.004
R48041 S.t41 S.n22823 0.004
R48042 S.n22336 S.n22335 0.004
R48043 S.t158 S.n1185 0.004
R48044 S.t9 S.n22291 0.004
R48045 S.t158 S.n1300 0.004
R48046 S.t79 S.n18062 0.004
R48047 S.t158 S.n1418 0.004
R48048 S.t150 S.n18946 0.004
R48049 S.t158 S.n1315 0.004
R48050 S.t209 S.n19817 0.004
R48051 S.t158 S.n1362 0.004
R48052 S.t64 S.n20454 0.004
R48053 S.t100 S.n21299 0.004
R48054 S.t158 S.n1379 0.004
R48055 S.t158 S.n1288 0.004
R48056 S.t167 S.n16235 0.004
R48057 S.t158 S.n1414 0.004
R48058 S.t218 S.n17154 0.004
R48059 S.t158 S.n1276 0.004
R48060 S.t0 S.n14338 0.004
R48061 S.t158 S.n1410 0.004
R48062 S.t60 S.n15292 0.004
R48063 S.t158 S.n1263 0.004
R48064 S.t357 S.n12371 0.004
R48065 S.t158 S.n1406 0.004
R48066 S.t73 S.n13360 0.004
R48067 S.t158 S.n1250 0.004
R48068 S.t31 S.n10334 0.004
R48069 S.t158 S.n1402 0.004
R48070 S.t54 S.n11358 0.004
R48071 S.t158 S.n1237 0.004
R48072 S.t19 S.n8227 0.004
R48073 S.t158 S.n1398 0.004
R48074 S.t366 S.n9286 0.004
R48075 S.t158 S.n1224 0.004
R48076 S.t83 S.n6050 0.004
R48077 S.t158 S.n1394 0.004
R48078 S.t47 S.n7144 0.004
R48079 S.t158 S.n1211 0.004
R48080 S.t176 S.n3802 0.004
R48081 S.t158 S.n1390 0.004
R48082 S.t214 S.n4931 0.004
R48083 S.t158 S.n1198 0.004
R48084 S.t75 S.n1463 0.004
R48085 S.t158 S.n1386 0.004
R48086 S.t14 S.n2656 0.004
R48087 S.t158 S.n1382 0.004
R48088 S.t137 S.n435 0.004
R48089 S.t41 S.n22957 0.004
R48090 S.t41 S.n22964 0.004
R48091 S.t41 S.n22950 0.004
R48092 S.t41 S.n22943 0.004
R48093 S.t41 S.n22936 0.004
R48094 S.t41 S.n22929 0.004
R48095 S.t41 S.n22922 0.004
R48096 S.t41 S.n22915 0.004
R48097 S.t41 S.n22908 0.004
R48098 S.t41 S.n22901 0.004
R48099 S.t41 S.n22894 0.004
R48100 S.t41 S.n22887 0.004
R48101 S.t41 S.n22880 0.004
R48102 S.t41 S.n22873 0.004
R48103 S.t41 S.n22866 0.004
R48104 S.t41 S.n22859 0.004
R48105 S.t41 S.n22852 0.004
R48106 S.t41 S.n22845 0.004
R48107 S.t41 S.n22838 0.004
R48108 S.t41 S.n22829 0.004
R48109 S.t41 S.n22820 0.004
R48110 S.t41 S.n22995 0.004
R48111 S.t41 S.n22812 0.004
R48112 S.n1432 S.n1427 0.004
R48113 S.t88 S.n22773 0.004
R48114 S.t41 S.n22815 0.004
R48115 S.t158 S.n46 0.004
R48116 S.t158 S.n77 0.004
R48117 S.t158 S.n109 0.004
R48118 S.t158 S.n996 0.004
R48119 S.t158 S.n1028 0.004
R48120 S.t158 S.n1060 0.004
R48121 S.t158 S.n1092 0.004
R48122 S.t158 S.n1124 0.004
R48123 S.t158 S.n1162 0.004
R48124 S.t158 S.n1174 0.004
R48125 S.n823 S.n822 0.004
R48126 S.n1432 S.n1426 0.004
R48127 S.t158 S.n1292 0.004
R48128 S.t158 S.n1280 0.004
R48129 S.t158 S.n1267 0.004
R48130 S.t158 S.n1254 0.004
R48131 S.t158 S.n1241 0.004
R48132 S.t158 S.n1228 0.004
R48133 S.t158 S.n1215 0.004
R48134 S.t158 S.n1202 0.004
R48135 S.t158 S.n1189 0.004
R48136 S.n21296 S.n21295 0.004
R48137 S.n18961 S.n18950 0.004
R48138 S.n18096 S.n18085 0.004
R48139 S.n17207 S.n17196 0.004
R48140 S.n16305 S.n16294 0.004
R48141 S.n15381 S.n15370 0.004
R48142 S.n14444 S.n14433 0.004
R48143 S.n13485 S.n13474 0.004
R48144 S.n12513 S.n12502 0.004
R48145 S.n11519 S.n11508 0.004
R48146 S.n10512 S.n10501 0.004
R48147 S.n9483 S.n9472 0.004
R48148 S.n8441 S.n8430 0.004
R48149 S.n7377 S.n7366 0.004
R48150 S.n6300 S.n6289 0.004
R48151 S.n5200 S.n5189 0.004
R48152 S.n4088 S.n4077 0.004
R48153 S.n2961 S.n2950 0.004
R48154 S.n1422 S.n1421 0.003
R48155 S.n22310 S.n22309 0.003
R48156 S.n20339 S.n20338 0.003
R48157 S.n20186 S.n20185 0.003
R48158 S.n21136 S.n21135 0.003
R48159 S.n22643 S.n22642 0.003
R48160 S.n22016 S.n22015 0.003
R48161 S.n21620 S.n21619 0.003
R48162 S.n21945 S.n21944 0.003
R48163 S.n20797 S.n20796 0.003
R48164 S.n21142 S.n21141 0.003
R48165 S.n22659 S.n22658 0.003
R48166 S.n22001 S.n22000 0.003
R48167 S.n21641 S.n21640 0.003
R48168 S.n21965 S.n21964 0.003
R48169 S.n20821 S.n20820 0.003
R48170 S.n19499 S.n19498 0.003
R48171 S.n19316 S.n19315 0.003
R48172 S.n19539 S.n19538 0.003
R48173 S.n22627 S.n22626 0.003
R48174 S.n22031 S.n22030 0.003
R48175 S.n21604 S.n21603 0.003
R48176 S.n21930 S.n21929 0.003
R48177 S.n20781 S.n20780 0.003
R48178 S.n21120 S.n21119 0.003
R48179 S.n20170 S.n20169 0.003
R48180 S.n18642 S.n18641 0.003
R48181 S.n18434 S.n18433 0.003
R48182 S.n18682 S.n18681 0.003
R48183 S.n22611 S.n22610 0.003
R48184 S.n22046 S.n22045 0.003
R48185 S.n21588 S.n21587 0.003
R48186 S.n21915 S.n21914 0.003
R48187 S.n20765 S.n20764 0.003
R48188 S.n21105 S.n21104 0.003
R48189 S.n20154 S.n20153 0.003
R48190 S.n19554 S.n19553 0.003
R48191 S.n19300 S.n19299 0.003
R48192 S.n17774 S.n17773 0.003
R48193 S.n17529 S.n17528 0.003
R48194 S.n17814 S.n17813 0.003
R48195 S.n22595 S.n22594 0.003
R48196 S.n22061 S.n22060 0.003
R48197 S.n21572 S.n21571 0.003
R48198 S.n21900 S.n21899 0.003
R48199 S.n20749 S.n20748 0.003
R48200 S.n21090 S.n21089 0.003
R48201 S.n20138 S.n20137 0.003
R48202 S.n19569 S.n19568 0.003
R48203 S.n19284 S.n19283 0.003
R48204 S.n18697 S.n18696 0.003
R48205 S.n18418 S.n18417 0.003
R48206 S.n16880 S.n16879 0.003
R48207 S.n16611 S.n16610 0.003
R48208 S.n16920 S.n16919 0.003
R48209 S.n22579 S.n22578 0.003
R48210 S.n22076 S.n22075 0.003
R48211 S.n21556 S.n21555 0.003
R48212 S.n21885 S.n21884 0.003
R48213 S.n20733 S.n20732 0.003
R48214 S.n21075 S.n21074 0.003
R48215 S.n20122 S.n20121 0.003
R48216 S.n19584 S.n19583 0.003
R48217 S.n19268 S.n19267 0.003
R48218 S.n18712 S.n18711 0.003
R48219 S.n18402 S.n18401 0.003
R48220 S.n17829 S.n17828 0.003
R48221 S.n17513 S.n17512 0.003
R48222 S.n15977 S.n15976 0.003
R48223 S.n15671 S.n15670 0.003
R48224 S.n16017 S.n16016 0.003
R48225 S.n22563 S.n22562 0.003
R48226 S.n22091 S.n22090 0.003
R48227 S.n21540 S.n21539 0.003
R48228 S.n21870 S.n21869 0.003
R48229 S.n20717 S.n20716 0.003
R48230 S.n21060 S.n21059 0.003
R48231 S.n20106 S.n20105 0.003
R48232 S.n19599 S.n19598 0.003
R48233 S.n19252 S.n19251 0.003
R48234 S.n18727 S.n18726 0.003
R48235 S.n18386 S.n18385 0.003
R48236 S.n17844 S.n17843 0.003
R48237 S.n17497 S.n17496 0.003
R48238 S.n16935 S.n16934 0.003
R48239 S.n16595 S.n16594 0.003
R48240 S.n15048 S.n15047 0.003
R48241 S.n14718 S.n14717 0.003
R48242 S.n15088 S.n15087 0.003
R48243 S.n22547 S.n22546 0.003
R48244 S.n22106 S.n22105 0.003
R48245 S.n21524 S.n21523 0.003
R48246 S.n21855 S.n21854 0.003
R48247 S.n20701 S.n20700 0.003
R48248 S.n21045 S.n21044 0.003
R48249 S.n20090 S.n20089 0.003
R48250 S.n19614 S.n19613 0.003
R48251 S.n19236 S.n19235 0.003
R48252 S.n18742 S.n18741 0.003
R48253 S.n18370 S.n18369 0.003
R48254 S.n17859 S.n17858 0.003
R48255 S.n17481 S.n17480 0.003
R48256 S.n16950 S.n16949 0.003
R48257 S.n16579 S.n16578 0.003
R48258 S.n16032 S.n16031 0.003
R48259 S.n15655 S.n15654 0.003
R48260 S.n14110 S.n14109 0.003
R48261 S.n13743 S.n13742 0.003
R48262 S.n14150 S.n14149 0.003
R48263 S.n22531 S.n22530 0.003
R48264 S.n22121 S.n22120 0.003
R48265 S.n21508 S.n21507 0.003
R48266 S.n21840 S.n21839 0.003
R48267 S.n20685 S.n20684 0.003
R48268 S.n21030 S.n21029 0.003
R48269 S.n20074 S.n20073 0.003
R48270 S.n19629 S.n19628 0.003
R48271 S.n19220 S.n19219 0.003
R48272 S.n18757 S.n18756 0.003
R48273 S.n18354 S.n18353 0.003
R48274 S.n17874 S.n17873 0.003
R48275 S.n17465 S.n17464 0.003
R48276 S.n16965 S.n16964 0.003
R48277 S.n16563 S.n16562 0.003
R48278 S.n16047 S.n16046 0.003
R48279 S.n15639 S.n15638 0.003
R48280 S.n15103 S.n15102 0.003
R48281 S.n14702 S.n14701 0.003
R48282 S.n13146 S.n13145 0.003
R48283 S.n12755 S.n12754 0.003
R48284 S.n13186 S.n13185 0.003
R48285 S.n22515 S.n22514 0.003
R48286 S.n22136 S.n22135 0.003
R48287 S.n21492 S.n21491 0.003
R48288 S.n21825 S.n21824 0.003
R48289 S.n20669 S.n20668 0.003
R48290 S.n21015 S.n21014 0.003
R48291 S.n20058 S.n20057 0.003
R48292 S.n19644 S.n19643 0.003
R48293 S.n19204 S.n19203 0.003
R48294 S.n18772 S.n18771 0.003
R48295 S.n18338 S.n18337 0.003
R48296 S.n17889 S.n17888 0.003
R48297 S.n17449 S.n17448 0.003
R48298 S.n16980 S.n16979 0.003
R48299 S.n16547 S.n16546 0.003
R48300 S.n16062 S.n16061 0.003
R48301 S.n15623 S.n15622 0.003
R48302 S.n15118 S.n15117 0.003
R48303 S.n14686 S.n14685 0.003
R48304 S.n14165 S.n14164 0.003
R48305 S.n13727 S.n13726 0.003
R48306 S.n12173 S.n12172 0.003
R48307 S.n11745 S.n11744 0.003
R48308 S.n12213 S.n12212 0.003
R48309 S.n22499 S.n22498 0.003
R48310 S.n22151 S.n22150 0.003
R48311 S.n21476 S.n21475 0.003
R48312 S.n21810 S.n21809 0.003
R48313 S.n20653 S.n20652 0.003
R48314 S.n21000 S.n20999 0.003
R48315 S.n20042 S.n20041 0.003
R48316 S.n19659 S.n19658 0.003
R48317 S.n19188 S.n19187 0.003
R48318 S.n18787 S.n18786 0.003
R48319 S.n18322 S.n18321 0.003
R48320 S.n17904 S.n17903 0.003
R48321 S.n17433 S.n17432 0.003
R48322 S.n16995 S.n16994 0.003
R48323 S.n16531 S.n16530 0.003
R48324 S.n16077 S.n16076 0.003
R48325 S.n15607 S.n15606 0.003
R48326 S.n15133 S.n15132 0.003
R48327 S.n14670 S.n14669 0.003
R48328 S.n14180 S.n14179 0.003
R48329 S.n13711 S.n13710 0.003
R48330 S.n13201 S.n13200 0.003
R48331 S.n12739 S.n12738 0.003
R48332 S.n11174 S.n11173 0.003
R48333 S.n10722 S.n10721 0.003
R48334 S.n11214 S.n11213 0.003
R48335 S.n22483 S.n22482 0.003
R48336 S.n22166 S.n22165 0.003
R48337 S.n21460 S.n21459 0.003
R48338 S.n21795 S.n21794 0.003
R48339 S.n20637 S.n20636 0.003
R48340 S.n20985 S.n20984 0.003
R48341 S.n20026 S.n20025 0.003
R48342 S.n19674 S.n19673 0.003
R48343 S.n19172 S.n19171 0.003
R48344 S.n18802 S.n18801 0.003
R48345 S.n18306 S.n18305 0.003
R48346 S.n17919 S.n17918 0.003
R48347 S.n17417 S.n17416 0.003
R48348 S.n17010 S.n17009 0.003
R48349 S.n16515 S.n16514 0.003
R48350 S.n16092 S.n16091 0.003
R48351 S.n15591 S.n15590 0.003
R48352 S.n15148 S.n15147 0.003
R48353 S.n14654 S.n14653 0.003
R48354 S.n14195 S.n14194 0.003
R48355 S.n13695 S.n13694 0.003
R48356 S.n13216 S.n13215 0.003
R48357 S.n12723 S.n12722 0.003
R48358 S.n12228 S.n12227 0.003
R48359 S.n11729 S.n11728 0.003
R48360 S.n10166 S.n10165 0.003
R48361 S.n9677 S.n9676 0.003
R48362 S.n10206 S.n10205 0.003
R48363 S.n22467 S.n22466 0.003
R48364 S.n22181 S.n22180 0.003
R48365 S.n21444 S.n21443 0.003
R48366 S.n21780 S.n21779 0.003
R48367 S.n20621 S.n20620 0.003
R48368 S.n20970 S.n20969 0.003
R48369 S.n20010 S.n20009 0.003
R48370 S.n19689 S.n19688 0.003
R48371 S.n19156 S.n19155 0.003
R48372 S.n18817 S.n18816 0.003
R48373 S.n18290 S.n18289 0.003
R48374 S.n17934 S.n17933 0.003
R48375 S.n17401 S.n17400 0.003
R48376 S.n17025 S.n17024 0.003
R48377 S.n16499 S.n16498 0.003
R48378 S.n16107 S.n16106 0.003
R48379 S.n15575 S.n15574 0.003
R48380 S.n15163 S.n15162 0.003
R48381 S.n14638 S.n14637 0.003
R48382 S.n14210 S.n14209 0.003
R48383 S.n13679 S.n13678 0.003
R48384 S.n13231 S.n13230 0.003
R48385 S.n12707 S.n12706 0.003
R48386 S.n12243 S.n12242 0.003
R48387 S.n11713 S.n11712 0.003
R48388 S.n11229 S.n11228 0.003
R48389 S.n10706 S.n10705 0.003
R48390 S.n9132 S.n9131 0.003
R48391 S.n8619 S.n8618 0.003
R48392 S.n9172 S.n9171 0.003
R48393 S.n22451 S.n22450 0.003
R48394 S.n22196 S.n22195 0.003
R48395 S.n21428 S.n21427 0.003
R48396 S.n21765 S.n21764 0.003
R48397 S.n20605 S.n20604 0.003
R48398 S.n20955 S.n20954 0.003
R48399 S.n19994 S.n19993 0.003
R48400 S.n19704 S.n19703 0.003
R48401 S.n19140 S.n19139 0.003
R48402 S.n18832 S.n18831 0.003
R48403 S.n18274 S.n18273 0.003
R48404 S.n17949 S.n17948 0.003
R48405 S.n17385 S.n17384 0.003
R48406 S.n17040 S.n17039 0.003
R48407 S.n16483 S.n16482 0.003
R48408 S.n16122 S.n16121 0.003
R48409 S.n15559 S.n15558 0.003
R48410 S.n15178 S.n15177 0.003
R48411 S.n14622 S.n14621 0.003
R48412 S.n14225 S.n14224 0.003
R48413 S.n13663 S.n13662 0.003
R48414 S.n13246 S.n13245 0.003
R48415 S.n12691 S.n12690 0.003
R48416 S.n12258 S.n12257 0.003
R48417 S.n11697 S.n11696 0.003
R48418 S.n11244 S.n11243 0.003
R48419 S.n10690 S.n10689 0.003
R48420 S.n10221 S.n10220 0.003
R48421 S.n9661 S.n9660 0.003
R48422 S.n8089 S.n8088 0.003
R48423 S.n7539 S.n7538 0.003
R48424 S.n8129 S.n8128 0.003
R48425 S.n22435 S.n22434 0.003
R48426 S.n22211 S.n22210 0.003
R48427 S.n21412 S.n21411 0.003
R48428 S.n21750 S.n21749 0.003
R48429 S.n20589 S.n20588 0.003
R48430 S.n20940 S.n20939 0.003
R48431 S.n19978 S.n19977 0.003
R48432 S.n19719 S.n19718 0.003
R48433 S.n19124 S.n19123 0.003
R48434 S.n18847 S.n18846 0.003
R48435 S.n18258 S.n18257 0.003
R48436 S.n17964 S.n17963 0.003
R48437 S.n17369 S.n17368 0.003
R48438 S.n17055 S.n17054 0.003
R48439 S.n16467 S.n16466 0.003
R48440 S.n16137 S.n16136 0.003
R48441 S.n15543 S.n15542 0.003
R48442 S.n15193 S.n15192 0.003
R48443 S.n14606 S.n14605 0.003
R48444 S.n14240 S.n14239 0.003
R48445 S.n13647 S.n13646 0.003
R48446 S.n13261 S.n13260 0.003
R48447 S.n12675 S.n12674 0.003
R48448 S.n12273 S.n12272 0.003
R48449 S.n11681 S.n11680 0.003
R48450 S.n11259 S.n11258 0.003
R48451 S.n10674 S.n10673 0.003
R48452 S.n10236 S.n10235 0.003
R48453 S.n9645 S.n9644 0.003
R48454 S.n9187 S.n9186 0.003
R48455 S.n8603 S.n8602 0.003
R48456 S.n7020 S.n7019 0.003
R48457 S.n6446 S.n6445 0.003
R48458 S.n7060 S.n7059 0.003
R48459 S.n22419 S.n22418 0.003
R48460 S.n22226 S.n22225 0.003
R48461 S.n21396 S.n21395 0.003
R48462 S.n21735 S.n21734 0.003
R48463 S.n20573 S.n20572 0.003
R48464 S.n20925 S.n20924 0.003
R48465 S.n19962 S.n19961 0.003
R48466 S.n19734 S.n19733 0.003
R48467 S.n19108 S.n19107 0.003
R48468 S.n18862 S.n18861 0.003
R48469 S.n18242 S.n18241 0.003
R48470 S.n17979 S.n17978 0.003
R48471 S.n17353 S.n17352 0.003
R48472 S.n17070 S.n17069 0.003
R48473 S.n16451 S.n16450 0.003
R48474 S.n16152 S.n16151 0.003
R48475 S.n15527 S.n15526 0.003
R48476 S.n15208 S.n15207 0.003
R48477 S.n14590 S.n14589 0.003
R48478 S.n14255 S.n14254 0.003
R48479 S.n13631 S.n13630 0.003
R48480 S.n13276 S.n13275 0.003
R48481 S.n12659 S.n12658 0.003
R48482 S.n12288 S.n12287 0.003
R48483 S.n11665 S.n11664 0.003
R48484 S.n11274 S.n11273 0.003
R48485 S.n10658 S.n10657 0.003
R48486 S.n10251 S.n10250 0.003
R48487 S.n9629 S.n9628 0.003
R48488 S.n9202 S.n9201 0.003
R48489 S.n8587 S.n8586 0.003
R48490 S.n8144 S.n8143 0.003
R48491 S.n7523 S.n7522 0.003
R48492 S.n5942 S.n5941 0.003
R48493 S.n5330 S.n5329 0.003
R48494 S.n5982 S.n5981 0.003
R48495 S.n22403 S.n22402 0.003
R48496 S.n22241 S.n22240 0.003
R48497 S.n21380 S.n21379 0.003
R48498 S.n21720 S.n21719 0.003
R48499 S.n20557 S.n20556 0.003
R48500 S.n20910 S.n20909 0.003
R48501 S.n19946 S.n19945 0.003
R48502 S.n19749 S.n19748 0.003
R48503 S.n19092 S.n19091 0.003
R48504 S.n18877 S.n18876 0.003
R48505 S.n18226 S.n18225 0.003
R48506 S.n17994 S.n17993 0.003
R48507 S.n17337 S.n17336 0.003
R48508 S.n17085 S.n17084 0.003
R48509 S.n16435 S.n16434 0.003
R48510 S.n16167 S.n16166 0.003
R48511 S.n15511 S.n15510 0.003
R48512 S.n15223 S.n15222 0.003
R48513 S.n14574 S.n14573 0.003
R48514 S.n14270 S.n14269 0.003
R48515 S.n13615 S.n13614 0.003
R48516 S.n13291 S.n13290 0.003
R48517 S.n12643 S.n12642 0.003
R48518 S.n12303 S.n12302 0.003
R48519 S.n11649 S.n11648 0.003
R48520 S.n11289 S.n11288 0.003
R48521 S.n10642 S.n10641 0.003
R48522 S.n10266 S.n10265 0.003
R48523 S.n9613 S.n9612 0.003
R48524 S.n9217 S.n9216 0.003
R48525 S.n8571 S.n8570 0.003
R48526 S.n8159 S.n8158 0.003
R48527 S.n7507 S.n7506 0.003
R48528 S.n7075 S.n7074 0.003
R48529 S.n6430 S.n6429 0.003
R48530 S.n4836 S.n4835 0.003
R48531 S.n4201 S.n4200 0.003
R48532 S.n4877 S.n4876 0.003
R48533 S.n22387 S.n22386 0.003
R48534 S.n22256 S.n22255 0.003
R48535 S.n21364 S.n21363 0.003
R48536 S.n21705 S.n21704 0.003
R48537 S.n20541 S.n20540 0.003
R48538 S.n20895 S.n20894 0.003
R48539 S.n19930 S.n19929 0.003
R48540 S.n19764 S.n19763 0.003
R48541 S.n19076 S.n19075 0.003
R48542 S.n18892 S.n18891 0.003
R48543 S.n18210 S.n18209 0.003
R48544 S.n18009 S.n18008 0.003
R48545 S.n17321 S.n17320 0.003
R48546 S.n17100 S.n17099 0.003
R48547 S.n16419 S.n16418 0.003
R48548 S.n16182 S.n16181 0.003
R48549 S.n15495 S.n15494 0.003
R48550 S.n15238 S.n15237 0.003
R48551 S.n14558 S.n14557 0.003
R48552 S.n14285 S.n14284 0.003
R48553 S.n13599 S.n13598 0.003
R48554 S.n13306 S.n13305 0.003
R48555 S.n12627 S.n12626 0.003
R48556 S.n12318 S.n12317 0.003
R48557 S.n11633 S.n11632 0.003
R48558 S.n11304 S.n11303 0.003
R48559 S.n10626 S.n10625 0.003
R48560 S.n10281 S.n10280 0.003
R48561 S.n9597 S.n9596 0.003
R48562 S.n9232 S.n9231 0.003
R48563 S.n8555 S.n8554 0.003
R48564 S.n8174 S.n8173 0.003
R48565 S.n7491 S.n7490 0.003
R48566 S.n7090 S.n7089 0.003
R48567 S.n6414 S.n6413 0.003
R48568 S.n5997 S.n5996 0.003
R48569 S.n5314 S.n5313 0.003
R48570 S.n3723 S.n3722 0.003
R48571 S.n3060 S.n3059 0.003
R48572 S.n3765 S.n3764 0.003
R48573 S.n22668 S.n22667 0.003
R48574 S.n22681 S.n22680 0.003
R48575 S.n21681 S.n21680 0.003
R48576 S.n21690 S.n21689 0.003
R48577 S.n20525 S.n20524 0.003
R48578 S.n20880 S.n20879 0.003
R48579 S.n19914 S.n19913 0.003
R48580 S.n19780 S.n19779 0.003
R48581 S.n19060 S.n19059 0.003
R48582 S.n18908 S.n18907 0.003
R48583 S.n18194 S.n18193 0.003
R48584 S.n18025 S.n18024 0.003
R48585 S.n17305 S.n17304 0.003
R48586 S.n17116 S.n17115 0.003
R48587 S.n16403 S.n16402 0.003
R48588 S.n16198 S.n16197 0.003
R48589 S.n15479 S.n15478 0.003
R48590 S.n15254 S.n15253 0.003
R48591 S.n14542 S.n14541 0.003
R48592 S.n14301 S.n14300 0.003
R48593 S.n13583 S.n13582 0.003
R48594 S.n13322 S.n13321 0.003
R48595 S.n12611 S.n12610 0.003
R48596 S.n12334 S.n12333 0.003
R48597 S.n11617 S.n11616 0.003
R48598 S.n11320 S.n11319 0.003
R48599 S.n10610 S.n10609 0.003
R48600 S.n10297 S.n10296 0.003
R48601 S.n9581 S.n9580 0.003
R48602 S.n9248 S.n9247 0.003
R48603 S.n8539 S.n8538 0.003
R48604 S.n8190 S.n8189 0.003
R48605 S.n7475 S.n7474 0.003
R48606 S.n7106 S.n7105 0.003
R48607 S.n6398 S.n6397 0.003
R48608 S.n6013 S.n6012 0.003
R48609 S.n5298 S.n5297 0.003
R48610 S.n4893 S.n4892 0.003
R48611 S.n4185 S.n4184 0.003
R48612 S.n2592 S.n2591 0.003
R48613 S.n1891 S.n1890 0.003
R48614 S.n2634 S.n2633 0.003
R48615 S.n22371 S.n22370 0.003
R48616 S.n22700 S.n22699 0.003
R48617 S.n21650 S.n21649 0.003
R48618 S.n21659 S.n21658 0.003
R48619 S.n20510 S.n20509 0.003
R48620 S.n20864 S.n20863 0.003
R48621 S.n19899 S.n19898 0.003
R48622 S.n19796 S.n19795 0.003
R48623 S.n19045 S.n19044 0.003
R48624 S.n18924 S.n18923 0.003
R48625 S.n18179 S.n18178 0.003
R48626 S.n18041 S.n18040 0.003
R48627 S.n17290 S.n17289 0.003
R48628 S.n17132 S.n17131 0.003
R48629 S.n16388 S.n16387 0.003
R48630 S.n16214 S.n16213 0.003
R48631 S.n15464 S.n15463 0.003
R48632 S.n15270 S.n15269 0.003
R48633 S.n14527 S.n14526 0.003
R48634 S.n14317 S.n14316 0.003
R48635 S.n13568 S.n13567 0.003
R48636 S.n13338 S.n13337 0.003
R48637 S.n12596 S.n12595 0.003
R48638 S.n12350 S.n12349 0.003
R48639 S.n11602 S.n11601 0.003
R48640 S.n11336 S.n11335 0.003
R48641 S.n10595 S.n10594 0.003
R48642 S.n10313 S.n10312 0.003
R48643 S.n9566 S.n9565 0.003
R48644 S.n9264 S.n9263 0.003
R48645 S.n8524 S.n8523 0.003
R48646 S.n8206 S.n8205 0.003
R48647 S.n7460 S.n7459 0.003
R48648 S.n7122 S.n7121 0.003
R48649 S.n6383 S.n6382 0.003
R48650 S.n6029 S.n6028 0.003
R48651 S.n5283 S.n5282 0.003
R48652 S.n4909 S.n4908 0.003
R48653 S.n4170 S.n4169 0.003
R48654 S.n3781 S.n3780 0.003
R48655 S.n3044 S.n3043 0.003
R48656 S.n920 S.n919 0.003
R48657 S.n1988 S.n1987 0.003
R48658 S.n22747 S.n22746 0.003
R48659 S.n21320 S.n21319 0.003
R48660 S.n21223 S.n21222 0.003
R48661 S.n20497 S.n20496 0.003
R48662 S.n20404 S.n20403 0.003
R48663 S.n19886 S.n19885 0.003
R48664 S.n20274 S.n20273 0.003
R48665 S.n19032 S.n19031 0.003
R48666 S.n19406 S.n19405 0.003
R48667 S.n18166 S.n18165 0.003
R48668 S.n18519 S.n18518 0.003
R48669 S.n17277 S.n17276 0.003
R48670 S.n17619 S.n17618 0.003
R48671 S.n16375 S.n16374 0.003
R48672 S.n16696 S.n16695 0.003
R48673 S.n15451 S.n15450 0.003
R48674 S.n15761 S.n15760 0.003
R48675 S.n14514 S.n14513 0.003
R48676 S.n14803 S.n14802 0.003
R48677 S.n13555 S.n13554 0.003
R48678 S.n13833 S.n13832 0.003
R48679 S.n12583 S.n12582 0.003
R48680 S.n12840 S.n12839 0.003
R48681 S.n11589 S.n11588 0.003
R48682 S.n11835 S.n11834 0.003
R48683 S.n10582 S.n10581 0.003
R48684 S.n10807 S.n10806 0.003
R48685 S.n9553 S.n9552 0.003
R48686 S.n9767 S.n9766 0.003
R48687 S.n8511 S.n8510 0.003
R48688 S.n8704 S.n8703 0.003
R48689 S.n7447 S.n7446 0.003
R48690 S.n7629 S.n7628 0.003
R48691 S.n6370 S.n6369 0.003
R48692 S.n6531 S.n6530 0.003
R48693 S.n5270 S.n5269 0.003
R48694 S.n5420 S.n5419 0.003
R48695 S.n4157 S.n4156 0.003
R48696 S.n4286 S.n4285 0.003
R48697 S.n3031 S.n3030 0.003
R48698 S.n3149 S.n3148 0.003
R48699 S.n1871 S.n1870 0.003
R48700 S.n877 S.n876 0.003
R48701 S.n809 S.n808 0.003
R48702 S.n977 S.n976 0.003
R48703 S.n22354 S.n22353 0.003
R48704 S.n22719 S.n22718 0.003
R48705 S.n21348 S.n21347 0.003
R48706 S.n21264 S.n21263 0.003
R48707 S.n20827 S.n20826 0.003
R48708 S.n20848 S.n20847 0.003
R48709 S.n20192 S.n20191 0.003
R48710 S.n20216 S.n20215 0.003
R48711 S.n19322 S.n19321 0.003
R48712 S.n19346 S.n19345 0.003
R48713 S.n18440 S.n18439 0.003
R48714 S.n18464 S.n18463 0.003
R48715 S.n17535 S.n17534 0.003
R48716 S.n17559 S.n17558 0.003
R48717 S.n16617 S.n16616 0.003
R48718 S.n16641 S.n16640 0.003
R48719 S.n15677 S.n15676 0.003
R48720 S.n15701 S.n15700 0.003
R48721 S.n14724 S.n14723 0.003
R48722 S.n14748 S.n14747 0.003
R48723 S.n13749 S.n13748 0.003
R48724 S.n13773 S.n13772 0.003
R48725 S.n12761 S.n12760 0.003
R48726 S.n12785 S.n12784 0.003
R48727 S.n11751 S.n11750 0.003
R48728 S.n11775 S.n11774 0.003
R48729 S.n10728 S.n10727 0.003
R48730 S.n10752 S.n10751 0.003
R48731 S.n9683 S.n9682 0.003
R48732 S.n9707 S.n9706 0.003
R48733 S.n8625 S.n8624 0.003
R48734 S.n8649 S.n8648 0.003
R48735 S.n7545 S.n7544 0.003
R48736 S.n7569 S.n7568 0.003
R48737 S.n6452 S.n6451 0.003
R48738 S.n6476 S.n6475 0.003
R48739 S.n5336 S.n5335 0.003
R48740 S.n5360 S.n5359 0.003
R48741 S.n4207 S.n4206 0.003
R48742 S.n4231 S.n4230 0.003
R48743 S.n3066 S.n3065 0.003
R48744 S.n3090 S.n3089 0.003
R48745 S.n1885 S.n1884 0.003
R48746 S.n1937 S.n1936 0.003
R48747 S.n412 S.n411 0.003
R48748 S.n2140 S.n2139 0.003
R48749 S.n18489 S.n18488 0.003
R48750 S.n17175 S.n17174 0.003
R48751 S.n17768 S.n17767 0.003
R48752 S.n16275 S.n16274 0.003
R48753 S.n16841 S.n16840 0.003
R48754 S.n15351 S.n15350 0.003
R48755 S.n15906 S.n15905 0.003
R48756 S.n14414 S.n14413 0.003
R48757 S.n14948 S.n14947 0.003
R48758 S.n13455 S.n13454 0.003
R48759 S.n13978 S.n13977 0.003
R48760 S.n12483 S.n12482 0.003
R48761 S.n12985 S.n12984 0.003
R48762 S.n11489 S.n11488 0.003
R48763 S.n11980 S.n11979 0.003
R48764 S.n10482 S.n10481 0.003
R48765 S.n10952 S.n10951 0.003
R48766 S.n9453 S.n9452 0.003
R48767 S.n9912 S.n9911 0.003
R48768 S.n8411 S.n8410 0.003
R48769 S.n8849 S.n8848 0.003
R48770 S.n7347 S.n7346 0.003
R48771 S.n7774 S.n7773 0.003
R48772 S.n6270 S.n6269 0.003
R48773 S.n6676 S.n6675 0.003
R48774 S.n5170 S.n5169 0.003
R48775 S.n5566 S.n5565 0.003
R48776 S.n4058 S.n4057 0.003
R48777 S.n4431 S.n4430 0.003
R48778 S.n2931 S.n2930 0.003
R48779 S.n3293 S.n3292 0.003
R48780 S.n1763 S.n1762 0.003
R48781 S.n16 S.n15 0.003
R48782 S.n19376 S.n19375 0.003
R48783 S.n18083 S.n18082 0.003
R48784 S.n18636 S.n18635 0.003
R48785 S.n17194 S.n17193 0.003
R48786 S.n17736 S.n17735 0.003
R48787 S.n16292 S.n16291 0.003
R48788 S.n16809 S.n16808 0.003
R48789 S.n15368 S.n15367 0.003
R48790 S.n15874 S.n15873 0.003
R48791 S.n14431 S.n14430 0.003
R48792 S.n14916 S.n14915 0.003
R48793 S.n13472 S.n13471 0.003
R48794 S.n13946 S.n13945 0.003
R48795 S.n12500 S.n12499 0.003
R48796 S.n12953 S.n12952 0.003
R48797 S.n11506 S.n11505 0.003
R48798 S.n11948 S.n11947 0.003
R48799 S.n10499 S.n10498 0.003
R48800 S.n10920 S.n10919 0.003
R48801 S.n9470 S.n9469 0.003
R48802 S.n9880 S.n9879 0.003
R48803 S.n8428 S.n8427 0.003
R48804 S.n8817 S.n8816 0.003
R48805 S.n7364 S.n7363 0.003
R48806 S.n7742 S.n7741 0.003
R48807 S.n6287 S.n6286 0.003
R48808 S.n6644 S.n6643 0.003
R48809 S.n5187 S.n5186 0.003
R48810 S.n5534 S.n5533 0.003
R48811 S.n4075 S.n4074 0.003
R48812 S.n4399 S.n4398 0.003
R48813 S.n2948 S.n2947 0.003
R48814 S.n3262 S.n3261 0.003
R48815 S.n1782 S.n1781 0.003
R48816 S.n1805 S.n1804 0.003
R48817 S.n2082 S.n2081 0.003
R48818 S.n815 S.n814 0.003
R48819 S.n844 S.n843 0.003
R48820 S.n3233 S.n3232 0.003
R48821 S.n4370 S.n4369 0.003
R48822 S.n5505 S.n5504 0.003
R48823 S.n6615 S.n6614 0.003
R48824 S.n7713 S.n7712 0.003
R48825 S.n8788 S.n8787 0.003
R48826 S.n9851 S.n9850 0.003
R48827 S.n10891 S.n10890 0.003
R48828 S.n11919 S.n11918 0.003
R48829 S.n12924 S.n12923 0.003
R48830 S.n13917 S.n13916 0.003
R48831 S.n14887 S.n14886 0.003
R48832 S.n15845 S.n15844 0.003
R48833 S.n16780 S.n16779 0.003
R48834 S.n17703 S.n17702 0.003
R48835 S.n18603 S.n18602 0.003
R48836 S.n19493 S.n19492 0.003
R48837 S.n20244 S.n20243 0.003
R48838 S.n18967 S.n18966 0.003
R48839 S.n18102 S.n18101 0.003
R48840 S.n17213 S.n17212 0.003
R48841 S.n16311 S.n16310 0.003
R48842 S.n15387 S.n15386 0.003
R48843 S.n14450 S.n14449 0.003
R48844 S.n13491 S.n13490 0.003
R48845 S.n12519 S.n12518 0.003
R48846 S.n11525 S.n11524 0.003
R48847 S.n10518 S.n10517 0.003
R48848 S.n9489 S.n9488 0.003
R48849 S.n8447 S.n8446 0.003
R48850 S.n7383 S.n7382 0.003
R48851 S.n6306 S.n6305 0.003
R48852 S.n5206 S.n5205 0.003
R48853 S.n4094 S.n4093 0.003
R48854 S.n2967 S.n2966 0.003
R48855 S.n2048 S.n2047 0.003
R48856 S.n773 S.n772 0.003
R48857 S.n1328 S.n1327 0.003
R48858 S.n20427 S.n20426 0.003
R48859 S.n19845 S.n19844 0.003
R48860 S.n20333 S.n20332 0.003
R48861 S.n18993 S.n18992 0.003
R48862 S.n19461 S.n19460 0.003
R48863 S.n18127 S.n18126 0.003
R48864 S.n18571 S.n18570 0.003
R48865 S.n17238 S.n17237 0.003
R48866 S.n17671 S.n17670 0.003
R48867 S.n16336 S.n16335 0.003
R48868 S.n16748 S.n16747 0.003
R48869 S.n15412 S.n15411 0.003
R48870 S.n15813 S.n15812 0.003
R48871 S.n14475 S.n14474 0.003
R48872 S.n14855 S.n14854 0.003
R48873 S.n13516 S.n13515 0.003
R48874 S.n13885 S.n13884 0.003
R48875 S.n12544 S.n12543 0.003
R48876 S.n12892 S.n12891 0.003
R48877 S.n11550 S.n11549 0.003
R48878 S.n11887 S.n11886 0.003
R48879 S.n10543 S.n10542 0.003
R48880 S.n10859 S.n10858 0.003
R48881 S.n9514 S.n9513 0.003
R48882 S.n9819 S.n9818 0.003
R48883 S.n8472 S.n8471 0.003
R48884 S.n8756 S.n8755 0.003
R48885 S.n7408 S.n7407 0.003
R48886 S.n7681 S.n7680 0.003
R48887 S.n6331 S.n6330 0.003
R48888 S.n6583 S.n6582 0.003
R48889 S.n5231 S.n5230 0.003
R48890 S.n5473 S.n5472 0.003
R48891 S.n4119 S.n4118 0.003
R48892 S.n4338 S.n4337 0.003
R48893 S.n2992 S.n2991 0.003
R48894 S.n3201 S.n3200 0.003
R48895 S.n1829 S.n1828 0.003
R48896 S.n2015 S.n2014 0.003
R48897 S.n792 S.n791 0.003
R48898 S.n1851 S.n1850 0.003
R48899 S.n3169 S.n3168 0.003
R48900 S.n3012 S.n3011 0.003
R48901 S.n4306 S.n4305 0.003
R48902 S.n4138 S.n4137 0.003
R48903 S.n5441 S.n5440 0.003
R48904 S.n5251 S.n5250 0.003
R48905 S.n6551 S.n6550 0.003
R48906 S.n6351 S.n6350 0.003
R48907 S.n7649 S.n7648 0.003
R48908 S.n7428 S.n7427 0.003
R48909 S.n8724 S.n8723 0.003
R48910 S.n8492 S.n8491 0.003
R48911 S.n9787 S.n9786 0.003
R48912 S.n9534 S.n9533 0.003
R48913 S.n10827 S.n10826 0.003
R48914 S.n10563 S.n10562 0.003
R48915 S.n11855 S.n11854 0.003
R48916 S.n11570 S.n11569 0.003
R48917 S.n12860 S.n12859 0.003
R48918 S.n12564 S.n12563 0.003
R48919 S.n13853 S.n13852 0.003
R48920 S.n13536 S.n13535 0.003
R48921 S.n14823 S.n14822 0.003
R48922 S.n14495 S.n14494 0.003
R48923 S.n15781 S.n15780 0.003
R48924 S.n15432 S.n15431 0.003
R48925 S.n16716 S.n16715 0.003
R48926 S.n16356 S.n16355 0.003
R48927 S.n17639 S.n17638 0.003
R48928 S.n17258 S.n17257 0.003
R48929 S.n18539 S.n18538 0.003
R48930 S.n18147 S.n18146 0.003
R48931 S.n19426 S.n19425 0.003
R48932 S.n19013 S.n19012 0.003
R48933 S.n20298 S.n20297 0.003
R48934 S.n19867 S.n19866 0.003
R48935 S.n20372 S.n20371 0.003
R48936 S.n20478 S.n20477 0.003
R48937 S.n21245 S.n21244 0.003
R48938 S.n870 S.n869 0.003
R48939 S.n2110 S.n2109 0.003
R48940 S.n749 S.n748 0.003
R48941 S.n732 S.n731 0.003
R48942 S.n380 S.n379 0.003
R48943 S.n2199 S.n2198 0.003
R48944 S.n16666 S.n16665 0.003
R48945 S.n15313 S.n15312 0.003
R48946 S.n15971 S.n15970 0.003
R48947 S.n14378 S.n14377 0.003
R48948 S.n15009 S.n15008 0.003
R48949 S.n13419 S.n13418 0.003
R48950 S.n14039 S.n14038 0.003
R48951 S.n12447 S.n12446 0.003
R48952 S.n13046 S.n13045 0.003
R48953 S.n11453 S.n11452 0.003
R48954 S.n12041 S.n12040 0.003
R48955 S.n10446 S.n10445 0.003
R48956 S.n11013 S.n11012 0.003
R48957 S.n9417 S.n9416 0.003
R48958 S.n9973 S.n9972 0.003
R48959 S.n8375 S.n8374 0.003
R48960 S.n8910 S.n8909 0.003
R48961 S.n7311 S.n7310 0.003
R48962 S.n7835 S.n7834 0.003
R48963 S.n6234 S.n6233 0.003
R48964 S.n6737 S.n6736 0.003
R48965 S.n5134 S.n5133 0.003
R48966 S.n5627 S.n5626 0.003
R48967 S.n4022 S.n4021 0.003
R48968 S.n4492 S.n4491 0.003
R48969 S.n2895 S.n2894 0.003
R48970 S.n3353 S.n3352 0.003
R48971 S.n1726 S.n1725 0.003
R48972 S.n63 S.n62 0.003
R48973 S.n17589 S.n17588 0.003
R48974 S.n16256 S.n16255 0.003
R48975 S.n16874 S.n16873 0.003
R48976 S.n15332 S.n15331 0.003
R48977 S.n15939 S.n15938 0.003
R48978 S.n14395 S.n14394 0.003
R48979 S.n14977 S.n14976 0.003
R48980 S.n13436 S.n13435 0.003
R48981 S.n14007 S.n14006 0.003
R48982 S.n12464 S.n12463 0.003
R48983 S.n13014 S.n13013 0.003
R48984 S.n11470 S.n11469 0.003
R48985 S.n12009 S.n12008 0.003
R48986 S.n10463 S.n10462 0.003
R48987 S.n10981 S.n10980 0.003
R48988 S.n9434 S.n9433 0.003
R48989 S.n9941 S.n9940 0.003
R48990 S.n8392 S.n8391 0.003
R48991 S.n8878 S.n8877 0.003
R48992 S.n7328 S.n7327 0.003
R48993 S.n7803 S.n7802 0.003
R48994 S.n6251 S.n6250 0.003
R48995 S.n6705 S.n6704 0.003
R48996 S.n5151 S.n5150 0.003
R48997 S.n5595 S.n5594 0.003
R48998 S.n4039 S.n4038 0.003
R48999 S.n4460 S.n4459 0.003
R49000 S.n2912 S.n2911 0.003
R49001 S.n3322 S.n3321 0.003
R49002 S.n1743 S.n1742 0.003
R49003 S.n2169 S.n2168 0.003
R49004 S.n714 S.n713 0.003
R49005 S.n697 S.n696 0.003
R49006 S.n348 S.n347 0.003
R49007 S.n2258 S.n2257 0.003
R49008 S.n14773 S.n14772 0.003
R49009 S.n13381 S.n13380 0.003
R49010 S.n14104 S.n14103 0.003
R49011 S.n12411 S.n12410 0.003
R49012 S.n13107 S.n13106 0.003
R49013 S.n11417 S.n11416 0.003
R49014 S.n12102 S.n12101 0.003
R49015 S.n10410 S.n10409 0.003
R49016 S.n11074 S.n11073 0.003
R49017 S.n9381 S.n9380 0.003
R49018 S.n10034 S.n10033 0.003
R49019 S.n8339 S.n8338 0.003
R49020 S.n8971 S.n8970 0.003
R49021 S.n7275 S.n7274 0.003
R49022 S.n7896 S.n7895 0.003
R49023 S.n6198 S.n6197 0.003
R49024 S.n6798 S.n6797 0.003
R49025 S.n5098 S.n5097 0.003
R49026 S.n5688 S.n5687 0.003
R49027 S.n3986 S.n3985 0.003
R49028 S.n4553 S.n4552 0.003
R49029 S.n2859 S.n2858 0.003
R49030 S.n3413 S.n3412 0.003
R49031 S.n1689 S.n1688 0.003
R49032 S.n95 S.n94 0.003
R49033 S.n15731 S.n15730 0.003
R49034 S.n14359 S.n14358 0.003
R49035 S.n15042 S.n15041 0.003
R49036 S.n13400 S.n13399 0.003
R49037 S.n14072 S.n14071 0.003
R49038 S.n12428 S.n12427 0.003
R49039 S.n13075 S.n13074 0.003
R49040 S.n11434 S.n11433 0.003
R49041 S.n12070 S.n12069 0.003
R49042 S.n10427 S.n10426 0.003
R49043 S.n11042 S.n11041 0.003
R49044 S.n9398 S.n9397 0.003
R49045 S.n10002 S.n10001 0.003
R49046 S.n8356 S.n8355 0.003
R49047 S.n8939 S.n8938 0.003
R49048 S.n7292 S.n7291 0.003
R49049 S.n7864 S.n7863 0.003
R49050 S.n6215 S.n6214 0.003
R49051 S.n6766 S.n6765 0.003
R49052 S.n5115 S.n5114 0.003
R49053 S.n5656 S.n5655 0.003
R49054 S.n4003 S.n4002 0.003
R49055 S.n4521 S.n4520 0.003
R49056 S.n2876 S.n2875 0.003
R49057 S.n3382 S.n3381 0.003
R49058 S.n1706 S.n1705 0.003
R49059 S.n2228 S.n2227 0.003
R49060 S.n679 S.n678 0.003
R49061 S.n662 S.n661 0.003
R49062 S.n316 S.n315 0.003
R49063 S.n2317 S.n2316 0.003
R49064 S.n12810 S.n12809 0.003
R49065 S.n11379 S.n11378 0.003
R49066 S.n12167 S.n12166 0.003
R49067 S.n10374 S.n10373 0.003
R49068 S.n11135 S.n11134 0.003
R49069 S.n9345 S.n9344 0.003
R49070 S.n10095 S.n10094 0.003
R49071 S.n8303 S.n8302 0.003
R49072 S.n9032 S.n9031 0.003
R49073 S.n7239 S.n7238 0.003
R49074 S.n7957 S.n7956 0.003
R49075 S.n6162 S.n6161 0.003
R49076 S.n6859 S.n6858 0.003
R49077 S.n5062 S.n5061 0.003
R49078 S.n5749 S.n5748 0.003
R49079 S.n3950 S.n3949 0.003
R49080 S.n4614 S.n4613 0.003
R49081 S.n2823 S.n2822 0.003
R49082 S.n3473 S.n3472 0.003
R49083 S.n1652 S.n1651 0.003
R49084 S.n982 S.n981 0.003
R49085 S.n13803 S.n13802 0.003
R49086 S.n12392 S.n12391 0.003
R49087 S.n13140 S.n13139 0.003
R49088 S.n11398 S.n11397 0.003
R49089 S.n12135 S.n12134 0.003
R49090 S.n10391 S.n10390 0.003
R49091 S.n11103 S.n11102 0.003
R49092 S.n9362 S.n9361 0.003
R49093 S.n10063 S.n10062 0.003
R49094 S.n8320 S.n8319 0.003
R49095 S.n9000 S.n8999 0.003
R49096 S.n7256 S.n7255 0.003
R49097 S.n7925 S.n7924 0.003
R49098 S.n6179 S.n6178 0.003
R49099 S.n6827 S.n6826 0.003
R49100 S.n5079 S.n5078 0.003
R49101 S.n5717 S.n5716 0.003
R49102 S.n3967 S.n3966 0.003
R49103 S.n4582 S.n4581 0.003
R49104 S.n2840 S.n2839 0.003
R49105 S.n3442 S.n3441 0.003
R49106 S.n1669 S.n1668 0.003
R49107 S.n2287 S.n2286 0.003
R49108 S.n644 S.n643 0.003
R49109 S.n627 S.n626 0.003
R49110 S.n284 S.n283 0.003
R49111 S.n2376 S.n2375 0.003
R49112 S.n10777 S.n10776 0.003
R49113 S.n9307 S.n9306 0.003
R49114 S.n10160 S.n10159 0.003
R49115 S.n8267 S.n8266 0.003
R49116 S.n9093 S.n9092 0.003
R49117 S.n7203 S.n7202 0.003
R49118 S.n8018 S.n8017 0.003
R49119 S.n6126 S.n6125 0.003
R49120 S.n6920 S.n6919 0.003
R49121 S.n5026 S.n5025 0.003
R49122 S.n5810 S.n5809 0.003
R49123 S.n3914 S.n3913 0.003
R49124 S.n4675 S.n4674 0.003
R49125 S.n2787 S.n2786 0.003
R49126 S.n3533 S.n3532 0.003
R49127 S.n1615 S.n1614 0.003
R49128 S.n1014 S.n1013 0.003
R49129 S.n11805 S.n11804 0.003
R49130 S.n10355 S.n10354 0.003
R49131 S.n11168 S.n11167 0.003
R49132 S.n9326 S.n9325 0.003
R49133 S.n10128 S.n10127 0.003
R49134 S.n8284 S.n8283 0.003
R49135 S.n9061 S.n9060 0.003
R49136 S.n7220 S.n7219 0.003
R49137 S.n7986 S.n7985 0.003
R49138 S.n6143 S.n6142 0.003
R49139 S.n6888 S.n6887 0.003
R49140 S.n5043 S.n5042 0.003
R49141 S.n5778 S.n5777 0.003
R49142 S.n3931 S.n3930 0.003
R49143 S.n4643 S.n4642 0.003
R49144 S.n2804 S.n2803 0.003
R49145 S.n3502 S.n3501 0.003
R49146 S.n1632 S.n1631 0.003
R49147 S.n2346 S.n2345 0.003
R49148 S.n609 S.n608 0.003
R49149 S.n592 S.n591 0.003
R49150 S.n252 S.n251 0.003
R49151 S.n2435 S.n2434 0.003
R49152 S.n8674 S.n8673 0.003
R49153 S.n7165 S.n7164 0.003
R49154 S.n8083 S.n8082 0.003
R49155 S.n6090 S.n6089 0.003
R49156 S.n6981 S.n6980 0.003
R49157 S.n4990 S.n4989 0.003
R49158 S.n5871 S.n5870 0.003
R49159 S.n3878 S.n3877 0.003
R49160 S.n4736 S.n4735 0.003
R49161 S.n2751 S.n2750 0.003
R49162 S.n3593 S.n3592 0.003
R49163 S.n1578 S.n1577 0.003
R49164 S.n1046 S.n1045 0.003
R49165 S.n9737 S.n9736 0.003
R49166 S.n8248 S.n8247 0.003
R49167 S.n9126 S.n9125 0.003
R49168 S.n7184 S.n7183 0.003
R49169 S.n8051 S.n8050 0.003
R49170 S.n6107 S.n6106 0.003
R49171 S.n6949 S.n6948 0.003
R49172 S.n5007 S.n5006 0.003
R49173 S.n5839 S.n5838 0.003
R49174 S.n3895 S.n3894 0.003
R49175 S.n4704 S.n4703 0.003
R49176 S.n2768 S.n2767 0.003
R49177 S.n3562 S.n3561 0.003
R49178 S.n1595 S.n1594 0.003
R49179 S.n2405 S.n2404 0.003
R49180 S.n574 S.n573 0.003
R49181 S.n557 S.n556 0.003
R49182 S.n220 S.n219 0.003
R49183 S.n2494 S.n2493 0.003
R49184 S.n6501 S.n6500 0.003
R49185 S.n4952 S.n4951 0.003
R49186 S.n5936 S.n5935 0.003
R49187 S.n3842 S.n3841 0.003
R49188 S.n4797 S.n4796 0.003
R49189 S.n2715 S.n2714 0.003
R49190 S.n3653 S.n3652 0.003
R49191 S.n1541 S.n1540 0.003
R49192 S.n1078 S.n1077 0.003
R49193 S.n7599 S.n7598 0.003
R49194 S.n6071 S.n6070 0.003
R49195 S.n7014 S.n7013 0.003
R49196 S.n4971 S.n4970 0.003
R49197 S.n5904 S.n5903 0.003
R49198 S.n3859 S.n3858 0.003
R49199 S.n4765 S.n4764 0.003
R49200 S.n2732 S.n2731 0.003
R49201 S.n3622 S.n3621 0.003
R49202 S.n1558 S.n1557 0.003
R49203 S.n2464 S.n2463 0.003
R49204 S.n539 S.n538 0.003
R49205 S.n522 S.n521 0.003
R49206 S.n188 S.n187 0.003
R49207 S.n2553 S.n2552 0.003
R49208 S.n4256 S.n4255 0.003
R49209 S.n2677 S.n2676 0.003
R49210 S.n3717 S.n3716 0.003
R49211 S.n1504 S.n1503 0.003
R49212 S.n1110 S.n1109 0.003
R49213 S.n5390 S.n5389 0.003
R49214 S.n3823 S.n3822 0.003
R49215 S.n4830 S.n4829 0.003
R49216 S.n2696 S.n2695 0.003
R49217 S.n3686 S.n3685 0.003
R49218 S.n1521 S.n1520 0.003
R49219 S.n2523 S.n2522 0.003
R49220 S.n504 S.n503 0.003
R49221 S.n487 S.n486 0.003
R49222 S.n156 S.n155 0.003
R49223 S.n1960 S.n1959 0.003
R49224 S.n1148 S.n1147 0.003
R49225 S.n3120 S.n3119 0.003
R49226 S.n1484 S.n1483 0.003
R49227 S.n2586 S.n2585 0.003
R49228 S.n469 S.n468 0.003
R49229 S.n453 S.n452 0.003
R49230 S.n945 S.n944 0.003
R49231 S.n22313 S.n22312 0.003
R49232 S.n21971 S.n21970 0.003
R49233 S.n22768 S.n22767 0.003
R49234 S.n21334 S.n21333 0.003
R49235 S.n22339 S.n22338 0.003
R49236 S.n1776 S.n1775 0.003
R49237 S.n20183 S.n20178 0.003
R49238 S.n21133 S.n21132 0.003
R49239 S.n22640 S.n22638 0.003
R49240 S.n22010 S.n22009 0.003
R49241 S.n21617 S.n21615 0.003
R49242 S.n21942 S.n21941 0.003
R49243 S.n20794 S.n20792 0.003
R49244 S.n22656 S.n22651 0.003
R49245 S.n21995 S.n21990 0.003
R49246 S.n21638 S.n21633 0.003
R49247 S.n21962 S.n21956 0.003
R49248 S.n20818 S.n20810 0.003
R49249 S.n19313 S.n19308 0.003
R49250 S.n19533 S.n19532 0.003
R49251 S.n22624 S.n22622 0.003
R49252 S.n22025 S.n22024 0.003
R49253 S.n21601 S.n21599 0.003
R49254 S.n21927 S.n21926 0.003
R49255 S.n20778 S.n20776 0.003
R49256 S.n21117 S.n21116 0.003
R49257 S.n20167 S.n20165 0.003
R49258 S.n18431 S.n18426 0.003
R49259 S.n18676 S.n18675 0.003
R49260 S.n22608 S.n22606 0.003
R49261 S.n22040 S.n22039 0.003
R49262 S.n21585 S.n21583 0.003
R49263 S.n21912 S.n21911 0.003
R49264 S.n20762 S.n20760 0.003
R49265 S.n21102 S.n21101 0.003
R49266 S.n20151 S.n20149 0.003
R49267 S.n19548 S.n19547 0.003
R49268 S.n19297 S.n19295 0.003
R49269 S.n17526 S.n17521 0.003
R49270 S.n17808 S.n17807 0.003
R49271 S.n22592 S.n22590 0.003
R49272 S.n22055 S.n22054 0.003
R49273 S.n21569 S.n21567 0.003
R49274 S.n21897 S.n21896 0.003
R49275 S.n20746 S.n20744 0.003
R49276 S.n21087 S.n21086 0.003
R49277 S.n20135 S.n20133 0.003
R49278 S.n19563 S.n19562 0.003
R49279 S.n19281 S.n19279 0.003
R49280 S.n18691 S.n18690 0.003
R49281 S.n18415 S.n18413 0.003
R49282 S.n16608 S.n16603 0.003
R49283 S.n16914 S.n16913 0.003
R49284 S.n22576 S.n22574 0.003
R49285 S.n22070 S.n22069 0.003
R49286 S.n21553 S.n21551 0.003
R49287 S.n21882 S.n21881 0.003
R49288 S.n20730 S.n20728 0.003
R49289 S.n21072 S.n21071 0.003
R49290 S.n20119 S.n20117 0.003
R49291 S.n19578 S.n19577 0.003
R49292 S.n19265 S.n19263 0.003
R49293 S.n18706 S.n18705 0.003
R49294 S.n18399 S.n18397 0.003
R49295 S.n17823 S.n17822 0.003
R49296 S.n17510 S.n17508 0.003
R49297 S.n15668 S.n15663 0.003
R49298 S.n16011 S.n16010 0.003
R49299 S.n22560 S.n22558 0.003
R49300 S.n22085 S.n22084 0.003
R49301 S.n21537 S.n21535 0.003
R49302 S.n21867 S.n21866 0.003
R49303 S.n20714 S.n20712 0.003
R49304 S.n21057 S.n21056 0.003
R49305 S.n20103 S.n20101 0.003
R49306 S.n19593 S.n19592 0.003
R49307 S.n19249 S.n19247 0.003
R49308 S.n18721 S.n18720 0.003
R49309 S.n18383 S.n18381 0.003
R49310 S.n17838 S.n17837 0.003
R49311 S.n17494 S.n17492 0.003
R49312 S.n16929 S.n16928 0.003
R49313 S.n16592 S.n16590 0.003
R49314 S.n14715 S.n14710 0.003
R49315 S.n15082 S.n15081 0.003
R49316 S.n22544 S.n22542 0.003
R49317 S.n22100 S.n22099 0.003
R49318 S.n21521 S.n21519 0.003
R49319 S.n21852 S.n21851 0.003
R49320 S.n20698 S.n20696 0.003
R49321 S.n21042 S.n21041 0.003
R49322 S.n20087 S.n20085 0.003
R49323 S.n19608 S.n19607 0.003
R49324 S.n19233 S.n19231 0.003
R49325 S.n18736 S.n18735 0.003
R49326 S.n18367 S.n18365 0.003
R49327 S.n17853 S.n17852 0.003
R49328 S.n17478 S.n17476 0.003
R49329 S.n16944 S.n16943 0.003
R49330 S.n16576 S.n16574 0.003
R49331 S.n16026 S.n16025 0.003
R49332 S.n15652 S.n15650 0.003
R49333 S.n13740 S.n13735 0.003
R49334 S.n14144 S.n14143 0.003
R49335 S.n22528 S.n22526 0.003
R49336 S.n22115 S.n22114 0.003
R49337 S.n21505 S.n21503 0.003
R49338 S.n21837 S.n21836 0.003
R49339 S.n20682 S.n20680 0.003
R49340 S.n21027 S.n21026 0.003
R49341 S.n20071 S.n20069 0.003
R49342 S.n19623 S.n19622 0.003
R49343 S.n19217 S.n19215 0.003
R49344 S.n18751 S.n18750 0.003
R49345 S.n18351 S.n18349 0.003
R49346 S.n17868 S.n17867 0.003
R49347 S.n17462 S.n17460 0.003
R49348 S.n16959 S.n16958 0.003
R49349 S.n16560 S.n16558 0.003
R49350 S.n16041 S.n16040 0.003
R49351 S.n15636 S.n15634 0.003
R49352 S.n15097 S.n15096 0.003
R49353 S.n14699 S.n14697 0.003
R49354 S.n12752 S.n12747 0.003
R49355 S.n13180 S.n13179 0.003
R49356 S.n22512 S.n22510 0.003
R49357 S.n22130 S.n22129 0.003
R49358 S.n21489 S.n21487 0.003
R49359 S.n21822 S.n21821 0.003
R49360 S.n20666 S.n20664 0.003
R49361 S.n21012 S.n21011 0.003
R49362 S.n20055 S.n20053 0.003
R49363 S.n19638 S.n19637 0.003
R49364 S.n19201 S.n19199 0.003
R49365 S.n18766 S.n18765 0.003
R49366 S.n18335 S.n18333 0.003
R49367 S.n17883 S.n17882 0.003
R49368 S.n17446 S.n17444 0.003
R49369 S.n16974 S.n16973 0.003
R49370 S.n16544 S.n16542 0.003
R49371 S.n16056 S.n16055 0.003
R49372 S.n15620 S.n15618 0.003
R49373 S.n15112 S.n15111 0.003
R49374 S.n14683 S.n14681 0.003
R49375 S.n14159 S.n14158 0.003
R49376 S.n13724 S.n13722 0.003
R49377 S.n11742 S.n11737 0.003
R49378 S.n12207 S.n12206 0.003
R49379 S.n22496 S.n22494 0.003
R49380 S.n22145 S.n22144 0.003
R49381 S.n21473 S.n21471 0.003
R49382 S.n21807 S.n21806 0.003
R49383 S.n20650 S.n20648 0.003
R49384 S.n20997 S.n20996 0.003
R49385 S.n20039 S.n20037 0.003
R49386 S.n19653 S.n19652 0.003
R49387 S.n19185 S.n19183 0.003
R49388 S.n18781 S.n18780 0.003
R49389 S.n18319 S.n18317 0.003
R49390 S.n17898 S.n17897 0.003
R49391 S.n17430 S.n17428 0.003
R49392 S.n16989 S.n16988 0.003
R49393 S.n16528 S.n16526 0.003
R49394 S.n16071 S.n16070 0.003
R49395 S.n15604 S.n15602 0.003
R49396 S.n15127 S.n15126 0.003
R49397 S.n14667 S.n14665 0.003
R49398 S.n14174 S.n14173 0.003
R49399 S.n13708 S.n13706 0.003
R49400 S.n13195 S.n13194 0.003
R49401 S.n12736 S.n12734 0.003
R49402 S.n10719 S.n10714 0.003
R49403 S.n11208 S.n11207 0.003
R49404 S.n22480 S.n22478 0.003
R49405 S.n22160 S.n22159 0.003
R49406 S.n21457 S.n21455 0.003
R49407 S.n21792 S.n21791 0.003
R49408 S.n20634 S.n20632 0.003
R49409 S.n20982 S.n20981 0.003
R49410 S.n20023 S.n20021 0.003
R49411 S.n19668 S.n19667 0.003
R49412 S.n19169 S.n19167 0.003
R49413 S.n18796 S.n18795 0.003
R49414 S.n18303 S.n18301 0.003
R49415 S.n17913 S.n17912 0.003
R49416 S.n17414 S.n17412 0.003
R49417 S.n17004 S.n17003 0.003
R49418 S.n16512 S.n16510 0.003
R49419 S.n16086 S.n16085 0.003
R49420 S.n15588 S.n15586 0.003
R49421 S.n15142 S.n15141 0.003
R49422 S.n14651 S.n14649 0.003
R49423 S.n14189 S.n14188 0.003
R49424 S.n13692 S.n13690 0.003
R49425 S.n13210 S.n13209 0.003
R49426 S.n12720 S.n12718 0.003
R49427 S.n12222 S.n12221 0.003
R49428 S.n11726 S.n11724 0.003
R49429 S.n9674 S.n9669 0.003
R49430 S.n10200 S.n10199 0.003
R49431 S.n22464 S.n22462 0.003
R49432 S.n22175 S.n22174 0.003
R49433 S.n21441 S.n21439 0.003
R49434 S.n21777 S.n21776 0.003
R49435 S.n20618 S.n20616 0.003
R49436 S.n20967 S.n20966 0.003
R49437 S.n20007 S.n20005 0.003
R49438 S.n19683 S.n19682 0.003
R49439 S.n19153 S.n19151 0.003
R49440 S.n18811 S.n18810 0.003
R49441 S.n18287 S.n18285 0.003
R49442 S.n17928 S.n17927 0.003
R49443 S.n17398 S.n17396 0.003
R49444 S.n17019 S.n17018 0.003
R49445 S.n16496 S.n16494 0.003
R49446 S.n16101 S.n16100 0.003
R49447 S.n15572 S.n15570 0.003
R49448 S.n15157 S.n15156 0.003
R49449 S.n14635 S.n14633 0.003
R49450 S.n14204 S.n14203 0.003
R49451 S.n13676 S.n13674 0.003
R49452 S.n13225 S.n13224 0.003
R49453 S.n12704 S.n12702 0.003
R49454 S.n12237 S.n12236 0.003
R49455 S.n11710 S.n11708 0.003
R49456 S.n11223 S.n11222 0.003
R49457 S.n10703 S.n10701 0.003
R49458 S.n8616 S.n8611 0.003
R49459 S.n9166 S.n9165 0.003
R49460 S.n22448 S.n22446 0.003
R49461 S.n22190 S.n22189 0.003
R49462 S.n21425 S.n21423 0.003
R49463 S.n21762 S.n21761 0.003
R49464 S.n20602 S.n20600 0.003
R49465 S.n20952 S.n20951 0.003
R49466 S.n19991 S.n19989 0.003
R49467 S.n19698 S.n19697 0.003
R49468 S.n19137 S.n19135 0.003
R49469 S.n18826 S.n18825 0.003
R49470 S.n18271 S.n18269 0.003
R49471 S.n17943 S.n17942 0.003
R49472 S.n17382 S.n17380 0.003
R49473 S.n17034 S.n17033 0.003
R49474 S.n16480 S.n16478 0.003
R49475 S.n16116 S.n16115 0.003
R49476 S.n15556 S.n15554 0.003
R49477 S.n15172 S.n15171 0.003
R49478 S.n14619 S.n14617 0.003
R49479 S.n14219 S.n14218 0.003
R49480 S.n13660 S.n13658 0.003
R49481 S.n13240 S.n13239 0.003
R49482 S.n12688 S.n12686 0.003
R49483 S.n12252 S.n12251 0.003
R49484 S.n11694 S.n11692 0.003
R49485 S.n11238 S.n11237 0.003
R49486 S.n10687 S.n10685 0.003
R49487 S.n10215 S.n10214 0.003
R49488 S.n9658 S.n9656 0.003
R49489 S.n7536 S.n7531 0.003
R49490 S.n8123 S.n8122 0.003
R49491 S.n22432 S.n22430 0.003
R49492 S.n22205 S.n22204 0.003
R49493 S.n21409 S.n21407 0.003
R49494 S.n21747 S.n21746 0.003
R49495 S.n20586 S.n20584 0.003
R49496 S.n20937 S.n20936 0.003
R49497 S.n19975 S.n19973 0.003
R49498 S.n19713 S.n19712 0.003
R49499 S.n19121 S.n19119 0.003
R49500 S.n18841 S.n18840 0.003
R49501 S.n18255 S.n18253 0.003
R49502 S.n17958 S.n17957 0.003
R49503 S.n17366 S.n17364 0.003
R49504 S.n17049 S.n17048 0.003
R49505 S.n16464 S.n16462 0.003
R49506 S.n16131 S.n16130 0.003
R49507 S.n15540 S.n15538 0.003
R49508 S.n15187 S.n15186 0.003
R49509 S.n14603 S.n14601 0.003
R49510 S.n14234 S.n14233 0.003
R49511 S.n13644 S.n13642 0.003
R49512 S.n13255 S.n13254 0.003
R49513 S.n12672 S.n12670 0.003
R49514 S.n12267 S.n12266 0.003
R49515 S.n11678 S.n11676 0.003
R49516 S.n11253 S.n11252 0.003
R49517 S.n10671 S.n10669 0.003
R49518 S.n10230 S.n10229 0.003
R49519 S.n9642 S.n9640 0.003
R49520 S.n9181 S.n9180 0.003
R49521 S.n8600 S.n8598 0.003
R49522 S.n6443 S.n6438 0.003
R49523 S.n7054 S.n7053 0.003
R49524 S.n22416 S.n22414 0.003
R49525 S.n22220 S.n22219 0.003
R49526 S.n21393 S.n21391 0.003
R49527 S.n21732 S.n21731 0.003
R49528 S.n20570 S.n20568 0.003
R49529 S.n20922 S.n20921 0.003
R49530 S.n19959 S.n19957 0.003
R49531 S.n19728 S.n19727 0.003
R49532 S.n19105 S.n19103 0.003
R49533 S.n18856 S.n18855 0.003
R49534 S.n18239 S.n18237 0.003
R49535 S.n17973 S.n17972 0.003
R49536 S.n17350 S.n17348 0.003
R49537 S.n17064 S.n17063 0.003
R49538 S.n16448 S.n16446 0.003
R49539 S.n16146 S.n16145 0.003
R49540 S.n15524 S.n15522 0.003
R49541 S.n15202 S.n15201 0.003
R49542 S.n14587 S.n14585 0.003
R49543 S.n14249 S.n14248 0.003
R49544 S.n13628 S.n13626 0.003
R49545 S.n13270 S.n13269 0.003
R49546 S.n12656 S.n12654 0.003
R49547 S.n12282 S.n12281 0.003
R49548 S.n11662 S.n11660 0.003
R49549 S.n11268 S.n11267 0.003
R49550 S.n10655 S.n10653 0.003
R49551 S.n10245 S.n10244 0.003
R49552 S.n9626 S.n9624 0.003
R49553 S.n9196 S.n9195 0.003
R49554 S.n8584 S.n8582 0.003
R49555 S.n8138 S.n8137 0.003
R49556 S.n7520 S.n7518 0.003
R49557 S.n5327 S.n5322 0.003
R49558 S.n5976 S.n5975 0.003
R49559 S.n22400 S.n22398 0.003
R49560 S.n22235 S.n22234 0.003
R49561 S.n21377 S.n21375 0.003
R49562 S.n21717 S.n21716 0.003
R49563 S.n20554 S.n20552 0.003
R49564 S.n20907 S.n20906 0.003
R49565 S.n19943 S.n19941 0.003
R49566 S.n19743 S.n19742 0.003
R49567 S.n19089 S.n19087 0.003
R49568 S.n18871 S.n18870 0.003
R49569 S.n18223 S.n18221 0.003
R49570 S.n17988 S.n17987 0.003
R49571 S.n17334 S.n17332 0.003
R49572 S.n17079 S.n17078 0.003
R49573 S.n16432 S.n16430 0.003
R49574 S.n16161 S.n16160 0.003
R49575 S.n15508 S.n15506 0.003
R49576 S.n15217 S.n15216 0.003
R49577 S.n14571 S.n14569 0.003
R49578 S.n14264 S.n14263 0.003
R49579 S.n13612 S.n13610 0.003
R49580 S.n13285 S.n13284 0.003
R49581 S.n12640 S.n12638 0.003
R49582 S.n12297 S.n12296 0.003
R49583 S.n11646 S.n11644 0.003
R49584 S.n11283 S.n11282 0.003
R49585 S.n10639 S.n10637 0.003
R49586 S.n10260 S.n10259 0.003
R49587 S.n9610 S.n9608 0.003
R49588 S.n9211 S.n9210 0.003
R49589 S.n8568 S.n8566 0.003
R49590 S.n8153 S.n8152 0.003
R49591 S.n7504 S.n7502 0.003
R49592 S.n7069 S.n7068 0.003
R49593 S.n6427 S.n6425 0.003
R49594 S.n4198 S.n4193 0.003
R49595 S.n4871 S.n4870 0.003
R49596 S.n22384 S.n22382 0.003
R49597 S.n22250 S.n22249 0.003
R49598 S.n21361 S.n21359 0.003
R49599 S.n21702 S.n21701 0.003
R49600 S.n20538 S.n20536 0.003
R49601 S.n20892 S.n20891 0.003
R49602 S.n19927 S.n19925 0.003
R49603 S.n19758 S.n19757 0.003
R49604 S.n19073 S.n19071 0.003
R49605 S.n18886 S.n18885 0.003
R49606 S.n18207 S.n18205 0.003
R49607 S.n18003 S.n18002 0.003
R49608 S.n17318 S.n17316 0.003
R49609 S.n17094 S.n17093 0.003
R49610 S.n16416 S.n16414 0.003
R49611 S.n16176 S.n16175 0.003
R49612 S.n15492 S.n15490 0.003
R49613 S.n15232 S.n15231 0.003
R49614 S.n14555 S.n14553 0.003
R49615 S.n14279 S.n14278 0.003
R49616 S.n13596 S.n13594 0.003
R49617 S.n13300 S.n13299 0.003
R49618 S.n12624 S.n12622 0.003
R49619 S.n12312 S.n12311 0.003
R49620 S.n11630 S.n11628 0.003
R49621 S.n11298 S.n11297 0.003
R49622 S.n10623 S.n10621 0.003
R49623 S.n10275 S.n10274 0.003
R49624 S.n9594 S.n9592 0.003
R49625 S.n9229 S.n9228 0.003
R49626 S.n8552 S.n8550 0.003
R49627 S.n8168 S.n8167 0.003
R49628 S.n7488 S.n7486 0.003
R49629 S.n7084 S.n7083 0.003
R49630 S.n6411 S.n6409 0.003
R49631 S.n5991 S.n5990 0.003
R49632 S.n5311 S.n5309 0.003
R49633 S.n3057 S.n3052 0.003
R49634 S.n3759 S.n3757 0.003
R49635 S.n22672 S.n22671 0.003
R49636 S.n22675 S.n22264 0.003
R49637 S.n21685 S.n21684 0.003
R49638 S.n21687 S.n21670 0.003
R49639 S.n20522 S.n20521 0.003
R49640 S.n20877 S.n20875 0.003
R49641 S.n19911 S.n19910 0.003
R49642 S.n19774 S.n19772 0.003
R49643 S.n19057 S.n19056 0.003
R49644 S.n18902 S.n18900 0.003
R49645 S.n18191 S.n18190 0.003
R49646 S.n18019 S.n18017 0.003
R49647 S.n17302 S.n17301 0.003
R49648 S.n17110 S.n17108 0.003
R49649 S.n16400 S.n16399 0.003
R49650 S.n16192 S.n16190 0.003
R49651 S.n15476 S.n15475 0.003
R49652 S.n15248 S.n15246 0.003
R49653 S.n14539 S.n14538 0.003
R49654 S.n14295 S.n14293 0.003
R49655 S.n13580 S.n13579 0.003
R49656 S.n13316 S.n13314 0.003
R49657 S.n12608 S.n12607 0.003
R49658 S.n12328 S.n12326 0.003
R49659 S.n11614 S.n11613 0.003
R49660 S.n11314 S.n11312 0.003
R49661 S.n10607 S.n10606 0.003
R49662 S.n10291 S.n10289 0.003
R49663 S.n9578 S.n9577 0.003
R49664 S.n9242 S.n9240 0.003
R49665 S.n8536 S.n8535 0.003
R49666 S.n8184 S.n8182 0.003
R49667 S.n7472 S.n7471 0.003
R49668 S.n7100 S.n7098 0.003
R49669 S.n6395 S.n6394 0.003
R49670 S.n6007 S.n6005 0.003
R49671 S.n5295 S.n5294 0.003
R49672 S.n4887 S.n4885 0.003
R49673 S.n4182 S.n4181 0.003
R49674 S.n1899 S.n1445 0.003
R49675 S.n2628 S.n2626 0.003
R49676 S.n22368 S.n22365 0.003
R49677 S.n22694 S.n22689 0.003
R49678 S.n21654 S.n21653 0.003
R49679 S.n21656 S.n21275 0.003
R49680 S.n20507 S.n20506 0.003
R49681 S.n20861 S.n20859 0.003
R49682 S.n19896 S.n19895 0.003
R49683 S.n19790 S.n19788 0.003
R49684 S.n19042 S.n19041 0.003
R49685 S.n18918 S.n18916 0.003
R49686 S.n18176 S.n18175 0.003
R49687 S.n18035 S.n18033 0.003
R49688 S.n17287 S.n17286 0.003
R49689 S.n17126 S.n17124 0.003
R49690 S.n16385 S.n16384 0.003
R49691 S.n16208 S.n16206 0.003
R49692 S.n15461 S.n15460 0.003
R49693 S.n15264 S.n15262 0.003
R49694 S.n14524 S.n14523 0.003
R49695 S.n14311 S.n14309 0.003
R49696 S.n13565 S.n13564 0.003
R49697 S.n13332 S.n13330 0.003
R49698 S.n12593 S.n12592 0.003
R49699 S.n12344 S.n12342 0.003
R49700 S.n11599 S.n11598 0.003
R49701 S.n11330 S.n11328 0.003
R49702 S.n10592 S.n10591 0.003
R49703 S.n10307 S.n10305 0.003
R49704 S.n9563 S.n9562 0.003
R49705 S.n9258 S.n9256 0.003
R49706 S.n8521 S.n8520 0.003
R49707 S.n8200 S.n8198 0.003
R49708 S.n7457 S.n7456 0.003
R49709 S.n7116 S.n7114 0.003
R49710 S.n6380 S.n6379 0.003
R49711 S.n6023 S.n6021 0.003
R49712 S.n5280 S.n5279 0.003
R49713 S.n4903 S.n4901 0.003
R49714 S.n4167 S.n4166 0.003
R49715 S.n3775 S.n3773 0.003
R49716 S.n3041 S.n3040 0.003
R49717 S.n914 S.n896 0.003
R49718 S.n1985 S.n1978 0.003
R49719 S.n22741 S.n22729 0.003
R49720 S.n21314 S.n21309 0.003
R49721 S.n21217 S.n21208 0.003
R49722 S.n20491 S.n20486 0.003
R49723 S.n20398 S.n20389 0.003
R49724 S.n19880 S.n19875 0.003
R49725 S.n20271 S.n20262 0.003
R49726 S.n19026 S.n19021 0.003
R49727 S.n19403 S.n19394 0.003
R49728 S.n18160 S.n18155 0.003
R49729 S.n18516 S.n18507 0.003
R49730 S.n17271 S.n17266 0.003
R49731 S.n17616 S.n17607 0.003
R49732 S.n16369 S.n16364 0.003
R49733 S.n16693 S.n16684 0.003
R49734 S.n15445 S.n15440 0.003
R49735 S.n15758 S.n15749 0.003
R49736 S.n14508 S.n14503 0.003
R49737 S.n14800 S.n14791 0.003
R49738 S.n13549 S.n13544 0.003
R49739 S.n13830 S.n13821 0.003
R49740 S.n12577 S.n12572 0.003
R49741 S.n12837 S.n12828 0.003
R49742 S.n11583 S.n11578 0.003
R49743 S.n11832 S.n11823 0.003
R49744 S.n10576 S.n10571 0.003
R49745 S.n10804 S.n10795 0.003
R49746 S.n9547 S.n9542 0.003
R49747 S.n9764 S.n9755 0.003
R49748 S.n8505 S.n8500 0.003
R49749 S.n8701 S.n8692 0.003
R49750 S.n7441 S.n7436 0.003
R49751 S.n7626 S.n7617 0.003
R49752 S.n6364 S.n6359 0.003
R49753 S.n6528 S.n6519 0.003
R49754 S.n5264 S.n5259 0.003
R49755 S.n5417 S.n5408 0.003
R49756 S.n4151 S.n4146 0.003
R49757 S.n4283 S.n4274 0.003
R49758 S.n3025 S.n3020 0.003
R49759 S.n3146 S.n3138 0.003
R49760 S.n1865 S.n1859 0.003
R49761 S.n890 S.n874 0.003
R49762 S.n806 S.n798 0.003
R49763 S.n22351 S.n22346 0.003
R49764 S.n22713 S.n22708 0.003
R49765 S.n21345 S.n21340 0.003
R49766 S.n21261 S.n21256 0.003
R49767 S.n20835 S.n20434 0.003
R49768 S.n20845 S.n20840 0.003
R49769 S.n20200 S.n19800 0.003
R49770 S.n20210 S.n20205 0.003
R49771 S.n19330 S.n18928 0.003
R49772 S.n19340 S.n19335 0.003
R49773 S.n18448 S.n18045 0.003
R49774 S.n18458 S.n18453 0.003
R49775 S.n17543 S.n17136 0.003
R49776 S.n17553 S.n17548 0.003
R49777 S.n16625 S.n16218 0.003
R49778 S.n16635 S.n16630 0.003
R49779 S.n15685 S.n15274 0.003
R49780 S.n15695 S.n15690 0.003
R49781 S.n14732 S.n14321 0.003
R49782 S.n14742 S.n14737 0.003
R49783 S.n13757 S.n13342 0.003
R49784 S.n13767 S.n13762 0.003
R49785 S.n12769 S.n12354 0.003
R49786 S.n12779 S.n12774 0.003
R49787 S.n11759 S.n11340 0.003
R49788 S.n11769 S.n11764 0.003
R49789 S.n10736 S.n10317 0.003
R49790 S.n10746 S.n10741 0.003
R49791 S.n9691 S.n9268 0.003
R49792 S.n9701 S.n9696 0.003
R49793 S.n8633 S.n8210 0.003
R49794 S.n8643 S.n8638 0.003
R49795 S.n7553 S.n7126 0.003
R49796 S.n7563 S.n7558 0.003
R49797 S.n6460 S.n6033 0.003
R49798 S.n6470 S.n6465 0.003
R49799 S.n5344 S.n4913 0.003
R49800 S.n5354 S.n5349 0.003
R49801 S.n4215 S.n3785 0.003
R49802 S.n4225 S.n4220 0.003
R49803 S.n3074 S.n2638 0.003
R49804 S.n3084 S.n3079 0.003
R49805 S.n1882 S.n1877 0.003
R49806 S.n1931 S.n1922 0.003
R49807 S.n406 S.n401 0.003
R49808 S.n2137 S.n2130 0.003
R49809 S.n18483 S.n18472 0.003
R49810 S.n17169 S.n17164 0.003
R49811 S.n17765 S.n17756 0.003
R49812 S.n16269 S.n16264 0.003
R49813 S.n16838 S.n16829 0.003
R49814 S.n15345 S.n15340 0.003
R49815 S.n15903 S.n15894 0.003
R49816 S.n14408 S.n14403 0.003
R49817 S.n14945 S.n14936 0.003
R49818 S.n13449 S.n13444 0.003
R49819 S.n13975 S.n13966 0.003
R49820 S.n12477 S.n12472 0.003
R49821 S.n12982 S.n12973 0.003
R49822 S.n11483 S.n11478 0.003
R49823 S.n11977 S.n11968 0.003
R49824 S.n10476 S.n10471 0.003
R49825 S.n10949 S.n10940 0.003
R49826 S.n9447 S.n9442 0.003
R49827 S.n9909 S.n9900 0.003
R49828 S.n8405 S.n8400 0.003
R49829 S.n8846 S.n8837 0.003
R49830 S.n7341 S.n7336 0.003
R49831 S.n7771 S.n7762 0.003
R49832 S.n6264 S.n6259 0.003
R49833 S.n6673 S.n6664 0.003
R49834 S.n5164 S.n5159 0.003
R49835 S.n5563 S.n5554 0.003
R49836 S.n4052 S.n4047 0.003
R49837 S.n4428 S.n4419 0.003
R49838 S.n2925 S.n2920 0.003
R49839 S.n3290 S.n3282 0.003
R49840 S.n1757 S.n1751 0.003
R49841 S.n24 S.n13 0.003
R49842 S.n19370 S.n19358 0.003
R49843 S.n18077 S.n18072 0.003
R49844 S.n18633 S.n18619 0.003
R49845 S.n17188 S.n17183 0.003
R49846 S.n17733 S.n17719 0.003
R49847 S.n16286 S.n16281 0.003
R49848 S.n16806 S.n16792 0.003
R49849 S.n15362 S.n15357 0.003
R49850 S.n15871 S.n15857 0.003
R49851 S.n14425 S.n14420 0.003
R49852 S.n14913 S.n14899 0.003
R49853 S.n13466 S.n13461 0.003
R49854 S.n13943 S.n13929 0.003
R49855 S.n12494 S.n12489 0.003
R49856 S.n12950 S.n12936 0.003
R49857 S.n11500 S.n11495 0.003
R49858 S.n11945 S.n11931 0.003
R49859 S.n10493 S.n10488 0.003
R49860 S.n10917 S.n10903 0.003
R49861 S.n9464 S.n9459 0.003
R49862 S.n9877 S.n9863 0.003
R49863 S.n8422 S.n8417 0.003
R49864 S.n8814 S.n8800 0.003
R49865 S.n7358 S.n7353 0.003
R49866 S.n7739 S.n7725 0.003
R49867 S.n6281 S.n6276 0.003
R49868 S.n6641 S.n6627 0.003
R49869 S.n5181 S.n5176 0.003
R49870 S.n5531 S.n5517 0.003
R49871 S.n4069 S.n4064 0.003
R49872 S.n4396 S.n4382 0.003
R49873 S.n2942 S.n2937 0.003
R49874 S.n3259 S.n3245 0.003
R49875 S.n1776 S.n1769 0.003
R49876 S.n1799 S.n1791 0.003
R49877 S.n2079 S.n2061 0.003
R49878 S.n823 S.n416 0.003
R49879 S.n838 S.n829 0.003
R49880 S.n3230 S.n3222 0.003
R49881 S.n4367 S.n4358 0.003
R49882 S.n5502 S.n5493 0.003
R49883 S.n6612 S.n6603 0.003
R49884 S.n7710 S.n7701 0.003
R49885 S.n8785 S.n8776 0.003
R49886 S.n9848 S.n9839 0.003
R49887 S.n10888 S.n10879 0.003
R49888 S.n11916 S.n11907 0.003
R49889 S.n12921 S.n12912 0.003
R49890 S.n13914 S.n13905 0.003
R49891 S.n14884 S.n14875 0.003
R49892 S.n15842 S.n15833 0.003
R49893 S.n16777 S.n16768 0.003
R49894 S.n17700 S.n17691 0.003
R49895 S.n18600 S.n18591 0.003
R49896 S.n19490 S.n19481 0.003
R49897 S.n20238 S.n20227 0.003
R49898 S.n18961 S.n18956 0.003
R49899 S.n18096 S.n18091 0.003
R49900 S.n17207 S.n17202 0.003
R49901 S.n16305 S.n16300 0.003
R49902 S.n15381 S.n15376 0.003
R49903 S.n14444 S.n14439 0.003
R49904 S.n13485 S.n13480 0.003
R49905 S.n12513 S.n12508 0.003
R49906 S.n11519 S.n11514 0.003
R49907 S.n10512 S.n10507 0.003
R49908 S.n9483 S.n9478 0.003
R49909 S.n8441 S.n8436 0.003
R49910 S.n7377 S.n7372 0.003
R49911 S.n6300 S.n6295 0.003
R49912 S.n5200 S.n5195 0.003
R49913 S.n4088 S.n4083 0.003
R49914 S.n2961 S.n2956 0.003
R49915 S.n2045 S.n2033 0.003
R49916 S.n767 S.n754 0.003
R49917 S.n1337 S.n1325 0.003
R49918 S.n20424 S.n20419 0.003
R49919 S.n19839 S.n19836 0.003
R49920 S.n20330 S.n20315 0.003
R49921 S.n18987 S.n18984 0.003
R49922 S.n19458 S.n19443 0.003
R49923 S.n18121 S.n18119 0.003
R49924 S.n18568 S.n18556 0.003
R49925 S.n17232 S.n17230 0.003
R49926 S.n17668 S.n17656 0.003
R49927 S.n16330 S.n16328 0.003
R49928 S.n16745 S.n16733 0.003
R49929 S.n15406 S.n15404 0.003
R49930 S.n15810 S.n15798 0.003
R49931 S.n14469 S.n14467 0.003
R49932 S.n14852 S.n14840 0.003
R49933 S.n13510 S.n13508 0.003
R49934 S.n13882 S.n13870 0.003
R49935 S.n12538 S.n12536 0.003
R49936 S.n12889 S.n12877 0.003
R49937 S.n11544 S.n11542 0.003
R49938 S.n11884 S.n11872 0.003
R49939 S.n10537 S.n10535 0.003
R49940 S.n10856 S.n10844 0.003
R49941 S.n9508 S.n9506 0.003
R49942 S.n9816 S.n9804 0.003
R49943 S.n8466 S.n8464 0.003
R49944 S.n8753 S.n8741 0.003
R49945 S.n7402 S.n7400 0.003
R49946 S.n7678 S.n7666 0.003
R49947 S.n6325 S.n6323 0.003
R49948 S.n6580 S.n6568 0.003
R49949 S.n5225 S.n5223 0.003
R49950 S.n5470 S.n5458 0.003
R49951 S.n4113 S.n4111 0.003
R49952 S.n4335 S.n4323 0.003
R49953 S.n2986 S.n2984 0.003
R49954 S.n3198 S.n3186 0.003
R49955 S.n1823 S.n1821 0.003
R49956 S.n2012 S.n2000 0.003
R49957 S.n786 S.n778 0.003
R49958 S.n1845 S.n1842 0.003
R49959 S.n3166 S.n3161 0.003
R49960 S.n3006 S.n2998 0.003
R49961 S.n4303 S.n4298 0.003
R49962 S.n4132 S.n4125 0.003
R49963 S.n5438 S.n5432 0.003
R49964 S.n5245 S.n5237 0.003
R49965 S.n6548 S.n6543 0.003
R49966 S.n6345 S.n6337 0.003
R49967 S.n7646 S.n7641 0.003
R49968 S.n7422 S.n7414 0.003
R49969 S.n8721 S.n8716 0.003
R49970 S.n8486 S.n8478 0.003
R49971 S.n9784 S.n9779 0.003
R49972 S.n9528 S.n9520 0.003
R49973 S.n10824 S.n10819 0.003
R49974 S.n10557 S.n10549 0.003
R49975 S.n11852 S.n11847 0.003
R49976 S.n11564 S.n11556 0.003
R49977 S.n12857 S.n12852 0.003
R49978 S.n12558 S.n12550 0.003
R49979 S.n13850 S.n13845 0.003
R49980 S.n13530 S.n13522 0.003
R49981 S.n14820 S.n14815 0.003
R49982 S.n14489 S.n14481 0.003
R49983 S.n15778 S.n15773 0.003
R49984 S.n15426 S.n15418 0.003
R49985 S.n16713 S.n16708 0.003
R49986 S.n16350 S.n16342 0.003
R49987 S.n17636 S.n17631 0.003
R49988 S.n17252 S.n17244 0.003
R49989 S.n18536 S.n18531 0.003
R49990 S.n18141 S.n18133 0.003
R49991 S.n19423 S.n19418 0.003
R49992 S.n19007 S.n18999 0.003
R49993 S.n20295 S.n20290 0.003
R49994 S.n19861 S.n19853 0.003
R49995 S.n20366 S.n20361 0.003
R49996 S.n20472 S.n20464 0.003
R49997 S.n21242 S.n21237 0.003
R49998 S.n864 S.n853 0.003
R49999 S.n2107 S.n2094 0.003
R50000 S.n743 S.n738 0.003
R50001 S.n726 S.n721 0.003
R50002 S.n374 S.n369 0.003
R50003 S.n2196 S.n2189 0.003
R50004 S.n16660 S.n16649 0.003
R50005 S.n15307 S.n15302 0.003
R50006 S.n15968 S.n15959 0.003
R50007 S.n14372 S.n14367 0.003
R50008 S.n15006 S.n14997 0.003
R50009 S.n13413 S.n13408 0.003
R50010 S.n14036 S.n14027 0.003
R50011 S.n12441 S.n12436 0.003
R50012 S.n13043 S.n13034 0.003
R50013 S.n11447 S.n11442 0.003
R50014 S.n12038 S.n12029 0.003
R50015 S.n10440 S.n10435 0.003
R50016 S.n11010 S.n11001 0.003
R50017 S.n9411 S.n9406 0.003
R50018 S.n9970 S.n9961 0.003
R50019 S.n8369 S.n8364 0.003
R50020 S.n8907 S.n8898 0.003
R50021 S.n7305 S.n7300 0.003
R50022 S.n7832 S.n7823 0.003
R50023 S.n6228 S.n6223 0.003
R50024 S.n6734 S.n6725 0.003
R50025 S.n5128 S.n5123 0.003
R50026 S.n5624 S.n5615 0.003
R50027 S.n4016 S.n4011 0.003
R50028 S.n4489 S.n4480 0.003
R50029 S.n2889 S.n2884 0.003
R50030 S.n3350 S.n3342 0.003
R50031 S.n1720 S.n1714 0.003
R50032 S.n71 S.n60 0.003
R50033 S.n17583 S.n17571 0.003
R50034 S.n16250 S.n16245 0.003
R50035 S.n16871 S.n16857 0.003
R50036 S.n15326 S.n15321 0.003
R50037 S.n15936 S.n15922 0.003
R50038 S.n14389 S.n14384 0.003
R50039 S.n14974 S.n14960 0.003
R50040 S.n13430 S.n13425 0.003
R50041 S.n14004 S.n13990 0.003
R50042 S.n12458 S.n12453 0.003
R50043 S.n13011 S.n12997 0.003
R50044 S.n11464 S.n11459 0.003
R50045 S.n12006 S.n11992 0.003
R50046 S.n10457 S.n10452 0.003
R50047 S.n10978 S.n10964 0.003
R50048 S.n9428 S.n9423 0.003
R50049 S.n9938 S.n9924 0.003
R50050 S.n8386 S.n8381 0.003
R50051 S.n8875 S.n8861 0.003
R50052 S.n7322 S.n7317 0.003
R50053 S.n7800 S.n7786 0.003
R50054 S.n6245 S.n6240 0.003
R50055 S.n6702 S.n6688 0.003
R50056 S.n5145 S.n5140 0.003
R50057 S.n5592 S.n5578 0.003
R50058 S.n4033 S.n4028 0.003
R50059 S.n4457 S.n4443 0.003
R50060 S.n2906 S.n2901 0.003
R50061 S.n3319 S.n3305 0.003
R50062 S.n1737 S.n1732 0.003
R50063 S.n2166 S.n2152 0.003
R50064 S.n708 S.n703 0.003
R50065 S.n691 S.n686 0.003
R50066 S.n342 S.n337 0.003
R50067 S.n2255 S.n2248 0.003
R50068 S.n14767 S.n14756 0.003
R50069 S.n13375 S.n13370 0.003
R50070 S.n14101 S.n14092 0.003
R50071 S.n12405 S.n12400 0.003
R50072 S.n13104 S.n13095 0.003
R50073 S.n11411 S.n11406 0.003
R50074 S.n12099 S.n12090 0.003
R50075 S.n10404 S.n10399 0.003
R50076 S.n11071 S.n11062 0.003
R50077 S.n9375 S.n9370 0.003
R50078 S.n10031 S.n10022 0.003
R50079 S.n8333 S.n8328 0.003
R50080 S.n8968 S.n8959 0.003
R50081 S.n7269 S.n7264 0.003
R50082 S.n7893 S.n7884 0.003
R50083 S.n6192 S.n6187 0.003
R50084 S.n6795 S.n6786 0.003
R50085 S.n5092 S.n5087 0.003
R50086 S.n5685 S.n5676 0.003
R50087 S.n3980 S.n3975 0.003
R50088 S.n4550 S.n4541 0.003
R50089 S.n2853 S.n2848 0.003
R50090 S.n3410 S.n3402 0.003
R50091 S.n1683 S.n1677 0.003
R50092 S.n103 S.n92 0.003
R50093 S.n15725 S.n15713 0.003
R50094 S.n14353 S.n14348 0.003
R50095 S.n15039 S.n15025 0.003
R50096 S.n13394 S.n13389 0.003
R50097 S.n14069 S.n14055 0.003
R50098 S.n12422 S.n12417 0.003
R50099 S.n13072 S.n13058 0.003
R50100 S.n11428 S.n11423 0.003
R50101 S.n12067 S.n12053 0.003
R50102 S.n10421 S.n10416 0.003
R50103 S.n11039 S.n11025 0.003
R50104 S.n9392 S.n9387 0.003
R50105 S.n9999 S.n9985 0.003
R50106 S.n8350 S.n8345 0.003
R50107 S.n8936 S.n8922 0.003
R50108 S.n7286 S.n7281 0.003
R50109 S.n7861 S.n7847 0.003
R50110 S.n6209 S.n6204 0.003
R50111 S.n6763 S.n6749 0.003
R50112 S.n5109 S.n5104 0.003
R50113 S.n5653 S.n5639 0.003
R50114 S.n3997 S.n3992 0.003
R50115 S.n4518 S.n4504 0.003
R50116 S.n2870 S.n2865 0.003
R50117 S.n3379 S.n3365 0.003
R50118 S.n1700 S.n1695 0.003
R50119 S.n2225 S.n2211 0.003
R50120 S.n673 S.n668 0.003
R50121 S.n656 S.n651 0.003
R50122 S.n310 S.n305 0.003
R50123 S.n2314 S.n2307 0.003
R50124 S.n12804 S.n12793 0.003
R50125 S.n11373 S.n11368 0.003
R50126 S.n12164 S.n12155 0.003
R50127 S.n10368 S.n10363 0.003
R50128 S.n11132 S.n11123 0.003
R50129 S.n9339 S.n9334 0.003
R50130 S.n10092 S.n10083 0.003
R50131 S.n8297 S.n8292 0.003
R50132 S.n9029 S.n9020 0.003
R50133 S.n7233 S.n7228 0.003
R50134 S.n7954 S.n7945 0.003
R50135 S.n6156 S.n6151 0.003
R50136 S.n6856 S.n6847 0.003
R50137 S.n5056 S.n5051 0.003
R50138 S.n5746 S.n5737 0.003
R50139 S.n3944 S.n3939 0.003
R50140 S.n4611 S.n4602 0.003
R50141 S.n2817 S.n2812 0.003
R50142 S.n3470 S.n3462 0.003
R50143 S.n1646 S.n1640 0.003
R50144 S.n990 S.n124 0.003
R50145 S.n13797 S.n13785 0.003
R50146 S.n12386 S.n12381 0.003
R50147 S.n13137 S.n13123 0.003
R50148 S.n11392 S.n11387 0.003
R50149 S.n12132 S.n12118 0.003
R50150 S.n10385 S.n10380 0.003
R50151 S.n11100 S.n11086 0.003
R50152 S.n9356 S.n9351 0.003
R50153 S.n10060 S.n10046 0.003
R50154 S.n8314 S.n8309 0.003
R50155 S.n8997 S.n8983 0.003
R50156 S.n7250 S.n7245 0.003
R50157 S.n7922 S.n7908 0.003
R50158 S.n6173 S.n6168 0.003
R50159 S.n6824 S.n6810 0.003
R50160 S.n5073 S.n5068 0.003
R50161 S.n5714 S.n5700 0.003
R50162 S.n3961 S.n3956 0.003
R50163 S.n4579 S.n4565 0.003
R50164 S.n2834 S.n2829 0.003
R50165 S.n3439 S.n3425 0.003
R50166 S.n1663 S.n1658 0.003
R50167 S.n2284 S.n2270 0.003
R50168 S.n638 S.n633 0.003
R50169 S.n621 S.n616 0.003
R50170 S.n278 S.n273 0.003
R50171 S.n2373 S.n2366 0.003
R50172 S.n10771 S.n10760 0.003
R50173 S.n9301 S.n9296 0.003
R50174 S.n10157 S.n10148 0.003
R50175 S.n8261 S.n8256 0.003
R50176 S.n9090 S.n9081 0.003
R50177 S.n7197 S.n7192 0.003
R50178 S.n8015 S.n8006 0.003
R50179 S.n6120 S.n6115 0.003
R50180 S.n6917 S.n6908 0.003
R50181 S.n5020 S.n5015 0.003
R50182 S.n5807 S.n5798 0.003
R50183 S.n3908 S.n3903 0.003
R50184 S.n4672 S.n4663 0.003
R50185 S.n2781 S.n2776 0.003
R50186 S.n3530 S.n3522 0.003
R50187 S.n1609 S.n1603 0.003
R50188 S.n1022 S.n1011 0.003
R50189 S.n11799 S.n11787 0.003
R50190 S.n10349 S.n10344 0.003
R50191 S.n11165 S.n11151 0.003
R50192 S.n9320 S.n9315 0.003
R50193 S.n10125 S.n10111 0.003
R50194 S.n8278 S.n8273 0.003
R50195 S.n9058 S.n9044 0.003
R50196 S.n7214 S.n7209 0.003
R50197 S.n7983 S.n7969 0.003
R50198 S.n6137 S.n6132 0.003
R50199 S.n6885 S.n6871 0.003
R50200 S.n5037 S.n5032 0.003
R50201 S.n5775 S.n5761 0.003
R50202 S.n3925 S.n3920 0.003
R50203 S.n4640 S.n4626 0.003
R50204 S.n2798 S.n2793 0.003
R50205 S.n3499 S.n3485 0.003
R50206 S.n1626 S.n1621 0.003
R50207 S.n2343 S.n2329 0.003
R50208 S.n603 S.n598 0.003
R50209 S.n586 S.n581 0.003
R50210 S.n249 S.n244 0.003
R50211 S.n2432 S.n2425 0.003
R50212 S.n8668 S.n8657 0.003
R50213 S.n7159 S.n7154 0.003
R50214 S.n8080 S.n8071 0.003
R50215 S.n6084 S.n6079 0.003
R50216 S.n6978 S.n6969 0.003
R50217 S.n4984 S.n4979 0.003
R50218 S.n5868 S.n5859 0.003
R50219 S.n3872 S.n3867 0.003
R50220 S.n4733 S.n4724 0.003
R50221 S.n2745 S.n2740 0.003
R50222 S.n3590 S.n3582 0.003
R50223 S.n1572 S.n1566 0.003
R50224 S.n1054 S.n1043 0.003
R50225 S.n9731 S.n9719 0.003
R50226 S.n8242 S.n8237 0.003
R50227 S.n9123 S.n9109 0.003
R50228 S.n7178 S.n7173 0.003
R50229 S.n8048 S.n8034 0.003
R50230 S.n6101 S.n6096 0.003
R50231 S.n6946 S.n6932 0.003
R50232 S.n5001 S.n4996 0.003
R50233 S.n5836 S.n5822 0.003
R50234 S.n3889 S.n3884 0.003
R50235 S.n4701 S.n4687 0.003
R50236 S.n2762 S.n2757 0.003
R50237 S.n3559 S.n3545 0.003
R50238 S.n1589 S.n1584 0.003
R50239 S.n2402 S.n2388 0.003
R50240 S.n568 S.n563 0.003
R50241 S.n551 S.n546 0.003
R50242 S.n214 S.n209 0.003
R50243 S.n2491 S.n2484 0.003
R50244 S.n6495 S.n6484 0.003
R50245 S.n4946 S.n4941 0.003
R50246 S.n5933 S.n5924 0.003
R50247 S.n3836 S.n3831 0.003
R50248 S.n4794 S.n4785 0.003
R50249 S.n2709 S.n2704 0.003
R50250 S.n3650 S.n3642 0.003
R50251 S.n1535 S.n1529 0.003
R50252 S.n1086 S.n1075 0.003
R50253 S.n7593 S.n7581 0.003
R50254 S.n6065 S.n6060 0.003
R50255 S.n7011 S.n6997 0.003
R50256 S.n4965 S.n4960 0.003
R50257 S.n5901 S.n5887 0.003
R50258 S.n3853 S.n3848 0.003
R50259 S.n4762 S.n4748 0.003
R50260 S.n2726 S.n2721 0.003
R50261 S.n3619 S.n3605 0.003
R50262 S.n1552 S.n1547 0.003
R50263 S.n2461 S.n2447 0.003
R50264 S.n533 S.n528 0.003
R50265 S.n516 S.n511 0.003
R50266 S.n182 S.n177 0.003
R50267 S.n2550 S.n2543 0.003
R50268 S.n4250 S.n4239 0.003
R50269 S.n2671 S.n2666 0.003
R50270 S.n3714 S.n3706 0.003
R50271 S.n1498 S.n1492 0.003
R50272 S.n1118 S.n1107 0.003
R50273 S.n5384 S.n5372 0.003
R50274 S.n3817 S.n3812 0.003
R50275 S.n4827 S.n4813 0.003
R50276 S.n2690 S.n2685 0.003
R50277 S.n3683 S.n3669 0.003
R50278 S.n1515 S.n1510 0.003
R50279 S.n2520 S.n2506 0.003
R50280 S.n498 S.n493 0.003
R50281 S.n481 S.n476 0.003
R50282 S.n150 S.n145 0.003
R50283 S.n1954 S.n1945 0.003
R50284 S.n1156 S.n1145 0.003
R50285 S.n3114 S.n3102 0.003
R50286 S.n1478 S.n1473 0.003
R50287 S.n2583 S.n2569 0.003
R50288 S.n463 S.n458 0.003
R50289 S.n447 S.n442 0.003
R50290 S.n942 S.n932 0.003
R50291 S.n22765 S.n22760 0.003
R50292 S.n21328 S.n21323 0.003
R50293 S.n1373 S.n1371 0.003
R50294 S.n4 S.n2 0.003
R50295 S.n51 S.n49 0.003
R50296 S.n82 S.n80 0.003
R50297 S.n114 S.n112 0.003
R50298 S.n1001 S.n999 0.003
R50299 S.n1033 S.n1031 0.003
R50300 S.n1065 S.n1063 0.003
R50301 S.n1097 S.n1095 0.003
R50302 S.n1129 S.n1127 0.003
R50303 S.n1167 S.n1165 0.003
R50304 S.n23010 S.n23009 0.003
R50305 S.n23010 S.n22804 0.003
R50306 S.n20451 S.n20450 0.003
R50307 S.n1357 S.n1356 0.003
R50308 S.n850 S.n849 0.003
R50309 S.n10 S.n9 0.003
R50310 S.n57 S.n56 0.003
R50311 S.n89 S.n88 0.003
R50312 S.n121 S.n120 0.003
R50313 S.n1008 S.n1007 0.003
R50314 S.n1040 S.n1039 0.003
R50315 S.n1072 S.n1071 0.003
R50316 S.n1104 S.n1103 0.003
R50317 S.n1142 S.n1141 0.003
R50318 S.n21152 S.n21147 0.003
R50319 S.n836 S.n835 0.003
R50320 S.n20439 S.n20438 0.003
R50321 S.n18568 S.n18567 0.003
R50322 S.n17668 S.n17667 0.003
R50323 S.n16745 S.n16744 0.003
R50324 S.n15810 S.n15809 0.003
R50325 S.n14852 S.n14851 0.003
R50326 S.n13882 S.n13881 0.003
R50327 S.n12889 S.n12888 0.003
R50328 S.n11884 S.n11883 0.003
R50329 S.n10856 S.n10855 0.003
R50330 S.n9816 S.n9815 0.003
R50331 S.n8753 S.n8752 0.003
R50332 S.n7678 S.n7677 0.003
R50333 S.n6580 S.n6579 0.003
R50334 S.n5470 S.n5469 0.003
R50335 S.n4335 S.n4334 0.003
R50336 S.n3198 S.n3197 0.003
R50337 S.n2045 S.n2029 0.003
R50338 S.n397 S.n396 0.003
R50339 S.n365 S.n364 0.003
R50340 S.n333 S.n332 0.003
R50341 S.n301 S.n300 0.003
R50342 S.n269 S.n268 0.003
R50343 S.n240 S.n239 0.003
R50344 S.n205 S.n204 0.003
R50345 S.n173 S.n172 0.003
R50346 S.n1138 S.n1133 0.003
R50347 S.n1138 S.n1137 0.003
R50348 S.n141 S.n140 0.003
R50349 S.n20344 S.n19520 0.003
R50350 S.n19504 S.n18663 0.003
R50351 S.n18647 S.n17795 0.003
R50352 S.n17779 S.n16901 0.003
R50353 S.n16885 S.n15998 0.003
R50354 S.n15982 S.n15069 0.003
R50355 S.n15053 S.n14131 0.003
R50356 S.n14115 S.n13167 0.003
R50357 S.n13151 S.n12194 0.003
R50358 S.n12178 S.n11195 0.003
R50359 S.n11179 S.n10187 0.003
R50360 S.n10171 S.n9153 0.003
R50361 S.n9137 S.n8110 0.003
R50362 S.n8094 S.n7041 0.003
R50363 S.n7025 S.n5963 0.003
R50364 S.n5947 S.n4858 0.003
R50365 S.t41 S.n22997 0.003
R50366 S.n974 S.n973 0.003
R50367 S.n22288 S.n22271 0.003
R50368 S.n18059 S.n18058 0.003
R50369 S.n16232 S.n16231 0.003
R50370 S.n14335 S.n14334 0.003
R50371 S.n12368 S.n12367 0.003
R50372 S.n10331 S.n10330 0.003
R50373 S.n8224 S.n8223 0.003
R50374 S.n6047 S.n6046 0.003
R50375 S.n3799 S.n3798 0.003
R50376 S.n1460 S.n1459 0.003
R50377 S.n21133 S.n21126 0.003
R50378 S.t41 S.n22807 0.003
R50379 S.t41 S.n22982 0.003
R50380 S.n21233 S.n21232 0.003
R50381 S.n20357 S.n20356 0.003
R50382 S.n20286 S.n20285 0.003
R50383 S.n4841 S.n3745 0.003
R50384 S.n3728 S.n2614 0.003
R50385 S.n18077 S.n18068 0.003
R50386 S.n17188 S.n17179 0.003
R50387 S.n16286 S.n16277 0.003
R50388 S.n15362 S.n15353 0.003
R50389 S.n14425 S.n14416 0.003
R50390 S.n13466 S.n13457 0.003
R50391 S.n12494 S.n12485 0.003
R50392 S.n11500 S.n11491 0.003
R50393 S.n10493 S.n10484 0.003
R50394 S.n9464 S.n9455 0.003
R50395 S.n8422 S.n8413 0.003
R50396 S.n7358 S.n7349 0.003
R50397 S.n6281 S.n6272 0.003
R50398 S.n5181 S.n5172 0.003
R50399 S.n4069 S.n4060 0.003
R50400 S.n2942 S.n2933 0.003
R50401 S.n1776 S.n1765 0.003
R50402 S.n16250 S.n16241 0.003
R50403 S.n15326 S.n15317 0.003
R50404 S.n14389 S.n14380 0.003
R50405 S.n13430 S.n13421 0.003
R50406 S.n12458 S.n12449 0.003
R50407 S.n11464 S.n11455 0.003
R50408 S.n10457 S.n10448 0.003
R50409 S.n9428 S.n9419 0.003
R50410 S.n8386 S.n8377 0.003
R50411 S.n7322 S.n7313 0.003
R50412 S.n6245 S.n6236 0.003
R50413 S.n5145 S.n5136 0.003
R50414 S.n4033 S.n4024 0.003
R50415 S.n2906 S.n2897 0.003
R50416 S.n1737 S.n1728 0.003
R50417 S.n14353 S.n14344 0.003
R50418 S.n13394 S.n13385 0.003
R50419 S.n12422 S.n12413 0.003
R50420 S.n11428 S.n11419 0.003
R50421 S.n10421 S.n10412 0.003
R50422 S.n9392 S.n9383 0.003
R50423 S.n8350 S.n8341 0.003
R50424 S.n7286 S.n7277 0.003
R50425 S.n6209 S.n6200 0.003
R50426 S.n5109 S.n5100 0.003
R50427 S.n3997 S.n3988 0.003
R50428 S.n2870 S.n2861 0.003
R50429 S.n1700 S.n1691 0.003
R50430 S.n12386 S.n12377 0.003
R50431 S.n11392 S.n11383 0.003
R50432 S.n10385 S.n10376 0.003
R50433 S.n9356 S.n9347 0.003
R50434 S.n8314 S.n8305 0.003
R50435 S.n7250 S.n7241 0.003
R50436 S.n6173 S.n6164 0.003
R50437 S.n5073 S.n5064 0.003
R50438 S.n3961 S.n3952 0.003
R50439 S.n2834 S.n2825 0.003
R50440 S.n1663 S.n1654 0.003
R50441 S.n10349 S.n10340 0.003
R50442 S.n9320 S.n9311 0.003
R50443 S.n8278 S.n8269 0.003
R50444 S.n7214 S.n7205 0.003
R50445 S.n6137 S.n6128 0.003
R50446 S.n5037 S.n5028 0.003
R50447 S.n3925 S.n3916 0.003
R50448 S.n2798 S.n2789 0.003
R50449 S.n1626 S.n1617 0.003
R50450 S.n8242 S.n8233 0.003
R50451 S.n7178 S.n7169 0.003
R50452 S.n6101 S.n6092 0.003
R50453 S.n5001 S.n4992 0.003
R50454 S.n3889 S.n3880 0.003
R50455 S.n2762 S.n2753 0.003
R50456 S.n1589 S.n1580 0.003
R50457 S.n6065 S.n6056 0.003
R50458 S.n4965 S.n4956 0.003
R50459 S.n3853 S.n3844 0.003
R50460 S.n2726 S.n2717 0.003
R50461 S.n1552 S.n1543 0.003
R50462 S.n3817 S.n3808 0.003
R50463 S.n2690 S.n2681 0.003
R50464 S.n1515 S.n1506 0.003
R50465 S.n1478 S.n1469 0.003
R50466 S.n22791 S.n22790 0.003
R50467 S.n890 S.n889 0.003
R50468 S.n2547 S.n2546 0.003
R50469 S.n1948 S.n1947 0.003
R50470 S.n20325 S.n20324 0.003
R50471 S.n19453 S.n19452 0.003
R50472 S.n1350 S.n1349 0.003
R50473 S.n20818 S.n20807 0.002
R50474 S.n21962 S.n21953 0.002
R50475 S.n21638 S.n21630 0.002
R50476 S.n21995 S.n21987 0.002
R50477 S.n22656 S.n22648 0.002
R50478 S.n22640 S.n22631 0.002
R50479 S.n22010 S.n22002 0.002
R50480 S.n21617 S.n21608 0.002
R50481 S.n21942 S.n21934 0.002
R50482 S.n20794 S.n20785 0.002
R50483 S.n21133 S.n21124 0.002
R50484 S.n20183 S.n20175 0.002
R50485 S.n22624 S.n22615 0.002
R50486 S.n22025 S.n22017 0.002
R50487 S.n21601 S.n21592 0.002
R50488 S.n21927 S.n21919 0.002
R50489 S.n20778 S.n20769 0.002
R50490 S.n21117 S.n21109 0.002
R50491 S.n20167 S.n20158 0.002
R50492 S.n19533 S.n19525 0.002
R50493 S.n19313 S.n19305 0.002
R50494 S.n22608 S.n22599 0.002
R50495 S.n22040 S.n22032 0.002
R50496 S.n21585 S.n21576 0.002
R50497 S.n21912 S.n21904 0.002
R50498 S.n20762 S.n20753 0.002
R50499 S.n21102 S.n21094 0.002
R50500 S.n20151 S.n20142 0.002
R50501 S.n19548 S.n19540 0.002
R50502 S.n19297 S.n19288 0.002
R50503 S.n18676 S.n18668 0.002
R50504 S.n18431 S.n18423 0.002
R50505 S.n22592 S.n22583 0.002
R50506 S.n22055 S.n22047 0.002
R50507 S.n21569 S.n21560 0.002
R50508 S.n21897 S.n21889 0.002
R50509 S.n20746 S.n20737 0.002
R50510 S.n21087 S.n21079 0.002
R50511 S.n20135 S.n20126 0.002
R50512 S.n19563 S.n19555 0.002
R50513 S.n19281 S.n19272 0.002
R50514 S.n18691 S.n18683 0.002
R50515 S.n18415 S.n18406 0.002
R50516 S.n17808 S.n17800 0.002
R50517 S.n17526 S.n17518 0.002
R50518 S.n22576 S.n22567 0.002
R50519 S.n22070 S.n22062 0.002
R50520 S.n21553 S.n21544 0.002
R50521 S.n21882 S.n21874 0.002
R50522 S.n20730 S.n20721 0.002
R50523 S.n21072 S.n21064 0.002
R50524 S.n20119 S.n20110 0.002
R50525 S.n19578 S.n19570 0.002
R50526 S.n19265 S.n19256 0.002
R50527 S.n18706 S.n18698 0.002
R50528 S.n18399 S.n18390 0.002
R50529 S.n17823 S.n17815 0.002
R50530 S.n17510 S.n17501 0.002
R50531 S.n16914 S.n16906 0.002
R50532 S.n16608 S.n16600 0.002
R50533 S.n22560 S.n22551 0.002
R50534 S.n22085 S.n22077 0.002
R50535 S.n21537 S.n21528 0.002
R50536 S.n21867 S.n21859 0.002
R50537 S.n20714 S.n20705 0.002
R50538 S.n21057 S.n21049 0.002
R50539 S.n20103 S.n20094 0.002
R50540 S.n19593 S.n19585 0.002
R50541 S.n19249 S.n19240 0.002
R50542 S.n18721 S.n18713 0.002
R50543 S.n18383 S.n18374 0.002
R50544 S.n17838 S.n17830 0.002
R50545 S.n17494 S.n17485 0.002
R50546 S.n16929 S.n16921 0.002
R50547 S.n16592 S.n16583 0.002
R50548 S.n16011 S.n16003 0.002
R50549 S.n15668 S.n15660 0.002
R50550 S.n22544 S.n22535 0.002
R50551 S.n22100 S.n22092 0.002
R50552 S.n21521 S.n21512 0.002
R50553 S.n21852 S.n21844 0.002
R50554 S.n20698 S.n20689 0.002
R50555 S.n21042 S.n21034 0.002
R50556 S.n20087 S.n20078 0.002
R50557 S.n19608 S.n19600 0.002
R50558 S.n19233 S.n19224 0.002
R50559 S.n18736 S.n18728 0.002
R50560 S.n18367 S.n18358 0.002
R50561 S.n17853 S.n17845 0.002
R50562 S.n17478 S.n17469 0.002
R50563 S.n16944 S.n16936 0.002
R50564 S.n16576 S.n16567 0.002
R50565 S.n16026 S.n16018 0.002
R50566 S.n15652 S.n15643 0.002
R50567 S.n15082 S.n15074 0.002
R50568 S.n14715 S.n14707 0.002
R50569 S.n22528 S.n22519 0.002
R50570 S.n22115 S.n22107 0.002
R50571 S.n21505 S.n21496 0.002
R50572 S.n21837 S.n21829 0.002
R50573 S.n20682 S.n20673 0.002
R50574 S.n21027 S.n21019 0.002
R50575 S.n20071 S.n20062 0.002
R50576 S.n19623 S.n19615 0.002
R50577 S.n19217 S.n19208 0.002
R50578 S.n18751 S.n18743 0.002
R50579 S.n18351 S.n18342 0.002
R50580 S.n17868 S.n17860 0.002
R50581 S.n17462 S.n17453 0.002
R50582 S.n16959 S.n16951 0.002
R50583 S.n16560 S.n16551 0.002
R50584 S.n16041 S.n16033 0.002
R50585 S.n15636 S.n15627 0.002
R50586 S.n15097 S.n15089 0.002
R50587 S.n14699 S.n14690 0.002
R50588 S.n14144 S.n14136 0.002
R50589 S.n13740 S.n13732 0.002
R50590 S.n22512 S.n22503 0.002
R50591 S.n22130 S.n22122 0.002
R50592 S.n21489 S.n21480 0.002
R50593 S.n21822 S.n21814 0.002
R50594 S.n20666 S.n20657 0.002
R50595 S.n21012 S.n21004 0.002
R50596 S.n20055 S.n20046 0.002
R50597 S.n19638 S.n19630 0.002
R50598 S.n19201 S.n19192 0.002
R50599 S.n18766 S.n18758 0.002
R50600 S.n18335 S.n18326 0.002
R50601 S.n17883 S.n17875 0.002
R50602 S.n17446 S.n17437 0.002
R50603 S.n16974 S.n16966 0.002
R50604 S.n16544 S.n16535 0.002
R50605 S.n16056 S.n16048 0.002
R50606 S.n15620 S.n15611 0.002
R50607 S.n15112 S.n15104 0.002
R50608 S.n14683 S.n14674 0.002
R50609 S.n14159 S.n14151 0.002
R50610 S.n13724 S.n13715 0.002
R50611 S.n13180 S.n13172 0.002
R50612 S.n12752 S.n12744 0.002
R50613 S.n22496 S.n22487 0.002
R50614 S.n22145 S.n22137 0.002
R50615 S.n21473 S.n21464 0.002
R50616 S.n21807 S.n21799 0.002
R50617 S.n20650 S.n20641 0.002
R50618 S.n20997 S.n20989 0.002
R50619 S.n20039 S.n20030 0.002
R50620 S.n19653 S.n19645 0.002
R50621 S.n19185 S.n19176 0.002
R50622 S.n18781 S.n18773 0.002
R50623 S.n18319 S.n18310 0.002
R50624 S.n17898 S.n17890 0.002
R50625 S.n17430 S.n17421 0.002
R50626 S.n16989 S.n16981 0.002
R50627 S.n16528 S.n16519 0.002
R50628 S.n16071 S.n16063 0.002
R50629 S.n15604 S.n15595 0.002
R50630 S.n15127 S.n15119 0.002
R50631 S.n14667 S.n14658 0.002
R50632 S.n14174 S.n14166 0.002
R50633 S.n13708 S.n13699 0.002
R50634 S.n13195 S.n13187 0.002
R50635 S.n12736 S.n12727 0.002
R50636 S.n12207 S.n12199 0.002
R50637 S.n11742 S.n11734 0.002
R50638 S.n22480 S.n22471 0.002
R50639 S.n22160 S.n22152 0.002
R50640 S.n21457 S.n21448 0.002
R50641 S.n21792 S.n21784 0.002
R50642 S.n20634 S.n20625 0.002
R50643 S.n20982 S.n20974 0.002
R50644 S.n20023 S.n20014 0.002
R50645 S.n19668 S.n19660 0.002
R50646 S.n19169 S.n19160 0.002
R50647 S.n18796 S.n18788 0.002
R50648 S.n18303 S.n18294 0.002
R50649 S.n17913 S.n17905 0.002
R50650 S.n17414 S.n17405 0.002
R50651 S.n17004 S.n16996 0.002
R50652 S.n16512 S.n16503 0.002
R50653 S.n16086 S.n16078 0.002
R50654 S.n15588 S.n15579 0.002
R50655 S.n15142 S.n15134 0.002
R50656 S.n14651 S.n14642 0.002
R50657 S.n14189 S.n14181 0.002
R50658 S.n13692 S.n13683 0.002
R50659 S.n13210 S.n13202 0.002
R50660 S.n12720 S.n12711 0.002
R50661 S.n12222 S.n12214 0.002
R50662 S.n11726 S.n11717 0.002
R50663 S.n11208 S.n11200 0.002
R50664 S.n10719 S.n10711 0.002
R50665 S.n22464 S.n22455 0.002
R50666 S.n22175 S.n22167 0.002
R50667 S.n21441 S.n21432 0.002
R50668 S.n21777 S.n21769 0.002
R50669 S.n20618 S.n20609 0.002
R50670 S.n20967 S.n20959 0.002
R50671 S.n20007 S.n19998 0.002
R50672 S.n19683 S.n19675 0.002
R50673 S.n19153 S.n19144 0.002
R50674 S.n18811 S.n18803 0.002
R50675 S.n18287 S.n18278 0.002
R50676 S.n17928 S.n17920 0.002
R50677 S.n17398 S.n17389 0.002
R50678 S.n17019 S.n17011 0.002
R50679 S.n16496 S.n16487 0.002
R50680 S.n16101 S.n16093 0.002
R50681 S.n15572 S.n15563 0.002
R50682 S.n15157 S.n15149 0.002
R50683 S.n14635 S.n14626 0.002
R50684 S.n14204 S.n14196 0.002
R50685 S.n13676 S.n13667 0.002
R50686 S.n13225 S.n13217 0.002
R50687 S.n12704 S.n12695 0.002
R50688 S.n12237 S.n12229 0.002
R50689 S.n11710 S.n11701 0.002
R50690 S.n11223 S.n11215 0.002
R50691 S.n10703 S.n10694 0.002
R50692 S.n10200 S.n10192 0.002
R50693 S.n9674 S.n9666 0.002
R50694 S.n22448 S.n22439 0.002
R50695 S.n22190 S.n22182 0.002
R50696 S.n21425 S.n21416 0.002
R50697 S.n21762 S.n21754 0.002
R50698 S.n20602 S.n20593 0.002
R50699 S.n20952 S.n20944 0.002
R50700 S.n19991 S.n19982 0.002
R50701 S.n19698 S.n19690 0.002
R50702 S.n19137 S.n19128 0.002
R50703 S.n18826 S.n18818 0.002
R50704 S.n18271 S.n18262 0.002
R50705 S.n17943 S.n17935 0.002
R50706 S.n17382 S.n17373 0.002
R50707 S.n17034 S.n17026 0.002
R50708 S.n16480 S.n16471 0.002
R50709 S.n16116 S.n16108 0.002
R50710 S.n15556 S.n15547 0.002
R50711 S.n15172 S.n15164 0.002
R50712 S.n14619 S.n14610 0.002
R50713 S.n14219 S.n14211 0.002
R50714 S.n13660 S.n13651 0.002
R50715 S.n13240 S.n13232 0.002
R50716 S.n12688 S.n12679 0.002
R50717 S.n12252 S.n12244 0.002
R50718 S.n11694 S.n11685 0.002
R50719 S.n11238 S.n11230 0.002
R50720 S.n10687 S.n10678 0.002
R50721 S.n10215 S.n10207 0.002
R50722 S.n9658 S.n9649 0.002
R50723 S.n9166 S.n9158 0.002
R50724 S.n8616 S.n8608 0.002
R50725 S.n22432 S.n22423 0.002
R50726 S.n22205 S.n22197 0.002
R50727 S.n21409 S.n21400 0.002
R50728 S.n21747 S.n21739 0.002
R50729 S.n20586 S.n20577 0.002
R50730 S.n20937 S.n20929 0.002
R50731 S.n19975 S.n19966 0.002
R50732 S.n19713 S.n19705 0.002
R50733 S.n19121 S.n19112 0.002
R50734 S.n18841 S.n18833 0.002
R50735 S.n18255 S.n18246 0.002
R50736 S.n17958 S.n17950 0.002
R50737 S.n17366 S.n17357 0.002
R50738 S.n17049 S.n17041 0.002
R50739 S.n16464 S.n16455 0.002
R50740 S.n16131 S.n16123 0.002
R50741 S.n15540 S.n15531 0.002
R50742 S.n15187 S.n15179 0.002
R50743 S.n14603 S.n14594 0.002
R50744 S.n14234 S.n14226 0.002
R50745 S.n13644 S.n13635 0.002
R50746 S.n13255 S.n13247 0.002
R50747 S.n12672 S.n12663 0.002
R50748 S.n12267 S.n12259 0.002
R50749 S.n11678 S.n11669 0.002
R50750 S.n11253 S.n11245 0.002
R50751 S.n10671 S.n10662 0.002
R50752 S.n10230 S.n10222 0.002
R50753 S.n9642 S.n9633 0.002
R50754 S.n9181 S.n9173 0.002
R50755 S.n8600 S.n8591 0.002
R50756 S.n8123 S.n8115 0.002
R50757 S.n7536 S.n7528 0.002
R50758 S.n22416 S.n22407 0.002
R50759 S.n22220 S.n22212 0.002
R50760 S.n21393 S.n21384 0.002
R50761 S.n21732 S.n21724 0.002
R50762 S.n20570 S.n20561 0.002
R50763 S.n20922 S.n20914 0.002
R50764 S.n19959 S.n19950 0.002
R50765 S.n19728 S.n19720 0.002
R50766 S.n19105 S.n19096 0.002
R50767 S.n18856 S.n18848 0.002
R50768 S.n18239 S.n18230 0.002
R50769 S.n17973 S.n17965 0.002
R50770 S.n17350 S.n17341 0.002
R50771 S.n17064 S.n17056 0.002
R50772 S.n16448 S.n16439 0.002
R50773 S.n16146 S.n16138 0.002
R50774 S.n15524 S.n15515 0.002
R50775 S.n15202 S.n15194 0.002
R50776 S.n14587 S.n14578 0.002
R50777 S.n14249 S.n14241 0.002
R50778 S.n13628 S.n13619 0.002
R50779 S.n13270 S.n13262 0.002
R50780 S.n12656 S.n12647 0.002
R50781 S.n12282 S.n12274 0.002
R50782 S.n11662 S.n11653 0.002
R50783 S.n11268 S.n11260 0.002
R50784 S.n10655 S.n10646 0.002
R50785 S.n10245 S.n10237 0.002
R50786 S.n9626 S.n9617 0.002
R50787 S.n9196 S.n9188 0.002
R50788 S.n8584 S.n8575 0.002
R50789 S.n8138 S.n8130 0.002
R50790 S.n7520 S.n7511 0.002
R50791 S.n7054 S.n7046 0.002
R50792 S.n6443 S.n6435 0.002
R50793 S.n22400 S.n22391 0.002
R50794 S.n22235 S.n22227 0.002
R50795 S.n21377 S.n21368 0.002
R50796 S.n21717 S.n21709 0.002
R50797 S.n20554 S.n20545 0.002
R50798 S.n20907 S.n20899 0.002
R50799 S.n19943 S.n19934 0.002
R50800 S.n19743 S.n19735 0.002
R50801 S.n19089 S.n19080 0.002
R50802 S.n18871 S.n18863 0.002
R50803 S.n18223 S.n18214 0.002
R50804 S.n17988 S.n17980 0.002
R50805 S.n17334 S.n17325 0.002
R50806 S.n17079 S.n17071 0.002
R50807 S.n16432 S.n16423 0.002
R50808 S.n16161 S.n16153 0.002
R50809 S.n15508 S.n15499 0.002
R50810 S.n15217 S.n15209 0.002
R50811 S.n14571 S.n14562 0.002
R50812 S.n14264 S.n14256 0.002
R50813 S.n13612 S.n13603 0.002
R50814 S.n13285 S.n13277 0.002
R50815 S.n12640 S.n12631 0.002
R50816 S.n12297 S.n12289 0.002
R50817 S.n11646 S.n11637 0.002
R50818 S.n11283 S.n11275 0.002
R50819 S.n10639 S.n10630 0.002
R50820 S.n10260 S.n10252 0.002
R50821 S.n9610 S.n9601 0.002
R50822 S.n9211 S.n9203 0.002
R50823 S.n8568 S.n8559 0.002
R50824 S.n8153 S.n8145 0.002
R50825 S.n7504 S.n7495 0.002
R50826 S.n7069 S.n7061 0.002
R50827 S.n6427 S.n6418 0.002
R50828 S.n5976 S.n5968 0.002
R50829 S.n5327 S.n5319 0.002
R50830 S.n22384 S.n22375 0.002
R50831 S.n22250 S.n22242 0.002
R50832 S.n21361 S.n21352 0.002
R50833 S.n21702 S.n21694 0.002
R50834 S.n20538 S.n20529 0.002
R50835 S.n20892 S.n20884 0.002
R50836 S.n19927 S.n19918 0.002
R50837 S.n19758 S.n19750 0.002
R50838 S.n19073 S.n19064 0.002
R50839 S.n18886 S.n18878 0.002
R50840 S.n18207 S.n18198 0.002
R50841 S.n18003 S.n17995 0.002
R50842 S.n17318 S.n17309 0.002
R50843 S.n17094 S.n17086 0.002
R50844 S.n16416 S.n16407 0.002
R50845 S.n16176 S.n16168 0.002
R50846 S.n15492 S.n15483 0.002
R50847 S.n15232 S.n15224 0.002
R50848 S.n14555 S.n14546 0.002
R50849 S.n14279 S.n14271 0.002
R50850 S.n13596 S.n13587 0.002
R50851 S.n13300 S.n13292 0.002
R50852 S.n12624 S.n12615 0.002
R50853 S.n12312 S.n12304 0.002
R50854 S.n11630 S.n11621 0.002
R50855 S.n11298 S.n11290 0.002
R50856 S.n10623 S.n10614 0.002
R50857 S.n10275 S.n10267 0.002
R50858 S.n9594 S.n9585 0.002
R50859 S.n9229 S.n9221 0.002
R50860 S.n8552 S.n8543 0.002
R50861 S.n8168 S.n8160 0.002
R50862 S.n7488 S.n7479 0.002
R50863 S.n7084 S.n7076 0.002
R50864 S.n6411 S.n6402 0.002
R50865 S.n5991 S.n5983 0.002
R50866 S.n5311 S.n5302 0.002
R50867 S.n4871 S.n4863 0.002
R50868 S.n4198 S.n4190 0.002
R50869 S.n22672 S.n22265 0.002
R50870 S.n22675 S.n22257 0.002
R50871 S.n21685 S.n21671 0.002
R50872 S.n21687 S.n21663 0.002
R50873 S.n20522 S.n20514 0.002
R50874 S.n20877 S.n20868 0.002
R50875 S.n19911 S.n19903 0.002
R50876 S.n19774 S.n19765 0.002
R50877 S.n19057 S.n19049 0.002
R50878 S.n18902 S.n18893 0.002
R50879 S.n18191 S.n18183 0.002
R50880 S.n18019 S.n18010 0.002
R50881 S.n17302 S.n17294 0.002
R50882 S.n17110 S.n17101 0.002
R50883 S.n16400 S.n16392 0.002
R50884 S.n16192 S.n16183 0.002
R50885 S.n15476 S.n15468 0.002
R50886 S.n15248 S.n15239 0.002
R50887 S.n14539 S.n14531 0.002
R50888 S.n14295 S.n14286 0.002
R50889 S.n13580 S.n13572 0.002
R50890 S.n13316 S.n13307 0.002
R50891 S.n12608 S.n12600 0.002
R50892 S.n12328 S.n12319 0.002
R50893 S.n11614 S.n11606 0.002
R50894 S.n11314 S.n11305 0.002
R50895 S.n10607 S.n10599 0.002
R50896 S.n10291 S.n10282 0.002
R50897 S.n9578 S.n9570 0.002
R50898 S.n9242 S.n9233 0.002
R50899 S.n8536 S.n8528 0.002
R50900 S.n8184 S.n8175 0.002
R50901 S.n7472 S.n7464 0.002
R50902 S.n7100 S.n7091 0.002
R50903 S.n6395 S.n6387 0.002
R50904 S.n6007 S.n5998 0.002
R50905 S.n5295 S.n5287 0.002
R50906 S.n4887 S.n4878 0.002
R50907 S.n4182 S.n4174 0.002
R50908 S.n3759 S.n3750 0.002
R50909 S.n22368 S.n22358 0.002
R50910 S.n22694 S.n22682 0.002
R50911 S.n21654 S.n21276 0.002
R50912 S.n21656 S.n21268 0.002
R50913 S.n20507 S.n20499 0.002
R50914 S.n20861 S.n20852 0.002
R50915 S.n19896 S.n19888 0.002
R50916 S.n19790 S.n19781 0.002
R50917 S.n19042 S.n19034 0.002
R50918 S.n18918 S.n18909 0.002
R50919 S.n18176 S.n18168 0.002
R50920 S.n18035 S.n18026 0.002
R50921 S.n17287 S.n17279 0.002
R50922 S.n17126 S.n17117 0.002
R50923 S.n16385 S.n16377 0.002
R50924 S.n16208 S.n16199 0.002
R50925 S.n15461 S.n15453 0.002
R50926 S.n15264 S.n15255 0.002
R50927 S.n14524 S.n14516 0.002
R50928 S.n14311 S.n14302 0.002
R50929 S.n13565 S.n13557 0.002
R50930 S.n13332 S.n13323 0.002
R50931 S.n12593 S.n12585 0.002
R50932 S.n12344 S.n12335 0.002
R50933 S.n11599 S.n11591 0.002
R50934 S.n11330 S.n11321 0.002
R50935 S.n10592 S.n10584 0.002
R50936 S.n10307 S.n10298 0.002
R50937 S.n9563 S.n9555 0.002
R50938 S.n9258 S.n9249 0.002
R50939 S.n8521 S.n8513 0.002
R50940 S.n8200 S.n8191 0.002
R50941 S.n7457 S.n7449 0.002
R50942 S.n7116 S.n7107 0.002
R50943 S.n6380 S.n6372 0.002
R50944 S.n6023 S.n6014 0.002
R50945 S.n5280 S.n5272 0.002
R50946 S.n4903 S.n4894 0.002
R50947 S.n4167 S.n4159 0.002
R50948 S.n3775 S.n3766 0.002
R50949 S.n3041 S.n3033 0.002
R50950 S.n2628 S.n2619 0.002
R50951 S.n1931 S.n1919 0.002
R50952 S.n1882 S.n1874 0.002
R50953 S.n3084 S.n3076 0.002
R50954 S.n3074 S.n2635 0.002
R50955 S.n4225 S.n4217 0.002
R50956 S.n4215 S.n3782 0.002
R50957 S.n5354 S.n5346 0.002
R50958 S.n5344 S.n4910 0.002
R50959 S.n6470 S.n6462 0.002
R50960 S.n6460 S.n6030 0.002
R50961 S.n7563 S.n7555 0.002
R50962 S.n7553 S.n7123 0.002
R50963 S.n8643 S.n8635 0.002
R50964 S.n8633 S.n8207 0.002
R50965 S.n9701 S.n9693 0.002
R50966 S.n9691 S.n9265 0.002
R50967 S.n10746 S.n10738 0.002
R50968 S.n10736 S.n10314 0.002
R50969 S.n11769 S.n11761 0.002
R50970 S.n11759 S.n11337 0.002
R50971 S.n12779 S.n12771 0.002
R50972 S.n12769 S.n12351 0.002
R50973 S.n13767 S.n13759 0.002
R50974 S.n13757 S.n13339 0.002
R50975 S.n14742 S.n14734 0.002
R50976 S.n14732 S.n14318 0.002
R50977 S.n15695 S.n15687 0.002
R50978 S.n15685 S.n15271 0.002
R50979 S.n16635 S.n16627 0.002
R50980 S.n16625 S.n16215 0.002
R50981 S.n17553 S.n17545 0.002
R50982 S.n17543 S.n17133 0.002
R50983 S.n18458 S.n18450 0.002
R50984 S.n18448 S.n18042 0.002
R50985 S.n19340 S.n19332 0.002
R50986 S.n19330 S.n18925 0.002
R50987 S.n20210 S.n20202 0.002
R50988 S.n20200 S.n19797 0.002
R50989 S.n20845 S.n20837 0.002
R50990 S.n20835 S.n20431 0.002
R50991 S.n21261 S.n21253 0.002
R50992 S.n21345 S.n21337 0.002
R50993 S.n22713 S.n22705 0.002
R50994 S.n22351 S.n22343 0.002
R50995 S.n25 S.n24 0.002
R50996 S.n743 S.n735 0.002
R50997 S.n2107 S.n2086 0.002
R50998 S.n1776 S.n1766 0.002
R50999 S.n3259 S.n3242 0.002
R51000 S.n2942 S.n2934 0.002
R51001 S.n4396 S.n4379 0.002
R51002 S.n4069 S.n4061 0.002
R51003 S.n5531 S.n5514 0.002
R51004 S.n5181 S.n5173 0.002
R51005 S.n6641 S.n6624 0.002
R51006 S.n6281 S.n6273 0.002
R51007 S.n7739 S.n7722 0.002
R51008 S.n7358 S.n7350 0.002
R51009 S.n8814 S.n8797 0.002
R51010 S.n8422 S.n8414 0.002
R51011 S.n9877 S.n9860 0.002
R51012 S.n9464 S.n9456 0.002
R51013 S.n10917 S.n10900 0.002
R51014 S.n10493 S.n10485 0.002
R51015 S.n11945 S.n11928 0.002
R51016 S.n11500 S.n11492 0.002
R51017 S.n12950 S.n12933 0.002
R51018 S.n12494 S.n12486 0.002
R51019 S.n13943 S.n13926 0.002
R51020 S.n13466 S.n13458 0.002
R51021 S.n14913 S.n14896 0.002
R51022 S.n14425 S.n14417 0.002
R51023 S.n15871 S.n15854 0.002
R51024 S.n15362 S.n15354 0.002
R51025 S.n16806 S.n16789 0.002
R51026 S.n16286 S.n16278 0.002
R51027 S.n17733 S.n17716 0.002
R51028 S.n17188 S.n17180 0.002
R51029 S.n18633 S.n18616 0.002
R51030 S.n18077 S.n18069 0.002
R51031 S.n1338 S.n1337 0.002
R51032 S.n767 S.n751 0.002
R51033 S.n2045 S.n2030 0.002
R51034 S.n1823 S.n1806 0.002
R51035 S.n3198 S.n3173 0.002
R51036 S.n2986 S.n2968 0.002
R51037 S.n4335 S.n4310 0.002
R51038 S.n4113 S.n4095 0.002
R51039 S.n5470 S.n5445 0.002
R51040 S.n5225 S.n5207 0.002
R51041 S.n6580 S.n6555 0.002
R51042 S.n6325 S.n6307 0.002
R51043 S.n7678 S.n7653 0.002
R51044 S.n7402 S.n7384 0.002
R51045 S.n8753 S.n8728 0.002
R51046 S.n8466 S.n8448 0.002
R51047 S.n9816 S.n9791 0.002
R51048 S.n9508 S.n9490 0.002
R51049 S.n10856 S.n10831 0.002
R51050 S.n10537 S.n10519 0.002
R51051 S.n11884 S.n11859 0.002
R51052 S.n11544 S.n11526 0.002
R51053 S.n12889 S.n12864 0.002
R51054 S.n12538 S.n12520 0.002
R51055 S.n13882 S.n13857 0.002
R51056 S.n13510 S.n13492 0.002
R51057 S.n14852 S.n14827 0.002
R51058 S.n14469 S.n14451 0.002
R51059 S.n15810 S.n15785 0.002
R51060 S.n15406 S.n15388 0.002
R51061 S.n16745 S.n16720 0.002
R51062 S.n16330 S.n16312 0.002
R51063 S.n17668 S.n17643 0.002
R51064 S.n17232 S.n17214 0.002
R51065 S.n18568 S.n18543 0.002
R51066 S.n18121 S.n18103 0.002
R51067 S.n19458 S.n19430 0.002
R51068 S.n18987 S.n18968 0.002
R51069 S.n20330 S.n20302 0.002
R51070 S.n19839 S.n19820 0.002
R51071 S.n20472 S.n20461 0.002
R51072 S.n20366 S.n20358 0.002
R51073 S.n19861 S.n19850 0.002
R51074 S.n20295 S.n20287 0.002
R51075 S.n19007 S.n18996 0.002
R51076 S.n19423 S.n19415 0.002
R51077 S.n18141 S.n18130 0.002
R51078 S.n18536 S.n18528 0.002
R51079 S.n17252 S.n17241 0.002
R51080 S.n17636 S.n17628 0.002
R51081 S.n16350 S.n16339 0.002
R51082 S.n16713 S.n16705 0.002
R51083 S.n15426 S.n15415 0.002
R51084 S.n15778 S.n15770 0.002
R51085 S.n14489 S.n14478 0.002
R51086 S.n14820 S.n14812 0.002
R51087 S.n13530 S.n13519 0.002
R51088 S.n13850 S.n13842 0.002
R51089 S.n12558 S.n12547 0.002
R51090 S.n12857 S.n12849 0.002
R51091 S.n11564 S.n11553 0.002
R51092 S.n11852 S.n11844 0.002
R51093 S.n10557 S.n10546 0.002
R51094 S.n10824 S.n10816 0.002
R51095 S.n9528 S.n9517 0.002
R51096 S.n9784 S.n9776 0.002
R51097 S.n8486 S.n8475 0.002
R51098 S.n8721 S.n8713 0.002
R51099 S.n7422 S.n7411 0.002
R51100 S.n7646 S.n7638 0.002
R51101 S.n6345 S.n6334 0.002
R51102 S.n6548 S.n6540 0.002
R51103 S.n5245 S.n5234 0.002
R51104 S.n5438 S.n5429 0.002
R51105 S.n4132 S.n4122 0.002
R51106 S.n4303 S.n4295 0.002
R51107 S.n3006 S.n2995 0.002
R51108 S.n3166 S.n3158 0.002
R51109 S.n1845 S.n1830 0.002
R51110 S.n2012 S.n1997 0.002
R51111 S.n786 S.n775 0.002
R51112 S.n72 S.n71 0.002
R51113 S.n708 S.n700 0.002
R51114 S.n2166 S.n2144 0.002
R51115 S.n1737 S.n1729 0.002
R51116 S.n3319 S.n3302 0.002
R51117 S.n2906 S.n2898 0.002
R51118 S.n4457 S.n4440 0.002
R51119 S.n4033 S.n4025 0.002
R51120 S.n5592 S.n5575 0.002
R51121 S.n5145 S.n5137 0.002
R51122 S.n6702 S.n6685 0.002
R51123 S.n6245 S.n6237 0.002
R51124 S.n7800 S.n7783 0.002
R51125 S.n7322 S.n7314 0.002
R51126 S.n8875 S.n8858 0.002
R51127 S.n8386 S.n8378 0.002
R51128 S.n9938 S.n9921 0.002
R51129 S.n9428 S.n9420 0.002
R51130 S.n10978 S.n10961 0.002
R51131 S.n10457 S.n10449 0.002
R51132 S.n12006 S.n11989 0.002
R51133 S.n11464 S.n11456 0.002
R51134 S.n13011 S.n12994 0.002
R51135 S.n12458 S.n12450 0.002
R51136 S.n14004 S.n13987 0.002
R51137 S.n13430 S.n13422 0.002
R51138 S.n14974 S.n14957 0.002
R51139 S.n14389 S.n14381 0.002
R51140 S.n15936 S.n15919 0.002
R51141 S.n15326 S.n15318 0.002
R51142 S.n16871 S.n16854 0.002
R51143 S.n16250 S.n16242 0.002
R51144 S.n104 S.n103 0.002
R51145 S.n673 S.n665 0.002
R51146 S.n2225 S.n2203 0.002
R51147 S.n1700 S.n1692 0.002
R51148 S.n3379 S.n3362 0.002
R51149 S.n2870 S.n2862 0.002
R51150 S.n4518 S.n4501 0.002
R51151 S.n3997 S.n3989 0.002
R51152 S.n5653 S.n5636 0.002
R51153 S.n5109 S.n5101 0.002
R51154 S.n6763 S.n6746 0.002
R51155 S.n6209 S.n6201 0.002
R51156 S.n7861 S.n7844 0.002
R51157 S.n7286 S.n7278 0.002
R51158 S.n8936 S.n8919 0.002
R51159 S.n8350 S.n8342 0.002
R51160 S.n9999 S.n9982 0.002
R51161 S.n9392 S.n9384 0.002
R51162 S.n11039 S.n11022 0.002
R51163 S.n10421 S.n10413 0.002
R51164 S.n12067 S.n12050 0.002
R51165 S.n11428 S.n11420 0.002
R51166 S.n13072 S.n13055 0.002
R51167 S.n12422 S.n12414 0.002
R51168 S.n14069 S.n14052 0.002
R51169 S.n13394 S.n13386 0.002
R51170 S.n15039 S.n15022 0.002
R51171 S.n14353 S.n14345 0.002
R51172 S.n991 S.n990 0.002
R51173 S.n638 S.n630 0.002
R51174 S.n2284 S.n2262 0.002
R51175 S.n1663 S.n1655 0.002
R51176 S.n3439 S.n3422 0.002
R51177 S.n2834 S.n2826 0.002
R51178 S.n4579 S.n4562 0.002
R51179 S.n3961 S.n3953 0.002
R51180 S.n5714 S.n5697 0.002
R51181 S.n5073 S.n5065 0.002
R51182 S.n6824 S.n6807 0.002
R51183 S.n6173 S.n6165 0.002
R51184 S.n7922 S.n7905 0.002
R51185 S.n7250 S.n7242 0.002
R51186 S.n8997 S.n8980 0.002
R51187 S.n8314 S.n8306 0.002
R51188 S.n10060 S.n10043 0.002
R51189 S.n9356 S.n9348 0.002
R51190 S.n11100 S.n11083 0.002
R51191 S.n10385 S.n10377 0.002
R51192 S.n12132 S.n12115 0.002
R51193 S.n11392 S.n11384 0.002
R51194 S.n13137 S.n13120 0.002
R51195 S.n12386 S.n12378 0.002
R51196 S.n1023 S.n1022 0.002
R51197 S.n603 S.n595 0.002
R51198 S.n2343 S.n2321 0.002
R51199 S.n1626 S.n1618 0.002
R51200 S.n3499 S.n3482 0.002
R51201 S.n2798 S.n2790 0.002
R51202 S.n4640 S.n4623 0.002
R51203 S.n3925 S.n3917 0.002
R51204 S.n5775 S.n5758 0.002
R51205 S.n5037 S.n5029 0.002
R51206 S.n6885 S.n6868 0.002
R51207 S.n6137 S.n6129 0.002
R51208 S.n7983 S.n7966 0.002
R51209 S.n7214 S.n7206 0.002
R51210 S.n9058 S.n9041 0.002
R51211 S.n8278 S.n8270 0.002
R51212 S.n10125 S.n10108 0.002
R51213 S.n9320 S.n9312 0.002
R51214 S.n11165 S.n11148 0.002
R51215 S.n10349 S.n10341 0.002
R51216 S.n1055 S.n1054 0.002
R51217 S.n568 S.n560 0.002
R51218 S.n2402 S.n2380 0.002
R51219 S.n1589 S.n1581 0.002
R51220 S.n3559 S.n3542 0.002
R51221 S.n2762 S.n2754 0.002
R51222 S.n4701 S.n4684 0.002
R51223 S.n3889 S.n3881 0.002
R51224 S.n5836 S.n5819 0.002
R51225 S.n5001 S.n4993 0.002
R51226 S.n6946 S.n6929 0.002
R51227 S.n6101 S.n6093 0.002
R51228 S.n8048 S.n8031 0.002
R51229 S.n7178 S.n7170 0.002
R51230 S.n9123 S.n9106 0.002
R51231 S.n8242 S.n8234 0.002
R51232 S.n1087 S.n1086 0.002
R51233 S.n533 S.n525 0.002
R51234 S.n2461 S.n2439 0.002
R51235 S.n1552 S.n1544 0.002
R51236 S.n3619 S.n3602 0.002
R51237 S.n2726 S.n2718 0.002
R51238 S.n4762 S.n4745 0.002
R51239 S.n3853 S.n3845 0.002
R51240 S.n5901 S.n5884 0.002
R51241 S.n4965 S.n4957 0.002
R51242 S.n7011 S.n6994 0.002
R51243 S.n6065 S.n6057 0.002
R51244 S.n1119 S.n1118 0.002
R51245 S.n498 S.n490 0.002
R51246 S.n2520 S.n2498 0.002
R51247 S.n1515 S.n1507 0.002
R51248 S.n3683 S.n3666 0.002
R51249 S.n2690 S.n2682 0.002
R51250 S.n4827 S.n4810 0.002
R51251 S.n3817 S.n3809 0.002
R51252 S.n1157 S.n1156 0.002
R51253 S.n463 S.n454 0.002
R51254 S.n2583 S.n2566 0.002
R51255 S.n1478 S.n1470 0.002
R51256 S.n22765 S.n22757 0.002
R51257 S.n22307 S.n22295 0.002
R51258 S.n22978 S.n22977 0.002
R51259 S.n19370 S.n19355 0.002
R51260 S.n20424 S.n20406 0.002
R51261 S.n21242 S.n21234 0.002
R51262 S.n17583 S.n17568 0.002
R51263 S.n15725 S.n15710 0.002
R51264 S.n13797 S.n13782 0.002
R51265 S.n11799 S.n11784 0.002
R51266 S.n9731 S.n9716 0.002
R51267 S.n7593 S.n7578 0.002
R51268 S.n5384 S.n5369 0.002
R51269 S.n3114 S.n3099 0.002
R51270 S.n911 S.n910 0.002
R51271 S.n389 S.n388 0.002
R51272 S.n357 S.n356 0.002
R51273 S.n325 S.n324 0.002
R51274 S.n293 S.n292 0.002
R51275 S.n261 S.n260 0.002
R51276 S.n232 S.n231 0.002
R51277 S.n197 S.n196 0.002
R51278 S.n165 S.n164 0.002
R51279 S.n133 S.n132 0.002
R51280 S.n22298 S.n22297 0.002
R51281 S.n22320 S.n22319 0.002
R51282 S.n2038 S.n2037 0.002
R51283 S.n20395 S.n20394 0.002
R51284 S.n21214 S.n21213 0.002
R51285 S.n22735 S.n22734 0.002
R51286 S.n18597 S.n18596 0.002
R51287 S.n19487 S.n19486 0.002
R51288 S.n20232 S.n20231 0.002
R51289 S.n16835 S.n16834 0.002
R51290 S.n17762 S.n17761 0.002
R51291 S.n18477 S.n18476 0.002
R51292 S.n15003 S.n15002 0.002
R51293 S.n15965 S.n15964 0.002
R51294 S.n16654 S.n16653 0.002
R51295 S.n13101 S.n13100 0.002
R51296 S.n14098 S.n14097 0.002
R51297 S.n14761 S.n14760 0.002
R51298 S.n11129 S.n11128 0.002
R51299 S.n12161 S.n12160 0.002
R51300 S.n12798 S.n12797 0.002
R51301 S.n9087 S.n9086 0.002
R51302 S.n10154 S.n10153 0.002
R51303 S.n10765 S.n10764 0.002
R51304 S.n6975 S.n6974 0.002
R51305 S.n8077 S.n8076 0.002
R51306 S.n8662 S.n8661 0.002
R51307 S.n4791 S.n4790 0.002
R51308 S.n5930 S.n5929 0.002
R51309 S.n6489 S.n6488 0.002
R51310 S.n3711 S.n3710 0.002
R51311 S.n4244 S.n4243 0.002
R51312 S.n21962 S.n21961 0.002
R51313 S.n21638 S.n21637 0.002
R51314 S.n21995 S.n21994 0.002
R51315 S.n22656 S.n22655 0.002
R51316 S.n19533 S.n19526 0.002
R51317 S.n18676 S.n18669 0.002
R51318 S.n17808 S.n17801 0.002
R51319 S.n16914 S.n16907 0.002
R51320 S.n16011 S.n16004 0.002
R51321 S.n15082 S.n15075 0.002
R51322 S.n14144 S.n14137 0.002
R51323 S.n13180 S.n13173 0.002
R51324 S.n12207 S.n12200 0.002
R51325 S.n11208 S.n11201 0.002
R51326 S.n10200 S.n10193 0.002
R51327 S.n9166 S.n9159 0.002
R51328 S.n8123 S.n8116 0.002
R51329 S.n7054 S.n7047 0.002
R51330 S.n5976 S.n5969 0.002
R51331 S.n4871 S.n4864 0.002
R51332 S.n3759 S.n3751 0.002
R51333 S.n2628 S.n2620 0.002
R51334 S.n1985 S.n1972 0.002
R51335 S.n2137 S.n2124 0.002
R51336 S.n3259 S.n3258 0.002
R51337 S.n2942 S.n2941 0.002
R51338 S.n4396 S.n4395 0.002
R51339 S.n4069 S.n4068 0.002
R51340 S.n5531 S.n5530 0.002
R51341 S.n5181 S.n5180 0.002
R51342 S.n6641 S.n6640 0.002
R51343 S.n6281 S.n6280 0.002
R51344 S.n7739 S.n7738 0.002
R51345 S.n7358 S.n7357 0.002
R51346 S.n8814 S.n8813 0.002
R51347 S.n8422 S.n8421 0.002
R51348 S.n9877 S.n9876 0.002
R51349 S.n9464 S.n9463 0.002
R51350 S.n10917 S.n10916 0.002
R51351 S.n10493 S.n10492 0.002
R51352 S.n11945 S.n11944 0.002
R51353 S.n11500 S.n11499 0.002
R51354 S.n12950 S.n12949 0.002
R51355 S.n12494 S.n12493 0.002
R51356 S.n13943 S.n13942 0.002
R51357 S.n13466 S.n13465 0.002
R51358 S.n14913 S.n14912 0.002
R51359 S.n14425 S.n14424 0.002
R51360 S.n15871 S.n15870 0.002
R51361 S.n15362 S.n15361 0.002
R51362 S.n16806 S.n16805 0.002
R51363 S.n16286 S.n16285 0.002
R51364 S.n17733 S.n17732 0.002
R51365 S.n17188 S.n17187 0.002
R51366 S.n18633 S.n18632 0.002
R51367 S.n18077 S.n18076 0.002
R51368 S.n2196 S.n2183 0.002
R51369 S.n1737 S.n1736 0.002
R51370 S.n3319 S.n3318 0.002
R51371 S.n2906 S.n2905 0.002
R51372 S.n4457 S.n4456 0.002
R51373 S.n4033 S.n4032 0.002
R51374 S.n5592 S.n5591 0.002
R51375 S.n5145 S.n5144 0.002
R51376 S.n6702 S.n6701 0.002
R51377 S.n6245 S.n6244 0.002
R51378 S.n7800 S.n7799 0.002
R51379 S.n7322 S.n7321 0.002
R51380 S.n8875 S.n8874 0.002
R51381 S.n8386 S.n8385 0.002
R51382 S.n9938 S.n9937 0.002
R51383 S.n9428 S.n9427 0.002
R51384 S.n10978 S.n10977 0.002
R51385 S.n10457 S.n10456 0.002
R51386 S.n12006 S.n12005 0.002
R51387 S.n11464 S.n11463 0.002
R51388 S.n13011 S.n13010 0.002
R51389 S.n12458 S.n12457 0.002
R51390 S.n14004 S.n14003 0.002
R51391 S.n13430 S.n13429 0.002
R51392 S.n14974 S.n14973 0.002
R51393 S.n14389 S.n14388 0.002
R51394 S.n15936 S.n15935 0.002
R51395 S.n15326 S.n15325 0.002
R51396 S.n16871 S.n16870 0.002
R51397 S.n16250 S.n16249 0.002
R51398 S.n2255 S.n2242 0.002
R51399 S.n1700 S.n1699 0.002
R51400 S.n3379 S.n3378 0.002
R51401 S.n2870 S.n2869 0.002
R51402 S.n4518 S.n4517 0.002
R51403 S.n3997 S.n3996 0.002
R51404 S.n5653 S.n5652 0.002
R51405 S.n5109 S.n5108 0.002
R51406 S.n6763 S.n6762 0.002
R51407 S.n6209 S.n6208 0.002
R51408 S.n7861 S.n7860 0.002
R51409 S.n7286 S.n7285 0.002
R51410 S.n8936 S.n8935 0.002
R51411 S.n8350 S.n8349 0.002
R51412 S.n9999 S.n9998 0.002
R51413 S.n9392 S.n9391 0.002
R51414 S.n11039 S.n11038 0.002
R51415 S.n10421 S.n10420 0.002
R51416 S.n12067 S.n12066 0.002
R51417 S.n11428 S.n11427 0.002
R51418 S.n13072 S.n13071 0.002
R51419 S.n12422 S.n12421 0.002
R51420 S.n14069 S.n14068 0.002
R51421 S.n13394 S.n13393 0.002
R51422 S.n15039 S.n15038 0.002
R51423 S.n14353 S.n14352 0.002
R51424 S.n2314 S.n2301 0.002
R51425 S.n1663 S.n1662 0.002
R51426 S.n3439 S.n3438 0.002
R51427 S.n2834 S.n2833 0.002
R51428 S.n4579 S.n4578 0.002
R51429 S.n3961 S.n3960 0.002
R51430 S.n5714 S.n5713 0.002
R51431 S.n5073 S.n5072 0.002
R51432 S.n6824 S.n6823 0.002
R51433 S.n6173 S.n6172 0.002
R51434 S.n7922 S.n7921 0.002
R51435 S.n7250 S.n7249 0.002
R51436 S.n8997 S.n8996 0.002
R51437 S.n8314 S.n8313 0.002
R51438 S.n10060 S.n10059 0.002
R51439 S.n9356 S.n9355 0.002
R51440 S.n11100 S.n11099 0.002
R51441 S.n10385 S.n10384 0.002
R51442 S.n12132 S.n12131 0.002
R51443 S.n11392 S.n11391 0.002
R51444 S.n13137 S.n13136 0.002
R51445 S.n12386 S.n12385 0.002
R51446 S.n2373 S.n2360 0.002
R51447 S.n1626 S.n1625 0.002
R51448 S.n3499 S.n3498 0.002
R51449 S.n2798 S.n2797 0.002
R51450 S.n4640 S.n4639 0.002
R51451 S.n3925 S.n3924 0.002
R51452 S.n5775 S.n5774 0.002
R51453 S.n5037 S.n5036 0.002
R51454 S.n6885 S.n6884 0.002
R51455 S.n6137 S.n6136 0.002
R51456 S.n7983 S.n7982 0.002
R51457 S.n7214 S.n7213 0.002
R51458 S.n9058 S.n9057 0.002
R51459 S.n8278 S.n8277 0.002
R51460 S.n10125 S.n10124 0.002
R51461 S.n9320 S.n9319 0.002
R51462 S.n11165 S.n11164 0.002
R51463 S.n10349 S.n10348 0.002
R51464 S.n2432 S.n2419 0.002
R51465 S.n1589 S.n1588 0.002
R51466 S.n3559 S.n3558 0.002
R51467 S.n2762 S.n2761 0.002
R51468 S.n4701 S.n4700 0.002
R51469 S.n3889 S.n3888 0.002
R51470 S.n5836 S.n5835 0.002
R51471 S.n5001 S.n5000 0.002
R51472 S.n6946 S.n6945 0.002
R51473 S.n6101 S.n6100 0.002
R51474 S.n8048 S.n8047 0.002
R51475 S.n7178 S.n7177 0.002
R51476 S.n9123 S.n9122 0.002
R51477 S.n8242 S.n8241 0.002
R51478 S.n2491 S.n2478 0.002
R51479 S.n1552 S.n1551 0.002
R51480 S.n3619 S.n3618 0.002
R51481 S.n2726 S.n2725 0.002
R51482 S.n4762 S.n4761 0.002
R51483 S.n3853 S.n3852 0.002
R51484 S.n5901 S.n5900 0.002
R51485 S.n4965 S.n4964 0.002
R51486 S.n7011 S.n7010 0.002
R51487 S.n6065 S.n6064 0.002
R51488 S.n2550 S.n2537 0.002
R51489 S.n1515 S.n1514 0.002
R51490 S.n3683 S.n3682 0.002
R51491 S.n2690 S.n2689 0.002
R51492 S.n4827 S.n4826 0.002
R51493 S.n3817 S.n3816 0.002
R51494 S.n2583 S.n2582 0.002
R51495 S.n1478 S.n1477 0.002
R51496 S.n22328 S.n22327 0.002
R51497 S.n3178 S.n3177 0.002
R51498 S.n4315 S.n4314 0.002
R51499 S.n5450 S.n5449 0.002
R51500 S.n6560 S.n6559 0.002
R51501 S.n7658 S.n7657 0.002
R51502 S.n8733 S.n8732 0.002
R51503 S.n9796 S.n9795 0.002
R51504 S.n10836 S.n10835 0.002
R51505 S.n11864 S.n11863 0.002
R51506 S.n12869 S.n12868 0.002
R51507 S.n13862 S.n13861 0.002
R51508 S.n14832 S.n14831 0.002
R51509 S.n15790 S.n15789 0.002
R51510 S.n16725 S.n16724 0.002
R51511 S.n17648 S.n17647 0.002
R51512 S.n18548 S.n18547 0.002
R51513 S.n19435 S.n19434 0.002
R51514 S.n20307 S.n20306 0.002
R51515 S.n20411 S.n20410 0.002
R51516 S.n19354 S.n19353 0.002
R51517 S.n18615 S.n18614 0.002
R51518 S.n17715 S.n17714 0.002
R51519 S.n17567 S.n17566 0.002
R51520 S.n16853 S.n16852 0.002
R51521 S.n15918 S.n15917 0.002
R51522 S.n15709 S.n15708 0.002
R51523 S.n15021 S.n15020 0.002
R51524 S.n14051 S.n14050 0.002
R51525 S.n13781 S.n13780 0.002
R51526 S.n13119 S.n13118 0.002
R51527 S.n12114 S.n12113 0.002
R51528 S.n11783 S.n11782 0.002
R51529 S.n11147 S.n11146 0.002
R51530 S.n10107 S.n10106 0.002
R51531 S.n9715 S.n9714 0.002
R51532 S.n9105 S.n9104 0.002
R51533 S.n8030 S.n8029 0.002
R51534 S.n7577 S.n7576 0.002
R51535 S.n6993 S.n6992 0.002
R51536 S.n5883 S.n5882 0.002
R51537 S.n5368 S.n5367 0.002
R51538 S.n4809 S.n4808 0.002
R51539 S.n3665 S.n3664 0.002
R51540 S.n3098 S.n3097 0.002
R51541 S.n2565 S.n2564 0.002
R51542 S.n22640 S.n22632 0.002
R51543 S.n22010 S.n22003 0.002
R51544 S.n21617 S.n21609 0.002
R51545 S.n21942 S.n21935 0.002
R51546 S.n20794 S.n20786 0.002
R51547 S.n20183 S.n20182 0.002
R51548 S.n22624 S.n22616 0.002
R51549 S.n22025 S.n22018 0.002
R51550 S.n21601 S.n21593 0.002
R51551 S.n21927 S.n21920 0.002
R51552 S.n20778 S.n20770 0.002
R51553 S.n21117 S.n21110 0.002
R51554 S.n20167 S.n20159 0.002
R51555 S.n19313 S.n19312 0.002
R51556 S.n22608 S.n22600 0.002
R51557 S.n22040 S.n22033 0.002
R51558 S.n21585 S.n21577 0.002
R51559 S.n21912 S.n21905 0.002
R51560 S.n20762 S.n20754 0.002
R51561 S.n21102 S.n21095 0.002
R51562 S.n20151 S.n20143 0.002
R51563 S.n19548 S.n19541 0.002
R51564 S.n19297 S.n19289 0.002
R51565 S.n18431 S.n18430 0.002
R51566 S.n22592 S.n22584 0.002
R51567 S.n22055 S.n22048 0.002
R51568 S.n21569 S.n21561 0.002
R51569 S.n21897 S.n21890 0.002
R51570 S.n20746 S.n20738 0.002
R51571 S.n21087 S.n21080 0.002
R51572 S.n20135 S.n20127 0.002
R51573 S.n19563 S.n19556 0.002
R51574 S.n19281 S.n19273 0.002
R51575 S.n18691 S.n18684 0.002
R51576 S.n18415 S.n18407 0.002
R51577 S.n17526 S.n17525 0.002
R51578 S.n22576 S.n22568 0.002
R51579 S.n22070 S.n22063 0.002
R51580 S.n21553 S.n21545 0.002
R51581 S.n21882 S.n21875 0.002
R51582 S.n20730 S.n20722 0.002
R51583 S.n21072 S.n21065 0.002
R51584 S.n20119 S.n20111 0.002
R51585 S.n19578 S.n19571 0.002
R51586 S.n19265 S.n19257 0.002
R51587 S.n18706 S.n18699 0.002
R51588 S.n18399 S.n18391 0.002
R51589 S.n17823 S.n17816 0.002
R51590 S.n17510 S.n17502 0.002
R51591 S.n16608 S.n16607 0.002
R51592 S.n22560 S.n22552 0.002
R51593 S.n22085 S.n22078 0.002
R51594 S.n21537 S.n21529 0.002
R51595 S.n21867 S.n21860 0.002
R51596 S.n20714 S.n20706 0.002
R51597 S.n21057 S.n21050 0.002
R51598 S.n20103 S.n20095 0.002
R51599 S.n19593 S.n19586 0.002
R51600 S.n19249 S.n19241 0.002
R51601 S.n18721 S.n18714 0.002
R51602 S.n18383 S.n18375 0.002
R51603 S.n17838 S.n17831 0.002
R51604 S.n17494 S.n17486 0.002
R51605 S.n16929 S.n16922 0.002
R51606 S.n16592 S.n16584 0.002
R51607 S.n15668 S.n15667 0.002
R51608 S.n22544 S.n22536 0.002
R51609 S.n22100 S.n22093 0.002
R51610 S.n21521 S.n21513 0.002
R51611 S.n21852 S.n21845 0.002
R51612 S.n20698 S.n20690 0.002
R51613 S.n21042 S.n21035 0.002
R51614 S.n20087 S.n20079 0.002
R51615 S.n19608 S.n19601 0.002
R51616 S.n19233 S.n19225 0.002
R51617 S.n18736 S.n18729 0.002
R51618 S.n18367 S.n18359 0.002
R51619 S.n17853 S.n17846 0.002
R51620 S.n17478 S.n17470 0.002
R51621 S.n16944 S.n16937 0.002
R51622 S.n16576 S.n16568 0.002
R51623 S.n16026 S.n16019 0.002
R51624 S.n15652 S.n15644 0.002
R51625 S.n14715 S.n14714 0.002
R51626 S.n22528 S.n22520 0.002
R51627 S.n22115 S.n22108 0.002
R51628 S.n21505 S.n21497 0.002
R51629 S.n21837 S.n21830 0.002
R51630 S.n20682 S.n20674 0.002
R51631 S.n21027 S.n21020 0.002
R51632 S.n20071 S.n20063 0.002
R51633 S.n19623 S.n19616 0.002
R51634 S.n19217 S.n19209 0.002
R51635 S.n18751 S.n18744 0.002
R51636 S.n18351 S.n18343 0.002
R51637 S.n17868 S.n17861 0.002
R51638 S.n17462 S.n17454 0.002
R51639 S.n16959 S.n16952 0.002
R51640 S.n16560 S.n16552 0.002
R51641 S.n16041 S.n16034 0.002
R51642 S.n15636 S.n15628 0.002
R51643 S.n15097 S.n15090 0.002
R51644 S.n14699 S.n14691 0.002
R51645 S.n13740 S.n13739 0.002
R51646 S.n22512 S.n22504 0.002
R51647 S.n22130 S.n22123 0.002
R51648 S.n21489 S.n21481 0.002
R51649 S.n21822 S.n21815 0.002
R51650 S.n20666 S.n20658 0.002
R51651 S.n21012 S.n21005 0.002
R51652 S.n20055 S.n20047 0.002
R51653 S.n19638 S.n19631 0.002
R51654 S.n19201 S.n19193 0.002
R51655 S.n18766 S.n18759 0.002
R51656 S.n18335 S.n18327 0.002
R51657 S.n17883 S.n17876 0.002
R51658 S.n17446 S.n17438 0.002
R51659 S.n16974 S.n16967 0.002
R51660 S.n16544 S.n16536 0.002
R51661 S.n16056 S.n16049 0.002
R51662 S.n15620 S.n15612 0.002
R51663 S.n15112 S.n15105 0.002
R51664 S.n14683 S.n14675 0.002
R51665 S.n14159 S.n14152 0.002
R51666 S.n13724 S.n13716 0.002
R51667 S.n12752 S.n12751 0.002
R51668 S.n22496 S.n22488 0.002
R51669 S.n22145 S.n22138 0.002
R51670 S.n21473 S.n21465 0.002
R51671 S.n21807 S.n21800 0.002
R51672 S.n20650 S.n20642 0.002
R51673 S.n20997 S.n20990 0.002
R51674 S.n20039 S.n20031 0.002
R51675 S.n19653 S.n19646 0.002
R51676 S.n19185 S.n19177 0.002
R51677 S.n18781 S.n18774 0.002
R51678 S.n18319 S.n18311 0.002
R51679 S.n17898 S.n17891 0.002
R51680 S.n17430 S.n17422 0.002
R51681 S.n16989 S.n16982 0.002
R51682 S.n16528 S.n16520 0.002
R51683 S.n16071 S.n16064 0.002
R51684 S.n15604 S.n15596 0.002
R51685 S.n15127 S.n15120 0.002
R51686 S.n14667 S.n14659 0.002
R51687 S.n14174 S.n14167 0.002
R51688 S.n13708 S.n13700 0.002
R51689 S.n13195 S.n13188 0.002
R51690 S.n12736 S.n12728 0.002
R51691 S.n11742 S.n11741 0.002
R51692 S.n22480 S.n22472 0.002
R51693 S.n22160 S.n22153 0.002
R51694 S.n21457 S.n21449 0.002
R51695 S.n21792 S.n21785 0.002
R51696 S.n20634 S.n20626 0.002
R51697 S.n20982 S.n20975 0.002
R51698 S.n20023 S.n20015 0.002
R51699 S.n19668 S.n19661 0.002
R51700 S.n19169 S.n19161 0.002
R51701 S.n18796 S.n18789 0.002
R51702 S.n18303 S.n18295 0.002
R51703 S.n17913 S.n17906 0.002
R51704 S.n17414 S.n17406 0.002
R51705 S.n17004 S.n16997 0.002
R51706 S.n16512 S.n16504 0.002
R51707 S.n16086 S.n16079 0.002
R51708 S.n15588 S.n15580 0.002
R51709 S.n15142 S.n15135 0.002
R51710 S.n14651 S.n14643 0.002
R51711 S.n14189 S.n14182 0.002
R51712 S.n13692 S.n13684 0.002
R51713 S.n13210 S.n13203 0.002
R51714 S.n12720 S.n12712 0.002
R51715 S.n12222 S.n12215 0.002
R51716 S.n11726 S.n11718 0.002
R51717 S.n10719 S.n10718 0.002
R51718 S.n22464 S.n22456 0.002
R51719 S.n22175 S.n22168 0.002
R51720 S.n21441 S.n21433 0.002
R51721 S.n21777 S.n21770 0.002
R51722 S.n20618 S.n20610 0.002
R51723 S.n20967 S.n20960 0.002
R51724 S.n20007 S.n19999 0.002
R51725 S.n19683 S.n19676 0.002
R51726 S.n19153 S.n19145 0.002
R51727 S.n18811 S.n18804 0.002
R51728 S.n18287 S.n18279 0.002
R51729 S.n17928 S.n17921 0.002
R51730 S.n17398 S.n17390 0.002
R51731 S.n17019 S.n17012 0.002
R51732 S.n16496 S.n16488 0.002
R51733 S.n16101 S.n16094 0.002
R51734 S.n15572 S.n15564 0.002
R51735 S.n15157 S.n15150 0.002
R51736 S.n14635 S.n14627 0.002
R51737 S.n14204 S.n14197 0.002
R51738 S.n13676 S.n13668 0.002
R51739 S.n13225 S.n13218 0.002
R51740 S.n12704 S.n12696 0.002
R51741 S.n12237 S.n12230 0.002
R51742 S.n11710 S.n11702 0.002
R51743 S.n11223 S.n11216 0.002
R51744 S.n10703 S.n10695 0.002
R51745 S.n9674 S.n9673 0.002
R51746 S.n22448 S.n22440 0.002
R51747 S.n22190 S.n22183 0.002
R51748 S.n21425 S.n21417 0.002
R51749 S.n21762 S.n21755 0.002
R51750 S.n20602 S.n20594 0.002
R51751 S.n20952 S.n20945 0.002
R51752 S.n19991 S.n19983 0.002
R51753 S.n19698 S.n19691 0.002
R51754 S.n19137 S.n19129 0.002
R51755 S.n18826 S.n18819 0.002
R51756 S.n18271 S.n18263 0.002
R51757 S.n17943 S.n17936 0.002
R51758 S.n17382 S.n17374 0.002
R51759 S.n17034 S.n17027 0.002
R51760 S.n16480 S.n16472 0.002
R51761 S.n16116 S.n16109 0.002
R51762 S.n15556 S.n15548 0.002
R51763 S.n15172 S.n15165 0.002
R51764 S.n14619 S.n14611 0.002
R51765 S.n14219 S.n14212 0.002
R51766 S.n13660 S.n13652 0.002
R51767 S.n13240 S.n13233 0.002
R51768 S.n12688 S.n12680 0.002
R51769 S.n12252 S.n12245 0.002
R51770 S.n11694 S.n11686 0.002
R51771 S.n11238 S.n11231 0.002
R51772 S.n10687 S.n10679 0.002
R51773 S.n10215 S.n10208 0.002
R51774 S.n9658 S.n9650 0.002
R51775 S.n8616 S.n8615 0.002
R51776 S.n22432 S.n22424 0.002
R51777 S.n22205 S.n22198 0.002
R51778 S.n21409 S.n21401 0.002
R51779 S.n21747 S.n21740 0.002
R51780 S.n20586 S.n20578 0.002
R51781 S.n20937 S.n20930 0.002
R51782 S.n19975 S.n19967 0.002
R51783 S.n19713 S.n19706 0.002
R51784 S.n19121 S.n19113 0.002
R51785 S.n18841 S.n18834 0.002
R51786 S.n18255 S.n18247 0.002
R51787 S.n17958 S.n17951 0.002
R51788 S.n17366 S.n17358 0.002
R51789 S.n17049 S.n17042 0.002
R51790 S.n16464 S.n16456 0.002
R51791 S.n16131 S.n16124 0.002
R51792 S.n15540 S.n15532 0.002
R51793 S.n15187 S.n15180 0.002
R51794 S.n14603 S.n14595 0.002
R51795 S.n14234 S.n14227 0.002
R51796 S.n13644 S.n13636 0.002
R51797 S.n13255 S.n13248 0.002
R51798 S.n12672 S.n12664 0.002
R51799 S.n12267 S.n12260 0.002
R51800 S.n11678 S.n11670 0.002
R51801 S.n11253 S.n11246 0.002
R51802 S.n10671 S.n10663 0.002
R51803 S.n10230 S.n10223 0.002
R51804 S.n9642 S.n9634 0.002
R51805 S.n9181 S.n9174 0.002
R51806 S.n8600 S.n8592 0.002
R51807 S.n7536 S.n7535 0.002
R51808 S.n22416 S.n22408 0.002
R51809 S.n22220 S.n22213 0.002
R51810 S.n21393 S.n21385 0.002
R51811 S.n21732 S.n21725 0.002
R51812 S.n20570 S.n20562 0.002
R51813 S.n20922 S.n20915 0.002
R51814 S.n19959 S.n19951 0.002
R51815 S.n19728 S.n19721 0.002
R51816 S.n19105 S.n19097 0.002
R51817 S.n18856 S.n18849 0.002
R51818 S.n18239 S.n18231 0.002
R51819 S.n17973 S.n17966 0.002
R51820 S.n17350 S.n17342 0.002
R51821 S.n17064 S.n17057 0.002
R51822 S.n16448 S.n16440 0.002
R51823 S.n16146 S.n16139 0.002
R51824 S.n15524 S.n15516 0.002
R51825 S.n15202 S.n15195 0.002
R51826 S.n14587 S.n14579 0.002
R51827 S.n14249 S.n14242 0.002
R51828 S.n13628 S.n13620 0.002
R51829 S.n13270 S.n13263 0.002
R51830 S.n12656 S.n12648 0.002
R51831 S.n12282 S.n12275 0.002
R51832 S.n11662 S.n11654 0.002
R51833 S.n11268 S.n11261 0.002
R51834 S.n10655 S.n10647 0.002
R51835 S.n10245 S.n10238 0.002
R51836 S.n9626 S.n9618 0.002
R51837 S.n9196 S.n9189 0.002
R51838 S.n8584 S.n8576 0.002
R51839 S.n8138 S.n8131 0.002
R51840 S.n7520 S.n7512 0.002
R51841 S.n6443 S.n6442 0.002
R51842 S.n22400 S.n22392 0.002
R51843 S.n22235 S.n22228 0.002
R51844 S.n21377 S.n21369 0.002
R51845 S.n21717 S.n21710 0.002
R51846 S.n20554 S.n20546 0.002
R51847 S.n20907 S.n20900 0.002
R51848 S.n19943 S.n19935 0.002
R51849 S.n19743 S.n19736 0.002
R51850 S.n19089 S.n19081 0.002
R51851 S.n18871 S.n18864 0.002
R51852 S.n18223 S.n18215 0.002
R51853 S.n17988 S.n17981 0.002
R51854 S.n17334 S.n17326 0.002
R51855 S.n17079 S.n17072 0.002
R51856 S.n16432 S.n16424 0.002
R51857 S.n16161 S.n16154 0.002
R51858 S.n15508 S.n15500 0.002
R51859 S.n15217 S.n15210 0.002
R51860 S.n14571 S.n14563 0.002
R51861 S.n14264 S.n14257 0.002
R51862 S.n13612 S.n13604 0.002
R51863 S.n13285 S.n13278 0.002
R51864 S.n12640 S.n12632 0.002
R51865 S.n12297 S.n12290 0.002
R51866 S.n11646 S.n11638 0.002
R51867 S.n11283 S.n11276 0.002
R51868 S.n10639 S.n10631 0.002
R51869 S.n10260 S.n10253 0.002
R51870 S.n9610 S.n9602 0.002
R51871 S.n9211 S.n9204 0.002
R51872 S.n8568 S.n8560 0.002
R51873 S.n8153 S.n8146 0.002
R51874 S.n7504 S.n7496 0.002
R51875 S.n7069 S.n7062 0.002
R51876 S.n6427 S.n6419 0.002
R51877 S.n5327 S.n5326 0.002
R51878 S.n22384 S.n22376 0.002
R51879 S.n22250 S.n22243 0.002
R51880 S.n21361 S.n21353 0.002
R51881 S.n21702 S.n21695 0.002
R51882 S.n20538 S.n20530 0.002
R51883 S.n20892 S.n20885 0.002
R51884 S.n19927 S.n19919 0.002
R51885 S.n19758 S.n19751 0.002
R51886 S.n19073 S.n19065 0.002
R51887 S.n18886 S.n18879 0.002
R51888 S.n18207 S.n18199 0.002
R51889 S.n18003 S.n17996 0.002
R51890 S.n17318 S.n17310 0.002
R51891 S.n17094 S.n17087 0.002
R51892 S.n16416 S.n16408 0.002
R51893 S.n16176 S.n16169 0.002
R51894 S.n15492 S.n15484 0.002
R51895 S.n15232 S.n15225 0.002
R51896 S.n14555 S.n14547 0.002
R51897 S.n14279 S.n14272 0.002
R51898 S.n13596 S.n13588 0.002
R51899 S.n13300 S.n13293 0.002
R51900 S.n12624 S.n12616 0.002
R51901 S.n12312 S.n12305 0.002
R51902 S.n11630 S.n11622 0.002
R51903 S.n11298 S.n11291 0.002
R51904 S.n10623 S.n10615 0.002
R51905 S.n10275 S.n10268 0.002
R51906 S.n9594 S.n9586 0.002
R51907 S.n9229 S.n9222 0.002
R51908 S.n8552 S.n8544 0.002
R51909 S.n8168 S.n8161 0.002
R51910 S.n7488 S.n7480 0.002
R51911 S.n7084 S.n7077 0.002
R51912 S.n6411 S.n6403 0.002
R51913 S.n5991 S.n5984 0.002
R51914 S.n5311 S.n5303 0.002
R51915 S.n4198 S.n4197 0.002
R51916 S.n22672 S.n22266 0.002
R51917 S.n22675 S.n22258 0.002
R51918 S.n21685 S.n21672 0.002
R51919 S.n21687 S.n21664 0.002
R51920 S.n20522 S.n20515 0.002
R51921 S.n20877 S.n20869 0.002
R51922 S.n19911 S.n19904 0.002
R51923 S.n19774 S.n19766 0.002
R51924 S.n19057 S.n19050 0.002
R51925 S.n18902 S.n18894 0.002
R51926 S.n18191 S.n18184 0.002
R51927 S.n18019 S.n18011 0.002
R51928 S.n17302 S.n17295 0.002
R51929 S.n17110 S.n17102 0.002
R51930 S.n16400 S.n16393 0.002
R51931 S.n16192 S.n16184 0.002
R51932 S.n15476 S.n15469 0.002
R51933 S.n15248 S.n15240 0.002
R51934 S.n14539 S.n14532 0.002
R51935 S.n14295 S.n14287 0.002
R51936 S.n13580 S.n13573 0.002
R51937 S.n13316 S.n13308 0.002
R51938 S.n12608 S.n12601 0.002
R51939 S.n12328 S.n12320 0.002
R51940 S.n11614 S.n11607 0.002
R51941 S.n11314 S.n11306 0.002
R51942 S.n10607 S.n10600 0.002
R51943 S.n10291 S.n10283 0.002
R51944 S.n9578 S.n9571 0.002
R51945 S.n9242 S.n9234 0.002
R51946 S.n8536 S.n8529 0.002
R51947 S.n8184 S.n8176 0.002
R51948 S.n7472 S.n7465 0.002
R51949 S.n7100 S.n7092 0.002
R51950 S.n6395 S.n6388 0.002
R51951 S.n6007 S.n5999 0.002
R51952 S.n5295 S.n5288 0.002
R51953 S.n4887 S.n4879 0.002
R51954 S.n4182 S.n4175 0.002
R51955 S.n3057 S.n3056 0.002
R51956 S.n22368 S.n22359 0.002
R51957 S.n22694 S.n22683 0.002
R51958 S.n21654 S.n21277 0.002
R51959 S.n21656 S.n21269 0.002
R51960 S.n20507 S.n20500 0.002
R51961 S.n20861 S.n20853 0.002
R51962 S.n19896 S.n19889 0.002
R51963 S.n19790 S.n19782 0.002
R51964 S.n19042 S.n19035 0.002
R51965 S.n18918 S.n18910 0.002
R51966 S.n18176 S.n18169 0.002
R51967 S.n18035 S.n18027 0.002
R51968 S.n17287 S.n17280 0.002
R51969 S.n17126 S.n17118 0.002
R51970 S.n16385 S.n16378 0.002
R51971 S.n16208 S.n16200 0.002
R51972 S.n15461 S.n15454 0.002
R51973 S.n15264 S.n15256 0.002
R51974 S.n14524 S.n14517 0.002
R51975 S.n14311 S.n14303 0.002
R51976 S.n13565 S.n13558 0.002
R51977 S.n13332 S.n13324 0.002
R51978 S.n12593 S.n12586 0.002
R51979 S.n12344 S.n12336 0.002
R51980 S.n11599 S.n11592 0.002
R51981 S.n11330 S.n11322 0.002
R51982 S.n10592 S.n10585 0.002
R51983 S.n10307 S.n10299 0.002
R51984 S.n9563 S.n9556 0.002
R51985 S.n9258 S.n9250 0.002
R51986 S.n8521 S.n8514 0.002
R51987 S.n8200 S.n8192 0.002
R51988 S.n7457 S.n7450 0.002
R51989 S.n7116 S.n7108 0.002
R51990 S.n6380 S.n6373 0.002
R51991 S.n6023 S.n6015 0.002
R51992 S.n5280 S.n5273 0.002
R51993 S.n4903 S.n4895 0.002
R51994 S.n4167 S.n4160 0.002
R51995 S.n3775 S.n3767 0.002
R51996 S.n3041 S.n3034 0.002
R51997 S.n1899 S.n1898 0.002
R51998 S.n21314 S.n21303 0.002
R51999 S.n21217 S.n21202 0.002
R52000 S.n20491 S.n20480 0.002
R52001 S.n20398 S.n20383 0.002
R52002 S.n19880 S.n19869 0.002
R52003 S.n20271 S.n20256 0.002
R52004 S.n19026 S.n19015 0.002
R52005 S.n19403 S.n19388 0.002
R52006 S.n18160 S.n18149 0.002
R52007 S.n18516 S.n18501 0.002
R52008 S.n17271 S.n17260 0.002
R52009 S.n17616 S.n17601 0.002
R52010 S.n16369 S.n16358 0.002
R52011 S.n16693 S.n16678 0.002
R52012 S.n15445 S.n15434 0.002
R52013 S.n15758 S.n15743 0.002
R52014 S.n14508 S.n14497 0.002
R52015 S.n14800 S.n14785 0.002
R52016 S.n13549 S.n13538 0.002
R52017 S.n13830 S.n13815 0.002
R52018 S.n12577 S.n12566 0.002
R52019 S.n12837 S.n12822 0.002
R52020 S.n11583 S.n11572 0.002
R52021 S.n11832 S.n11817 0.002
R52022 S.n10576 S.n10565 0.002
R52023 S.n10804 S.n10789 0.002
R52024 S.n9547 S.n9536 0.002
R52025 S.n9764 S.n9749 0.002
R52026 S.n8505 S.n8494 0.002
R52027 S.n8701 S.n8686 0.002
R52028 S.n7441 S.n7430 0.002
R52029 S.n7626 S.n7611 0.002
R52030 S.n6364 S.n6353 0.002
R52031 S.n6528 S.n6513 0.002
R52032 S.n5264 S.n5253 0.002
R52033 S.n5417 S.n5402 0.002
R52034 S.n4151 S.n4140 0.002
R52035 S.n4283 S.n4268 0.002
R52036 S.n3025 S.n3014 0.002
R52037 S.n3146 S.n3132 0.002
R52038 S.n1865 S.n1853 0.002
R52039 S.n17169 S.n17158 0.002
R52040 S.n17765 S.n17750 0.002
R52041 S.n16269 S.n16258 0.002
R52042 S.n16838 S.n16823 0.002
R52043 S.n15345 S.n15334 0.002
R52044 S.n15903 S.n15888 0.002
R52045 S.n14408 S.n14397 0.002
R52046 S.n14945 S.n14930 0.002
R52047 S.n13449 S.n13438 0.002
R52048 S.n13975 S.n13960 0.002
R52049 S.n12477 S.n12466 0.002
R52050 S.n12982 S.n12967 0.002
R52051 S.n11483 S.n11472 0.002
R52052 S.n11977 S.n11962 0.002
R52053 S.n10476 S.n10465 0.002
R52054 S.n10949 S.n10934 0.002
R52055 S.n9447 S.n9436 0.002
R52056 S.n9909 S.n9894 0.002
R52057 S.n8405 S.n8394 0.002
R52058 S.n8846 S.n8831 0.002
R52059 S.n7341 S.n7330 0.002
R52060 S.n7771 S.n7756 0.002
R52061 S.n6264 S.n6253 0.002
R52062 S.n6673 S.n6658 0.002
R52063 S.n5164 S.n5153 0.002
R52064 S.n5563 S.n5548 0.002
R52065 S.n4052 S.n4041 0.002
R52066 S.n4428 S.n4413 0.002
R52067 S.n2925 S.n2914 0.002
R52068 S.n3290 S.n3276 0.002
R52069 S.n1757 S.n1745 0.002
R52070 S.n2107 S.n2106 0.002
R52071 S.n743 S.n742 0.002
R52072 S.n726 S.n725 0.002
R52073 S.n15307 S.n15296 0.002
R52074 S.n15968 S.n15953 0.002
R52075 S.n14372 S.n14361 0.002
R52076 S.n15006 S.n14991 0.002
R52077 S.n13413 S.n13402 0.002
R52078 S.n14036 S.n14021 0.002
R52079 S.n12441 S.n12430 0.002
R52080 S.n13043 S.n13028 0.002
R52081 S.n11447 S.n11436 0.002
R52082 S.n12038 S.n12023 0.002
R52083 S.n10440 S.n10429 0.002
R52084 S.n11010 S.n10995 0.002
R52085 S.n9411 S.n9400 0.002
R52086 S.n9970 S.n9955 0.002
R52087 S.n8369 S.n8358 0.002
R52088 S.n8907 S.n8892 0.002
R52089 S.n7305 S.n7294 0.002
R52090 S.n7832 S.n7817 0.002
R52091 S.n6228 S.n6217 0.002
R52092 S.n6734 S.n6719 0.002
R52093 S.n5128 S.n5117 0.002
R52094 S.n5624 S.n5609 0.002
R52095 S.n4016 S.n4005 0.002
R52096 S.n4489 S.n4474 0.002
R52097 S.n2889 S.n2878 0.002
R52098 S.n3350 S.n3336 0.002
R52099 S.n1720 S.n1708 0.002
R52100 S.n2166 S.n2165 0.002
R52101 S.n708 S.n707 0.002
R52102 S.n691 S.n690 0.002
R52103 S.n13375 S.n13364 0.002
R52104 S.n14101 S.n14086 0.002
R52105 S.n12405 S.n12394 0.002
R52106 S.n13104 S.n13089 0.002
R52107 S.n11411 S.n11400 0.002
R52108 S.n12099 S.n12084 0.002
R52109 S.n10404 S.n10393 0.002
R52110 S.n11071 S.n11056 0.002
R52111 S.n9375 S.n9364 0.002
R52112 S.n10031 S.n10016 0.002
R52113 S.n8333 S.n8322 0.002
R52114 S.n8968 S.n8953 0.002
R52115 S.n7269 S.n7258 0.002
R52116 S.n7893 S.n7878 0.002
R52117 S.n6192 S.n6181 0.002
R52118 S.n6795 S.n6780 0.002
R52119 S.n5092 S.n5081 0.002
R52120 S.n5685 S.n5670 0.002
R52121 S.n3980 S.n3969 0.002
R52122 S.n4550 S.n4535 0.002
R52123 S.n2853 S.n2842 0.002
R52124 S.n3410 S.n3396 0.002
R52125 S.n1683 S.n1671 0.002
R52126 S.n2225 S.n2224 0.002
R52127 S.n673 S.n672 0.002
R52128 S.n656 S.n655 0.002
R52129 S.n11373 S.n11362 0.002
R52130 S.n12164 S.n12149 0.002
R52131 S.n10368 S.n10357 0.002
R52132 S.n11132 S.n11117 0.002
R52133 S.n9339 S.n9328 0.002
R52134 S.n10092 S.n10077 0.002
R52135 S.n8297 S.n8286 0.002
R52136 S.n9029 S.n9014 0.002
R52137 S.n7233 S.n7222 0.002
R52138 S.n7954 S.n7939 0.002
R52139 S.n6156 S.n6145 0.002
R52140 S.n6856 S.n6841 0.002
R52141 S.n5056 S.n5045 0.002
R52142 S.n5746 S.n5731 0.002
R52143 S.n3944 S.n3933 0.002
R52144 S.n4611 S.n4596 0.002
R52145 S.n2817 S.n2806 0.002
R52146 S.n3470 S.n3456 0.002
R52147 S.n1646 S.n1634 0.002
R52148 S.n2284 S.n2283 0.002
R52149 S.n638 S.n637 0.002
R52150 S.n621 S.n620 0.002
R52151 S.n9301 S.n9290 0.002
R52152 S.n10157 S.n10142 0.002
R52153 S.n8261 S.n8250 0.002
R52154 S.n9090 S.n9075 0.002
R52155 S.n7197 S.n7186 0.002
R52156 S.n8015 S.n8000 0.002
R52157 S.n6120 S.n6109 0.002
R52158 S.n6917 S.n6902 0.002
R52159 S.n5020 S.n5009 0.002
R52160 S.n5807 S.n5792 0.002
R52161 S.n3908 S.n3897 0.002
R52162 S.n4672 S.n4657 0.002
R52163 S.n2781 S.n2770 0.002
R52164 S.n3530 S.n3516 0.002
R52165 S.n1609 S.n1597 0.002
R52166 S.n2343 S.n2342 0.002
R52167 S.n603 S.n602 0.002
R52168 S.n586 S.n585 0.002
R52169 S.n7159 S.n7148 0.002
R52170 S.n8080 S.n8065 0.002
R52171 S.n6084 S.n6073 0.002
R52172 S.n6978 S.n6963 0.002
R52173 S.n4984 S.n4973 0.002
R52174 S.n5868 S.n5853 0.002
R52175 S.n3872 S.n3861 0.002
R52176 S.n4733 S.n4718 0.002
R52177 S.n2745 S.n2734 0.002
R52178 S.n3590 S.n3576 0.002
R52179 S.n1572 S.n1560 0.002
R52180 S.n2402 S.n2401 0.002
R52181 S.n568 S.n567 0.002
R52182 S.n551 S.n550 0.002
R52183 S.n4946 S.n4935 0.002
R52184 S.n5933 S.n5918 0.002
R52185 S.n3836 S.n3825 0.002
R52186 S.n4794 S.n4779 0.002
R52187 S.n2709 S.n2698 0.002
R52188 S.n3650 S.n3636 0.002
R52189 S.n1535 S.n1523 0.002
R52190 S.n2461 S.n2460 0.002
R52191 S.n533 S.n532 0.002
R52192 S.n516 S.n515 0.002
R52193 S.n2671 S.n2660 0.002
R52194 S.n3714 S.n3700 0.002
R52195 S.n1498 S.n1486 0.002
R52196 S.n2520 S.n2519 0.002
R52197 S.n498 S.n497 0.002
R52198 S.n481 S.n480 0.002
R52199 S.n463 S.n462 0.002
R52200 S.n447 S.n446 0.002
R52201 S.n22307 S.n22294 0.002
R52202 S.n22765 S.n22764 0.002
R52203 S.n21328 S.n21327 0.002
R52204 S.n21149 S.n21148 0.002
R52205 S.n21638 S.n21629 0.002
R52206 S.n20818 S.n20806 0.002
R52207 S.n21152 S.n21151 0.002
R52208 S.n1337 S.n1322 0.002
R52209 S.n864 S.n863 0.002
R52210 S.n3729 S.n3728 0.002
R52211 S.n43 S.n42 0.002
R52212 S.t41 S.n22992 0.002
R52213 S.t41 S.n23007 0.002
R52214 S.n22741 S.n22723 0.002
R52215 S.n18483 S.n18466 0.002
R52216 S.n16660 S.n16643 0.002
R52217 S.n14767 S.n14750 0.002
R52218 S.n12804 S.n12787 0.002
R52219 S.n10771 S.n10754 0.002
R52220 S.n8668 S.n8651 0.002
R52221 S.n6495 S.n6478 0.002
R52222 S.n4250 S.n4233 0.002
R52223 S.n1954 S.n1939 0.002
R52224 S.n1183 S.n1182 0.002
R52225 S.n22713 S.n22712 0.002
R52226 S.n21345 S.n21344 0.002
R52227 S.n21261 S.n21260 0.002
R52228 S.n20835 S.n20834 0.002
R52229 S.n20845 S.n20844 0.002
R52230 S.n20200 S.n20199 0.002
R52231 S.n20210 S.n20209 0.002
R52232 S.n19330 S.n19329 0.002
R52233 S.n19340 S.n19339 0.002
R52234 S.n18448 S.n18447 0.002
R52235 S.n18458 S.n18457 0.002
R52236 S.n17543 S.n17542 0.002
R52237 S.n17553 S.n17552 0.002
R52238 S.n16625 S.n16624 0.002
R52239 S.n16635 S.n16634 0.002
R52240 S.n15685 S.n15684 0.002
R52241 S.n15695 S.n15694 0.002
R52242 S.n14732 S.n14731 0.002
R52243 S.n14742 S.n14741 0.002
R52244 S.n13757 S.n13756 0.002
R52245 S.n13767 S.n13766 0.002
R52246 S.n12769 S.n12768 0.002
R52247 S.n12779 S.n12778 0.002
R52248 S.n11759 S.n11758 0.002
R52249 S.n11769 S.n11768 0.002
R52250 S.n10736 S.n10735 0.002
R52251 S.n10746 S.n10745 0.002
R52252 S.n9691 S.n9690 0.002
R52253 S.n9701 S.n9700 0.002
R52254 S.n8633 S.n8632 0.002
R52255 S.n8643 S.n8642 0.002
R52256 S.n7553 S.n7552 0.002
R52257 S.n7563 S.n7562 0.002
R52258 S.n6460 S.n6459 0.002
R52259 S.n6470 S.n6469 0.002
R52260 S.n5344 S.n5343 0.002
R52261 S.n5354 S.n5353 0.002
R52262 S.n4215 S.n4214 0.002
R52263 S.n4225 S.n4224 0.002
R52264 S.n3074 S.n3073 0.002
R52265 S.n3084 S.n3083 0.002
R52266 S.n1882 S.n1881 0.002
R52267 S.n21242 S.n21241 0.002
R52268 S.n20366 S.n20365 0.002
R52269 S.n20295 S.n20294 0.002
R52270 S.n19423 S.n19422 0.002
R52271 S.n18536 S.n18535 0.002
R52272 S.n17636 S.n17635 0.002
R52273 S.n16713 S.n16712 0.002
R52274 S.n15778 S.n15777 0.002
R52275 S.n14820 S.n14819 0.002
R52276 S.n13850 S.n13849 0.002
R52277 S.n12857 S.n12856 0.002
R52278 S.n11852 S.n11851 0.002
R52279 S.n10824 S.n10823 0.002
R52280 S.n9784 S.n9783 0.002
R52281 S.n8721 S.n8720 0.002
R52282 S.n7646 S.n7645 0.002
R52283 S.n6548 S.n6547 0.002
R52284 S.n5438 S.n5437 0.002
R52285 S.n4303 S.n4302 0.002
R52286 S.n3166 S.n3165 0.002
R52287 S.n22351 S.n22350 0.002
R52288 S.n22656 S.n22647 0.002
R52289 S.n20183 S.n20174 0.002
R52290 S.n20794 S.n20793 0.002
R52291 S.n21617 S.n21616 0.002
R52292 S.n22640 S.n22639 0.002
R52293 S.n19313 S.n19304 0.002
R52294 S.n20167 S.n20166 0.002
R52295 S.n20778 S.n20777 0.002
R52296 S.n21601 S.n21600 0.002
R52297 S.n22624 S.n22623 0.002
R52298 S.n18431 S.n18422 0.002
R52299 S.n19297 S.n19296 0.002
R52300 S.n20151 S.n20150 0.002
R52301 S.n20762 S.n20761 0.002
R52302 S.n21585 S.n21584 0.002
R52303 S.n22608 S.n22607 0.002
R52304 S.n17526 S.n17517 0.002
R52305 S.n18415 S.n18414 0.002
R52306 S.n19281 S.n19280 0.002
R52307 S.n20135 S.n20134 0.002
R52308 S.n20746 S.n20745 0.002
R52309 S.n21569 S.n21568 0.002
R52310 S.n22592 S.n22591 0.002
R52311 S.n16608 S.n16599 0.002
R52312 S.n17510 S.n17509 0.002
R52313 S.n18399 S.n18398 0.002
R52314 S.n19265 S.n19264 0.002
R52315 S.n20119 S.n20118 0.002
R52316 S.n20730 S.n20729 0.002
R52317 S.n21553 S.n21552 0.002
R52318 S.n22576 S.n22575 0.002
R52319 S.n15668 S.n15659 0.002
R52320 S.n16592 S.n16591 0.002
R52321 S.n17494 S.n17493 0.002
R52322 S.n18383 S.n18382 0.002
R52323 S.n19249 S.n19248 0.002
R52324 S.n20103 S.n20102 0.002
R52325 S.n20714 S.n20713 0.002
R52326 S.n21537 S.n21536 0.002
R52327 S.n22560 S.n22559 0.002
R52328 S.n14715 S.n14706 0.002
R52329 S.n15652 S.n15651 0.002
R52330 S.n16576 S.n16575 0.002
R52331 S.n17478 S.n17477 0.002
R52332 S.n18367 S.n18366 0.002
R52333 S.n19233 S.n19232 0.002
R52334 S.n20087 S.n20086 0.002
R52335 S.n20698 S.n20697 0.002
R52336 S.n21521 S.n21520 0.002
R52337 S.n22544 S.n22543 0.002
R52338 S.n13740 S.n13731 0.002
R52339 S.n14699 S.n14698 0.002
R52340 S.n15636 S.n15635 0.002
R52341 S.n16560 S.n16559 0.002
R52342 S.n17462 S.n17461 0.002
R52343 S.n18351 S.n18350 0.002
R52344 S.n19217 S.n19216 0.002
R52345 S.n20071 S.n20070 0.002
R52346 S.n20682 S.n20681 0.002
R52347 S.n21505 S.n21504 0.002
R52348 S.n22528 S.n22527 0.002
R52349 S.n12752 S.n12743 0.002
R52350 S.n13724 S.n13723 0.002
R52351 S.n14683 S.n14682 0.002
R52352 S.n15620 S.n15619 0.002
R52353 S.n16544 S.n16543 0.002
R52354 S.n17446 S.n17445 0.002
R52355 S.n18335 S.n18334 0.002
R52356 S.n19201 S.n19200 0.002
R52357 S.n20055 S.n20054 0.002
R52358 S.n20666 S.n20665 0.002
R52359 S.n21489 S.n21488 0.002
R52360 S.n22512 S.n22511 0.002
R52361 S.n11742 S.n11733 0.002
R52362 S.n12736 S.n12735 0.002
R52363 S.n13708 S.n13707 0.002
R52364 S.n14667 S.n14666 0.002
R52365 S.n15604 S.n15603 0.002
R52366 S.n16528 S.n16527 0.002
R52367 S.n17430 S.n17429 0.002
R52368 S.n18319 S.n18318 0.002
R52369 S.n19185 S.n19184 0.002
R52370 S.n20039 S.n20038 0.002
R52371 S.n20650 S.n20649 0.002
R52372 S.n21473 S.n21472 0.002
R52373 S.n22496 S.n22495 0.002
R52374 S.n10719 S.n10710 0.002
R52375 S.n11726 S.n11725 0.002
R52376 S.n12720 S.n12719 0.002
R52377 S.n13692 S.n13691 0.002
R52378 S.n14651 S.n14650 0.002
R52379 S.n15588 S.n15587 0.002
R52380 S.n16512 S.n16511 0.002
R52381 S.n17414 S.n17413 0.002
R52382 S.n18303 S.n18302 0.002
R52383 S.n19169 S.n19168 0.002
R52384 S.n20023 S.n20022 0.002
R52385 S.n20634 S.n20633 0.002
R52386 S.n21457 S.n21456 0.002
R52387 S.n22480 S.n22479 0.002
R52388 S.n9674 S.n9665 0.002
R52389 S.n10703 S.n10702 0.002
R52390 S.n11710 S.n11709 0.002
R52391 S.n12704 S.n12703 0.002
R52392 S.n13676 S.n13675 0.002
R52393 S.n14635 S.n14634 0.002
R52394 S.n15572 S.n15571 0.002
R52395 S.n16496 S.n16495 0.002
R52396 S.n17398 S.n17397 0.002
R52397 S.n18287 S.n18286 0.002
R52398 S.n19153 S.n19152 0.002
R52399 S.n20007 S.n20006 0.002
R52400 S.n20618 S.n20617 0.002
R52401 S.n21441 S.n21440 0.002
R52402 S.n22464 S.n22463 0.002
R52403 S.n8616 S.n8607 0.002
R52404 S.n9658 S.n9657 0.002
R52405 S.n10687 S.n10686 0.002
R52406 S.n11694 S.n11693 0.002
R52407 S.n12688 S.n12687 0.002
R52408 S.n13660 S.n13659 0.002
R52409 S.n14619 S.n14618 0.002
R52410 S.n15556 S.n15555 0.002
R52411 S.n16480 S.n16479 0.002
R52412 S.n17382 S.n17381 0.002
R52413 S.n18271 S.n18270 0.002
R52414 S.n19137 S.n19136 0.002
R52415 S.n19991 S.n19990 0.002
R52416 S.n20602 S.n20601 0.002
R52417 S.n21425 S.n21424 0.002
R52418 S.n22448 S.n22447 0.002
R52419 S.n7536 S.n7527 0.002
R52420 S.n8600 S.n8599 0.002
R52421 S.n9642 S.n9641 0.002
R52422 S.n10671 S.n10670 0.002
R52423 S.n11678 S.n11677 0.002
R52424 S.n12672 S.n12671 0.002
R52425 S.n13644 S.n13643 0.002
R52426 S.n14603 S.n14602 0.002
R52427 S.n15540 S.n15539 0.002
R52428 S.n16464 S.n16463 0.002
R52429 S.n17366 S.n17365 0.002
R52430 S.n18255 S.n18254 0.002
R52431 S.n19121 S.n19120 0.002
R52432 S.n19975 S.n19974 0.002
R52433 S.n20586 S.n20585 0.002
R52434 S.n21409 S.n21408 0.002
R52435 S.n22432 S.n22431 0.002
R52436 S.n6443 S.n6434 0.002
R52437 S.n7520 S.n7519 0.002
R52438 S.n8584 S.n8583 0.002
R52439 S.n9626 S.n9625 0.002
R52440 S.n10655 S.n10654 0.002
R52441 S.n11662 S.n11661 0.002
R52442 S.n12656 S.n12655 0.002
R52443 S.n13628 S.n13627 0.002
R52444 S.n14587 S.n14586 0.002
R52445 S.n15524 S.n15523 0.002
R52446 S.n16448 S.n16447 0.002
R52447 S.n17350 S.n17349 0.002
R52448 S.n18239 S.n18238 0.002
R52449 S.n19105 S.n19104 0.002
R52450 S.n19959 S.n19958 0.002
R52451 S.n20570 S.n20569 0.002
R52452 S.n21393 S.n21392 0.002
R52453 S.n22416 S.n22415 0.002
R52454 S.n5327 S.n5318 0.002
R52455 S.n6427 S.n6426 0.002
R52456 S.n7504 S.n7503 0.002
R52457 S.n8568 S.n8567 0.002
R52458 S.n9610 S.n9609 0.002
R52459 S.n10639 S.n10638 0.002
R52460 S.n11646 S.n11645 0.002
R52461 S.n12640 S.n12639 0.002
R52462 S.n13612 S.n13611 0.002
R52463 S.n14571 S.n14570 0.002
R52464 S.n15508 S.n15507 0.002
R52465 S.n16432 S.n16431 0.002
R52466 S.n17334 S.n17333 0.002
R52467 S.n18223 S.n18222 0.002
R52468 S.n19089 S.n19088 0.002
R52469 S.n19943 S.n19942 0.002
R52470 S.n20554 S.n20553 0.002
R52471 S.n21377 S.n21376 0.002
R52472 S.n22400 S.n22399 0.002
R52473 S.n4198 S.n4189 0.002
R52474 S.n5311 S.n5310 0.002
R52475 S.n6411 S.n6410 0.002
R52476 S.n7488 S.n7487 0.002
R52477 S.n8552 S.n8551 0.002
R52478 S.n9594 S.n9593 0.002
R52479 S.n10623 S.n10622 0.002
R52480 S.n11630 S.n11629 0.002
R52481 S.n12624 S.n12623 0.002
R52482 S.n13596 S.n13595 0.002
R52483 S.n14555 S.n14554 0.002
R52484 S.n15492 S.n15491 0.002
R52485 S.n16416 S.n16415 0.002
R52486 S.n17318 S.n17317 0.002
R52487 S.n18207 S.n18206 0.002
R52488 S.n19073 S.n19072 0.002
R52489 S.n19927 S.n19926 0.002
R52490 S.n20538 S.n20537 0.002
R52491 S.n21361 S.n21360 0.002
R52492 S.n22384 S.n22383 0.002
R52493 S.n3057 S.n3048 0.002
R52494 S.n21686 S.n21685 0.002
R52495 S.n22674 S.n22672 0.002
R52496 S.n1899 S.n1442 0.002
R52497 S.n21655 S.n21654 0.002
R52498 S.n22368 S.n22367 0.002
R52499 S.n22351 S.n22342 0.002
R52500 S.n21345 S.n21336 0.002
R52501 S.n20836 S.n20835 0.002
R52502 S.n20201 S.n20200 0.002
R52503 S.n19331 S.n19330 0.002
R52504 S.n18449 S.n18448 0.002
R52505 S.n17544 S.n17543 0.002
R52506 S.n16626 S.n16625 0.002
R52507 S.n15686 S.n15685 0.002
R52508 S.n14733 S.n14732 0.002
R52509 S.n13758 S.n13757 0.002
R52510 S.n12770 S.n12769 0.002
R52511 S.n11760 S.n11759 0.002
R52512 S.n10737 S.n10736 0.002
R52513 S.n9692 S.n9691 0.002
R52514 S.n8634 S.n8633 0.002
R52515 S.n7554 S.n7553 0.002
R52516 S.n6461 S.n6460 0.002
R52517 S.n5345 S.n5344 0.002
R52518 S.n4216 S.n4215 0.002
R52519 S.n3075 S.n3074 0.002
R52520 S.n1882 S.n1873 0.002
R52521 S.n806 S.n794 0.002
R52522 S.n19839 S.n19838 0.002
R52523 S.n18987 S.n18986 0.002
R52524 S.n18121 S.n18120 0.002
R52525 S.n17232 S.n17231 0.002
R52526 S.n16330 S.n16329 0.002
R52527 S.n15406 S.n15405 0.002
R52528 S.n14469 S.n14468 0.002
R52529 S.n13510 S.n13509 0.002
R52530 S.n12538 S.n12537 0.002
R52531 S.n11544 S.n11543 0.002
R52532 S.n10537 S.n10536 0.002
R52533 S.n9508 S.n9507 0.002
R52534 S.n8466 S.n8465 0.002
R52535 S.n7402 S.n7401 0.002
R52536 S.n6325 S.n6324 0.002
R52537 S.n5225 S.n5224 0.002
R52538 S.n4113 S.n4112 0.002
R52539 S.n2986 S.n2985 0.002
R52540 S.n1823 S.n1822 0.002
R52541 S.n767 S.n750 0.002
R52542 S.n22328 S.n22326 0.002
R52543 S.n22741 S.n22722 0.002
R52544 S.n21314 S.n21302 0.002
R52545 S.n21217 S.n21192 0.002
R52546 S.n20491 S.n20479 0.002
R52547 S.n20398 S.n20373 0.002
R52548 S.n19880 S.n19868 0.002
R52549 S.n20271 S.n20246 0.002
R52550 S.n19026 S.n19014 0.002
R52551 S.n19403 S.n19378 0.002
R52552 S.n18160 S.n18148 0.002
R52553 S.n18516 S.n18491 0.002
R52554 S.n17271 S.n17259 0.002
R52555 S.n17616 S.n17591 0.002
R52556 S.n16369 S.n16357 0.002
R52557 S.n16693 S.n16668 0.002
R52558 S.n15445 S.n15433 0.002
R52559 S.n15758 S.n15733 0.002
R52560 S.n14508 S.n14496 0.002
R52561 S.n14800 S.n14775 0.002
R52562 S.n13549 S.n13537 0.002
R52563 S.n13830 S.n13805 0.002
R52564 S.n12577 S.n12565 0.002
R52565 S.n12837 S.n12812 0.002
R52566 S.n11583 S.n11571 0.002
R52567 S.n11832 S.n11807 0.002
R52568 S.n10576 S.n10564 0.002
R52569 S.n10804 S.n10779 0.002
R52570 S.n9547 S.n9535 0.002
R52571 S.n9764 S.n9739 0.002
R52572 S.n8505 S.n8493 0.002
R52573 S.n8701 S.n8676 0.002
R52574 S.n7441 S.n7429 0.002
R52575 S.n7626 S.n7601 0.002
R52576 S.n6364 S.n6352 0.002
R52577 S.n6528 S.n6503 0.002
R52578 S.n5264 S.n5252 0.002
R52579 S.n5417 S.n5392 0.002
R52580 S.n4151 S.n4139 0.002
R52581 S.n4283 S.n4258 0.002
R52582 S.n3025 S.n3013 0.002
R52583 S.n3146 S.n3122 0.002
R52584 S.n1865 S.n1852 0.002
R52585 S.n1985 S.n1962 0.002
R52586 S.n890 S.n871 0.002
R52587 S.n914 S.n893 0.002
R52588 S.n20238 S.n20217 0.002
R52589 S.n18961 S.n18949 0.002
R52590 S.n19490 S.n19465 0.002
R52591 S.n18096 S.n18084 0.002
R52592 S.n18600 S.n18575 0.002
R52593 S.n17207 S.n17195 0.002
R52594 S.n17700 S.n17675 0.002
R52595 S.n16305 S.n16293 0.002
R52596 S.n16777 S.n16752 0.002
R52597 S.n15381 S.n15369 0.002
R52598 S.n15842 S.n15817 0.002
R52599 S.n14444 S.n14432 0.002
R52600 S.n14884 S.n14859 0.002
R52601 S.n13485 S.n13473 0.002
R52602 S.n13914 S.n13889 0.002
R52603 S.n12513 S.n12501 0.002
R52604 S.n12921 S.n12896 0.002
R52605 S.n11519 S.n11507 0.002
R52606 S.n11916 S.n11891 0.002
R52607 S.n10512 S.n10500 0.002
R52608 S.n10888 S.n10863 0.002
R52609 S.n9483 S.n9471 0.002
R52610 S.n9848 S.n9823 0.002
R52611 S.n8441 S.n8429 0.002
R52612 S.n8785 S.n8760 0.002
R52613 S.n7377 S.n7365 0.002
R52614 S.n7710 S.n7685 0.002
R52615 S.n6300 S.n6288 0.002
R52616 S.n6612 S.n6587 0.002
R52617 S.n5200 S.n5188 0.002
R52618 S.n5502 S.n5477 0.002
R52619 S.n4088 S.n4076 0.002
R52620 S.n4367 S.n4342 0.002
R52621 S.n2961 S.n2949 0.002
R52622 S.n3230 S.n3205 0.002
R52623 S.n1799 S.n1788 0.002
R52624 S.n2079 S.n2058 0.002
R52625 S.n838 S.n826 0.002
R52626 S.n823 S.n413 0.002
R52627 S.n18483 S.n18465 0.002
R52628 S.n17169 S.n17157 0.002
R52629 S.n17765 S.n17740 0.002
R52630 S.n16269 S.n16257 0.002
R52631 S.n16838 S.n16813 0.002
R52632 S.n15345 S.n15333 0.002
R52633 S.n15903 S.n15878 0.002
R52634 S.n14408 S.n14396 0.002
R52635 S.n14945 S.n14920 0.002
R52636 S.n13449 S.n13437 0.002
R52637 S.n13975 S.n13950 0.002
R52638 S.n12477 S.n12465 0.002
R52639 S.n12982 S.n12957 0.002
R52640 S.n11483 S.n11471 0.002
R52641 S.n11977 S.n11952 0.002
R52642 S.n10476 S.n10464 0.002
R52643 S.n10949 S.n10924 0.002
R52644 S.n9447 S.n9435 0.002
R52645 S.n9909 S.n9884 0.002
R52646 S.n8405 S.n8393 0.002
R52647 S.n8846 S.n8821 0.002
R52648 S.n7341 S.n7329 0.002
R52649 S.n7771 S.n7746 0.002
R52650 S.n6264 S.n6252 0.002
R52651 S.n6673 S.n6648 0.002
R52652 S.n5164 S.n5152 0.002
R52653 S.n5563 S.n5538 0.002
R52654 S.n4052 S.n4040 0.002
R52655 S.n4428 S.n4403 0.002
R52656 S.n2925 S.n2913 0.002
R52657 S.n3290 S.n3266 0.002
R52658 S.n1757 S.n1744 0.002
R52659 S.n2137 S.n2114 0.002
R52660 S.n726 S.n715 0.002
R52661 S.n406 S.n398 0.002
R52662 S.n16660 S.n16642 0.002
R52663 S.n15307 S.n15295 0.002
R52664 S.n15968 S.n15943 0.002
R52665 S.n14372 S.n14360 0.002
R52666 S.n15006 S.n14981 0.002
R52667 S.n13413 S.n13401 0.002
R52668 S.n14036 S.n14011 0.002
R52669 S.n12441 S.n12429 0.002
R52670 S.n13043 S.n13018 0.002
R52671 S.n11447 S.n11435 0.002
R52672 S.n12038 S.n12013 0.002
R52673 S.n10440 S.n10428 0.002
R52674 S.n11010 S.n10985 0.002
R52675 S.n9411 S.n9399 0.002
R52676 S.n9970 S.n9945 0.002
R52677 S.n8369 S.n8357 0.002
R52678 S.n8907 S.n8882 0.002
R52679 S.n7305 S.n7293 0.002
R52680 S.n7832 S.n7807 0.002
R52681 S.n6228 S.n6216 0.002
R52682 S.n6734 S.n6709 0.002
R52683 S.n5128 S.n5116 0.002
R52684 S.n5624 S.n5599 0.002
R52685 S.n4016 S.n4004 0.002
R52686 S.n4489 S.n4464 0.002
R52687 S.n2889 S.n2877 0.002
R52688 S.n3350 S.n3326 0.002
R52689 S.n1720 S.n1707 0.002
R52690 S.n2196 S.n2173 0.002
R52691 S.n691 S.n680 0.002
R52692 S.n374 S.n366 0.002
R52693 S.n14767 S.n14749 0.002
R52694 S.n13375 S.n13363 0.002
R52695 S.n14101 S.n14076 0.002
R52696 S.n12405 S.n12393 0.002
R52697 S.n13104 S.n13079 0.002
R52698 S.n11411 S.n11399 0.002
R52699 S.n12099 S.n12074 0.002
R52700 S.n10404 S.n10392 0.002
R52701 S.n11071 S.n11046 0.002
R52702 S.n9375 S.n9363 0.002
R52703 S.n10031 S.n10006 0.002
R52704 S.n8333 S.n8321 0.002
R52705 S.n8968 S.n8943 0.002
R52706 S.n7269 S.n7257 0.002
R52707 S.n7893 S.n7868 0.002
R52708 S.n6192 S.n6180 0.002
R52709 S.n6795 S.n6770 0.002
R52710 S.n5092 S.n5080 0.002
R52711 S.n5685 S.n5660 0.002
R52712 S.n3980 S.n3968 0.002
R52713 S.n4550 S.n4525 0.002
R52714 S.n2853 S.n2841 0.002
R52715 S.n3410 S.n3386 0.002
R52716 S.n1683 S.n1670 0.002
R52717 S.n2255 S.n2232 0.002
R52718 S.n656 S.n645 0.002
R52719 S.n342 S.n334 0.002
R52720 S.n12804 S.n12786 0.002
R52721 S.n11373 S.n11361 0.002
R52722 S.n12164 S.n12139 0.002
R52723 S.n10368 S.n10356 0.002
R52724 S.n11132 S.n11107 0.002
R52725 S.n9339 S.n9327 0.002
R52726 S.n10092 S.n10067 0.002
R52727 S.n8297 S.n8285 0.002
R52728 S.n9029 S.n9004 0.002
R52729 S.n7233 S.n7221 0.002
R52730 S.n7954 S.n7929 0.002
R52731 S.n6156 S.n6144 0.002
R52732 S.n6856 S.n6831 0.002
R52733 S.n5056 S.n5044 0.002
R52734 S.n5746 S.n5721 0.002
R52735 S.n3944 S.n3932 0.002
R52736 S.n4611 S.n4586 0.002
R52737 S.n2817 S.n2805 0.002
R52738 S.n3470 S.n3446 0.002
R52739 S.n1646 S.n1633 0.002
R52740 S.n2314 S.n2291 0.002
R52741 S.n621 S.n610 0.002
R52742 S.n310 S.n302 0.002
R52743 S.n10771 S.n10753 0.002
R52744 S.n9301 S.n9289 0.002
R52745 S.n10157 S.n10132 0.002
R52746 S.n8261 S.n8249 0.002
R52747 S.n9090 S.n9065 0.002
R52748 S.n7197 S.n7185 0.002
R52749 S.n8015 S.n7990 0.002
R52750 S.n6120 S.n6108 0.002
R52751 S.n6917 S.n6892 0.002
R52752 S.n5020 S.n5008 0.002
R52753 S.n5807 S.n5782 0.002
R52754 S.n3908 S.n3896 0.002
R52755 S.n4672 S.n4647 0.002
R52756 S.n2781 S.n2769 0.002
R52757 S.n3530 S.n3506 0.002
R52758 S.n1609 S.n1596 0.002
R52759 S.n2373 S.n2350 0.002
R52760 S.n586 S.n575 0.002
R52761 S.n278 S.n270 0.002
R52762 S.n8668 S.n8650 0.002
R52763 S.n7159 S.n7147 0.002
R52764 S.n8080 S.n8055 0.002
R52765 S.n6084 S.n6072 0.002
R52766 S.n6978 S.n6953 0.002
R52767 S.n4984 S.n4972 0.002
R52768 S.n5868 S.n5843 0.002
R52769 S.n3872 S.n3860 0.002
R52770 S.n4733 S.n4708 0.002
R52771 S.n2745 S.n2733 0.002
R52772 S.n3590 S.n3566 0.002
R52773 S.n1572 S.n1559 0.002
R52774 S.n2432 S.n2409 0.002
R52775 S.n551 S.n540 0.002
R52776 S.n249 S.n241 0.002
R52777 S.n6495 S.n6477 0.002
R52778 S.n4946 S.n4934 0.002
R52779 S.n5933 S.n5908 0.002
R52780 S.n3836 S.n3824 0.002
R52781 S.n4794 S.n4769 0.002
R52782 S.n2709 S.n2697 0.002
R52783 S.n3650 S.n3626 0.002
R52784 S.n1535 S.n1522 0.002
R52785 S.n2491 S.n2468 0.002
R52786 S.n516 S.n505 0.002
R52787 S.n214 S.n206 0.002
R52788 S.n4250 S.n4232 0.002
R52789 S.n2671 S.n2659 0.002
R52790 S.n3714 S.n3690 0.002
R52791 S.n1498 S.n1485 0.002
R52792 S.n2550 S.n2527 0.002
R52793 S.n481 S.n470 0.002
R52794 S.n182 S.n174 0.002
R52795 S.n1954 S.n1938 0.002
R52796 S.n447 S.n438 0.002
R52797 S.n150 S.n142 0.002
R52798 S.n23010 S.n23008 0.002
R52799 S.n1432 S.n1431 0.001
R52800 S.n2057 S.n2056 0.001
R52801 S.n1982 S.n1981 0.001
R52802 S.n2134 S.n2133 0.001
R52803 S.n2193 S.n2192 0.001
R52804 S.n2252 S.n2251 0.001
R52805 S.n2311 S.n2310 0.001
R52806 S.n2370 S.n2369 0.001
R52807 S.n2429 S.n2428 0.001
R52808 S.n2488 S.n2487 0.001
R52809 S.n1184 S.n1183 0.001
R52810 S.t158 S.n1184 0.001
R52811 S.n21189 S.n21188 0.001
R52812 S.n19414 S.n19413 0.001
R52813 S.n18527 S.n18526 0.001
R52814 S.n17627 S.n17626 0.001
R52815 S.n16704 S.n16703 0.001
R52816 S.n15769 S.n15768 0.001
R52817 S.n14811 S.n14810 0.001
R52818 S.n13841 S.n13840 0.001
R52819 S.n12848 S.n12847 0.001
R52820 S.n11843 S.n11842 0.001
R52821 S.n10815 S.n10814 0.001
R52822 S.n9775 S.n9774 0.001
R52823 S.n8712 S.n8711 0.001
R52824 S.n7637 S.n7636 0.001
R52825 S.n6539 S.n6538 0.001
R52826 S.n5428 S.n5427 0.001
R52827 S.n4294 S.n4293 0.001
R52828 S.n3157 S.n3156 0.001
R52829 S.n1996 S.n1995 0.001
R52830 S.n22978 S.n22976 0.001
R52831 S.n23008 S.t41 0.001
R52832 S.n3230 S.n3216 0.001
R52833 S.n968 S.n967 0.001
R52834 S.n427 S.n426 0.001
R52835 S.n1908 S.n1907 0.001
R52836 S.n1455 S.n1454 0.001
R52837 S.n2609 S.n2608 0.001
R52838 S.n2649 S.n2648 0.001
R52839 S.n3740 S.n3739 0.001
R52840 S.n3794 S.n3793 0.001
R52841 S.n4853 S.n4852 0.001
R52842 S.n4924 S.n4923 0.001
R52843 S.n5958 S.n5957 0.001
R52844 S.n6042 S.n6041 0.001
R52845 S.n7036 S.n7035 0.001
R52846 S.n7137 S.n7136 0.001
R52847 S.n8105 S.n8104 0.001
R52848 S.n8219 S.n8218 0.001
R52849 S.n9148 S.n9147 0.001
R52850 S.n9279 S.n9278 0.001
R52851 S.n10182 S.n10181 0.001
R52852 S.n10326 S.n10325 0.001
R52853 S.n11190 S.n11189 0.001
R52854 S.n11351 S.n11350 0.001
R52855 S.n12189 S.n12188 0.001
R52856 S.n12363 S.n12362 0.001
R52857 S.n13162 S.n13161 0.001
R52858 S.n13353 S.n13352 0.001
R52859 S.n14126 S.n14125 0.001
R52860 S.n14330 S.n14329 0.001
R52861 S.n15064 S.n15063 0.001
R52862 S.n15285 S.n15284 0.001
R52863 S.n15993 S.n15992 0.001
R52864 S.n16227 S.n16226 0.001
R52865 S.n16896 S.n16895 0.001
R52866 S.n17147 S.n17146 0.001
R52867 S.n17790 S.n17789 0.001
R52868 S.n18054 S.n18053 0.001
R52869 S.n18658 S.n18657 0.001
R52870 S.n18939 S.n18938 0.001
R52871 S.n19515 S.n19514 0.001
R52872 S.n19809 S.n19808 0.001
R52873 S.n21165 S.n21164 0.001
R52874 S.n20447 S.n20446 0.001
R52875 S.n21183 S.n21182 0.001
R52876 S.n21291 S.n21290 0.001
R52877 S.n22781 S.n22780 0.001
R52878 S.n22283 S.n22281 0.001
R52879 S.n22796 S.n22795 0.001
R52880 S.n19369 S.n19368 0.001
R52881 S.n17582 S.n17581 0.001
R52882 S.n15724 S.n15723 0.001
R52883 S.n13796 S.n13795 0.001
R52884 S.n11798 S.n11797 0.001
R52885 S.n9730 S.n9729 0.001
R52886 S.n7592 S.n7591 0.001
R52887 S.n5383 S.n5382 0.001
R52888 S.n3113 S.n3112 0.001
R52889 S.n21311 S.n21310 0.001
R52890 S.n20488 S.n20487 0.001
R52891 S.n17166 S.n17165 0.001
R52892 S.n16266 S.n16265 0.001
R52893 S.n18958 S.n18957 0.001
R52894 S.n18093 S.n18092 0.001
R52895 S.n15304 S.n15303 0.001
R52896 S.n14369 S.n14368 0.001
R52897 S.n13372 S.n13371 0.001
R52898 S.n12402 S.n12401 0.001
R52899 S.n11370 S.n11369 0.001
R52900 S.n10365 S.n10364 0.001
R52901 S.n9298 S.n9297 0.001
R52902 S.n8258 S.n8257 0.001
R52903 S.n7156 S.n7155 0.001
R52904 S.n6081 S.n6080 0.001
R52905 S.n4943 S.n4942 0.001
R52906 S.n3833 S.n3832 0.001
R52907 S.n2668 S.n2667 0.001
R52908 S.n1495 S.n1494 0.001
R52909 S.n939 S.n938 0.001
R52910 S.n22973 S.n22972 0.001
R52911 S.n22975 S.n22974 0.001
R52912 S.n1862 S.n1861 0.001
R52913 S.n3143 S.n3142 0.001
R52914 S.n3022 S.n3021 0.001
R52915 S.n4280 S.n4279 0.001
R52916 S.n4148 S.n4147 0.001
R52917 S.n5414 S.n5413 0.001
R52918 S.n5261 S.n5260 0.001
R52919 S.n6525 S.n6524 0.001
R52920 S.n6361 S.n6360 0.001
R52921 S.n7623 S.n7622 0.001
R52922 S.n7438 S.n7437 0.001
R52923 S.n8698 S.n8697 0.001
R52924 S.n8502 S.n8501 0.001
R52925 S.n9761 S.n9760 0.001
R52926 S.n9544 S.n9543 0.001
R52927 S.n10801 S.n10800 0.001
R52928 S.n10573 S.n10572 0.001
R52929 S.n11829 S.n11828 0.001
R52930 S.n11580 S.n11579 0.001
R52931 S.n12834 S.n12833 0.001
R52932 S.n12574 S.n12573 0.001
R52933 S.n13827 S.n13826 0.001
R52934 S.n13546 S.n13545 0.001
R52935 S.n14797 S.n14796 0.001
R52936 S.n14505 S.n14504 0.001
R52937 S.n15755 S.n15754 0.001
R52938 S.n15442 S.n15441 0.001
R52939 S.n16690 S.n16689 0.001
R52940 S.n16366 S.n16365 0.001
R52941 S.n17613 S.n17612 0.001
R52942 S.n17268 S.n17267 0.001
R52943 S.n18513 S.n18512 0.001
R52944 S.n18157 S.n18156 0.001
R52945 S.n19400 S.n19399 0.001
R52946 S.n19023 S.n19022 0.001
R52947 S.n20268 S.n20267 0.001
R52948 S.n19877 S.n19876 0.001
R52949 S.n1787 S.n1786 0.001
R52950 S.n3227 S.n3226 0.001
R52951 S.n2958 S.n2957 0.001
R52952 S.n4364 S.n4363 0.001
R52953 S.n4085 S.n4084 0.001
R52954 S.n5499 S.n5498 0.001
R52955 S.n5197 S.n5196 0.001
R52956 S.n6609 S.n6608 0.001
R52957 S.n6297 S.n6296 0.001
R52958 S.n7707 S.n7706 0.001
R52959 S.n7374 S.n7373 0.001
R52960 S.n8782 S.n8781 0.001
R52961 S.n8438 S.n8437 0.001
R52962 S.n9845 S.n9844 0.001
R52963 S.n9480 S.n9479 0.001
R52964 S.n10885 S.n10884 0.001
R52965 S.n10509 S.n10508 0.001
R52966 S.n11913 S.n11912 0.001
R52967 S.n11516 S.n11515 0.001
R52968 S.n12918 S.n12917 0.001
R52969 S.n12510 S.n12509 0.001
R52970 S.n13911 S.n13910 0.001
R52971 S.n13482 S.n13481 0.001
R52972 S.n14881 S.n14880 0.001
R52973 S.n14441 S.n14440 0.001
R52974 S.n15839 S.n15838 0.001
R52975 S.n15378 S.n15377 0.001
R52976 S.n16774 S.n16773 0.001
R52977 S.n16302 S.n16301 0.001
R52978 S.n17697 S.n17696 0.001
R52979 S.n17204 S.n17203 0.001
R52980 S.n1754 S.n1753 0.001
R52981 S.n3287 S.n3286 0.001
R52982 S.n2922 S.n2921 0.001
R52983 S.n4425 S.n4424 0.001
R52984 S.n4049 S.n4048 0.001
R52985 S.n5560 S.n5559 0.001
R52986 S.n5161 S.n5160 0.001
R52987 S.n6670 S.n6669 0.001
R52988 S.n6261 S.n6260 0.001
R52989 S.n7768 S.n7767 0.001
R52990 S.n7338 S.n7337 0.001
R52991 S.n8843 S.n8842 0.001
R52992 S.n8402 S.n8401 0.001
R52993 S.n9906 S.n9905 0.001
R52994 S.n9444 S.n9443 0.001
R52995 S.n10946 S.n10945 0.001
R52996 S.n10473 S.n10472 0.001
R52997 S.n11974 S.n11973 0.001
R52998 S.n11480 S.n11479 0.001
R52999 S.n12979 S.n12978 0.001
R53000 S.n12474 S.n12473 0.001
R53001 S.n13972 S.n13971 0.001
R53002 S.n13446 S.n13445 0.001
R53003 S.n14942 S.n14941 0.001
R53004 S.n14405 S.n14404 0.001
R53005 S.n15900 S.n15899 0.001
R53006 S.n15342 S.n15341 0.001
R53007 S.n1717 S.n1716 0.001
R53008 S.n3347 S.n3346 0.001
R53009 S.n2886 S.n2885 0.001
R53010 S.n4486 S.n4485 0.001
R53011 S.n4013 S.n4012 0.001
R53012 S.n5621 S.n5620 0.001
R53013 S.n5125 S.n5124 0.001
R53014 S.n6731 S.n6730 0.001
R53015 S.n6225 S.n6224 0.001
R53016 S.n7829 S.n7828 0.001
R53017 S.n7302 S.n7301 0.001
R53018 S.n8904 S.n8903 0.001
R53019 S.n8366 S.n8365 0.001
R53020 S.n9967 S.n9966 0.001
R53021 S.n9408 S.n9407 0.001
R53022 S.n11007 S.n11006 0.001
R53023 S.n10437 S.n10436 0.001
R53024 S.n12035 S.n12034 0.001
R53025 S.n11444 S.n11443 0.001
R53026 S.n13040 S.n13039 0.001
R53027 S.n12438 S.n12437 0.001
R53028 S.n14033 S.n14032 0.001
R53029 S.n13410 S.n13409 0.001
R53030 S.n1680 S.n1679 0.001
R53031 S.n3407 S.n3406 0.001
R53032 S.n2850 S.n2849 0.001
R53033 S.n4547 S.n4546 0.001
R53034 S.n3977 S.n3976 0.001
R53035 S.n5682 S.n5681 0.001
R53036 S.n5089 S.n5088 0.001
R53037 S.n6792 S.n6791 0.001
R53038 S.n6189 S.n6188 0.001
R53039 S.n7890 S.n7889 0.001
R53040 S.n7266 S.n7265 0.001
R53041 S.n8965 S.n8964 0.001
R53042 S.n8330 S.n8329 0.001
R53043 S.n10028 S.n10027 0.001
R53044 S.n9372 S.n9371 0.001
R53045 S.n11068 S.n11067 0.001
R53046 S.n10401 S.n10400 0.001
R53047 S.n12096 S.n12095 0.001
R53048 S.n11408 S.n11407 0.001
R53049 S.n1643 S.n1642 0.001
R53050 S.n3467 S.n3466 0.001
R53051 S.n2814 S.n2813 0.001
R53052 S.n4608 S.n4607 0.001
R53053 S.n3941 S.n3940 0.001
R53054 S.n5743 S.n5742 0.001
R53055 S.n5053 S.n5052 0.001
R53056 S.n6853 S.n6852 0.001
R53057 S.n6153 S.n6152 0.001
R53058 S.n7951 S.n7950 0.001
R53059 S.n7230 S.n7229 0.001
R53060 S.n9026 S.n9025 0.001
R53061 S.n8294 S.n8293 0.001
R53062 S.n10089 S.n10088 0.001
R53063 S.n9336 S.n9335 0.001
R53064 S.n1606 S.n1605 0.001
R53065 S.n3527 S.n3526 0.001
R53066 S.n2778 S.n2777 0.001
R53067 S.n4669 S.n4668 0.001
R53068 S.n3905 S.n3904 0.001
R53069 S.n5804 S.n5803 0.001
R53070 S.n5017 S.n5016 0.001
R53071 S.n6914 S.n6913 0.001
R53072 S.n6117 S.n6116 0.001
R53073 S.n8012 S.n8011 0.001
R53074 S.n7194 S.n7193 0.001
R53075 S.n1569 S.n1568 0.001
R53076 S.n3587 S.n3586 0.001
R53077 S.n2742 S.n2741 0.001
R53078 S.n4730 S.n4729 0.001
R53079 S.n3869 S.n3868 0.001
R53080 S.n5865 S.n5864 0.001
R53081 S.n4981 S.n4980 0.001
R53082 S.n1532 S.n1531 0.001
R53083 S.n3647 S.n3646 0.001
R53084 S.n2706 S.n2705 0.001
R53085 S.n22750 S.n22749 0.001
R53086 S.n16788 S.n16787 0.001
R53087 S.n15853 S.n15852 0.001
R53088 S.n14895 S.n14894 0.001
R53089 S.n13925 S.n13924 0.001
R53090 S.n12932 S.n12931 0.001
R53091 S.n11927 S.n11926 0.001
R53092 S.n10899 S.n10898 0.001
R53093 S.n9859 S.n9858 0.001
R53094 S.n8796 S.n8795 0.001
R53095 S.n7721 S.n7720 0.001
R53096 S.n6623 S.n6622 0.001
R53097 S.n5513 S.n5512 0.001
R53098 S.n4378 S.n4377 0.001
R53099 S.n3241 S.n3240 0.001
R53100 S.n2091 S.n2090 0.001
R53101 S.n14956 S.n14955 0.001
R53102 S.n13986 S.n13985 0.001
R53103 S.n12993 S.n12992 0.001
R53104 S.n11988 S.n11987 0.001
R53105 S.n10960 S.n10959 0.001
R53106 S.n9920 S.n9919 0.001
R53107 S.n8857 S.n8856 0.001
R53108 S.n7782 S.n7781 0.001
R53109 S.n6684 S.n6683 0.001
R53110 S.n5574 S.n5573 0.001
R53111 S.n4439 S.n4438 0.001
R53112 S.n3301 S.n3300 0.001
R53113 S.n2149 S.n2148 0.001
R53114 S.n13054 S.n13053 0.001
R53115 S.n12049 S.n12048 0.001
R53116 S.n11021 S.n11020 0.001
R53117 S.n9981 S.n9980 0.001
R53118 S.n8918 S.n8917 0.001
R53119 S.n7843 S.n7842 0.001
R53120 S.n6745 S.n6744 0.001
R53121 S.n5635 S.n5634 0.001
R53122 S.n4500 S.n4499 0.001
R53123 S.n3361 S.n3360 0.001
R53124 S.n2208 S.n2207 0.001
R53125 S.n11082 S.n11081 0.001
R53126 S.n10042 S.n10041 0.001
R53127 S.n8979 S.n8978 0.001
R53128 S.n7904 S.n7903 0.001
R53129 S.n6806 S.n6805 0.001
R53130 S.n5696 S.n5695 0.001
R53131 S.n4561 S.n4560 0.001
R53132 S.n3421 S.n3420 0.001
R53133 S.n2267 S.n2266 0.001
R53134 S.n9040 S.n9039 0.001
R53135 S.n7965 S.n7964 0.001
R53136 S.n6867 S.n6866 0.001
R53137 S.n5757 S.n5756 0.001
R53138 S.n4622 S.n4621 0.001
R53139 S.n3481 S.n3480 0.001
R53140 S.n2326 S.n2325 0.001
R53141 S.n6928 S.n6927 0.001
R53142 S.n5818 S.n5817 0.001
R53143 S.n4683 S.n4682 0.001
R53144 S.n3541 S.n3540 0.001
R53145 S.n2385 S.n2384 0.001
R53146 S.n4744 S.n4743 0.001
R53147 S.n3601 S.n3600 0.001
R53148 S.n2444 S.n2443 0.001
R53149 S.n2503 S.n2502 0.001
R53150 S.n3057 S.n3049 0.001
R53151 S.n1900 S.n1899 0.001
R53152 S.n806 S.n795 0.001
R53153 S.n1433 S.n1432 0.001
R53154 S.t158 S.n26 0.001
R53155 S.t158 S.n1309 0.001
R53156 S.t158 S.n1339 0.001
R53157 S.t158 S.n73 0.001
R53158 S.t158 S.n105 0.001
R53159 S.t158 S.n992 0.001
R53160 S.t158 S.n1024 0.001
R53161 S.t158 S.n1056 0.001
R53162 S.t158 S.n1088 0.001
R53163 S.t158 S.n1120 0.001
R53164 S.t158 S.n1158 0.001
R53165 S.t158 S.n1369 0.001
R53166 S.t158 S.n1295 0.001
R53167 S.t158 S.n1283 0.001
R53168 S.t158 S.n1271 0.001
R53169 S.t158 S.n1258 0.001
R53170 S.t158 S.n1245 0.001
R53171 S.t158 S.n1232 0.001
R53172 S.t158 S.n1219 0.001
R53173 S.t158 S.n1206 0.001
R53174 S.t158 S.n1193 0.001
R53175 S.t158 S.n1170 0.001
R53176 S.n19490 S.n19475 0.001
R53177 S.n18600 S.n18585 0.001
R53178 S.n17700 S.n17685 0.001
R53179 S.n16777 S.n16762 0.001
R53180 S.n15842 S.n15827 0.001
R53181 S.n14884 S.n14869 0.001
R53182 S.n13914 S.n13899 0.001
R53183 S.n12921 S.n12906 0.001
R53184 S.n11916 S.n11901 0.001
R53185 S.n10888 S.n10873 0.001
R53186 S.n9848 S.n9833 0.001
R53187 S.n8785 S.n8770 0.001
R53188 S.n7710 S.n7695 0.001
R53189 S.n6612 S.n6597 0.001
R53190 S.n5502 S.n5487 0.001
R53191 S.n4367 S.n4352 0.001
R53192 S.n22289 S.n22288 0.001
R53193 S.n18060 S.n18059 0.001
R53194 S.n19815 S.n19814 0.001
R53195 S.n20452 S.n20451 0.001
R53196 S.n21297 S.n21296 0.001
R53197 S.n18944 S.n18943 0.001
R53198 S.n16233 S.n16232 0.001
R53199 S.n17152 S.n17151 0.001
R53200 S.n14336 S.n14335 0.001
R53201 S.n15290 S.n15289 0.001
R53202 S.n12369 S.n12368 0.001
R53203 S.n13358 S.n13357 0.001
R53204 S.n10332 S.n10331 0.001
R53205 S.n11356 S.n11355 0.001
R53206 S.n8225 S.n8224 0.001
R53207 S.n9284 S.n9283 0.001
R53208 S.n6048 S.n6047 0.001
R53209 S.n7142 S.n7141 0.001
R53210 S.n3800 S.n3799 0.001
R53211 S.n4929 S.n4928 0.001
R53212 S.n1461 S.n1460 0.001
R53213 S.n2654 S.n2653 0.001
R53214 S.n433 S.n432 0.001
R53215 S.n22791 S.n22774 0.001
R53216 S.n43 S.n41 0.001
R53217 S.n901 S.n900 0.001
R53218 S.n20238 S.n20219 0.001
R53219 S.n395 S.n394 0.001
R53220 S.n363 S.n362 0.001
R53221 S.n331 S.n330 0.001
R53222 S.n299 S.n298 0.001
R53223 S.n266 S.n265 0.001
R53224 S.n237 S.n236 0.001
R53225 S.n203 S.n202 0.001
R53226 S.n171 S.n170 0.001
R53227 S.n138 S.n137 0.001
R53228 S.n22324 S.n22323 0.001
R53229 S.n22336 S.n22333 0.001
R53230 S.t9 S.n22336 0.001
R53231 S.n22774 S.t88 0.001
R53232 S.t9 S.n22289 0.001
R53233 S.t79 S.n18060 0.001
R53234 S.t150 S.n18944 0.001
R53235 S.t209 S.n19815 0.001
R53236 S.t64 S.n20452 0.001
R53237 S.t100 S.n21297 0.001
R53238 S.t167 S.n16233 0.001
R53239 S.t218 S.n17152 0.001
R53240 S.t0 S.n14336 0.001
R53241 S.t60 S.n15290 0.001
R53242 S.t357 S.n12369 0.001
R53243 S.t73 S.n13358 0.001
R53244 S.t31 S.n10332 0.001
R53245 S.t54 S.n11356 0.001
R53246 S.t19 S.n8225 0.001
R53247 S.t366 S.n9284 0.001
R53248 S.t83 S.n6048 0.001
R53249 S.t47 S.n7142 0.001
R53250 S.t176 S.n3800 0.001
R53251 S.t214 S.n4929 0.001
R53252 S.t75 S.n1461 0.001
R53253 S.t14 S.n2654 0.001
R53254 S.t137 S.n433 0.001
R53255 S.n43 S.n40 0.001
R53256 S.n4842 S.n4841 0.001
R53257 S.n2598 S.n2597 0.001
R53258 S.n891 S.n890 0.001
R53259 S.n824 S.n823 0.001
R53260 S.n43 S.n37 0.001
R53261 S.n43 S.n36 0.001
R53262 S.n43 S.n35 0.001
R53263 S.n43 S.n34 0.001
R53264 S.n43 S.n33 0.001
R53265 S.n43 S.n32 0.001
R53266 S.n43 S.n31 0.001
R53267 S.n43 S.n30 0.001
R53268 S.n43 S.n29 0.001
R53269 S.n43 S.n39 0.001
R53270 S.n22978 S.n22975 0.001
R53271 S.n22978 S.n22973 0.001
R53272 S.n726 S.n718 0.001
R53273 S.n691 S.n683 0.001
R53274 S.n656 S.n648 0.001
R53275 S.n621 S.n613 0.001
R53276 S.n586 S.n578 0.001
R53277 S.n551 S.n543 0.001
R53278 S.n516 S.n508 0.001
R53279 S.n481 S.n473 0.001
R53280 S.n447 S.n439 0.001
R53281 S.n969 S.n968 0.001
R53282 S.n426 S.n425 0.001
R53283 S.n1909 S.n1908 0.001
R53284 S.n1454 S.n1453 0.001
R53285 S.n2610 S.n2609 0.001
R53286 S.n2648 S.n2647 0.001
R53287 S.n3741 S.n3740 0.001
R53288 S.n3793 S.n3792 0.001
R53289 S.n4854 S.n4853 0.001
R53290 S.n4923 S.n4922 0.001
R53291 S.n5959 S.n5958 0.001
R53292 S.n6041 S.n6040 0.001
R53293 S.n7037 S.n7036 0.001
R53294 S.n7136 S.n7135 0.001
R53295 S.n8106 S.n8105 0.001
R53296 S.n8218 S.n8217 0.001
R53297 S.n9149 S.n9148 0.001
R53298 S.n9278 S.n9277 0.001
R53299 S.n10183 S.n10182 0.001
R53300 S.n10325 S.n10324 0.001
R53301 S.n11191 S.n11190 0.001
R53302 S.n11350 S.n11349 0.001
R53303 S.n12190 S.n12189 0.001
R53304 S.n12362 S.n12361 0.001
R53305 S.n13163 S.n13162 0.001
R53306 S.n13352 S.n13351 0.001
R53307 S.n14127 S.n14126 0.001
R53308 S.n14329 S.n14328 0.001
R53309 S.n15065 S.n15064 0.001
R53310 S.n15284 S.n15283 0.001
R53311 S.n15994 S.n15993 0.001
R53312 S.n16226 S.n16225 0.001
R53313 S.n16897 S.n16896 0.001
R53314 S.n17146 S.n17145 0.001
R53315 S.n17791 S.n17790 0.001
R53316 S.n18053 S.n18052 0.001
R53317 S.n18659 S.n18658 0.001
R53318 S.n18938 S.n18937 0.001
R53319 S.n19516 S.n19515 0.001
R53320 S.n19808 S.n19807 0.001
R53321 S.n21166 S.n21165 0.001
R53322 S.n20446 S.n20445 0.001
R53323 S.n21184 S.n21183 0.001
R53324 S.n21290 S.n21289 0.001
R53325 S.n22782 S.n22781 0.001
R53326 S.n22281 S.n22280 0.001
R53327 S.n22797 S.n22796 0.001
R53328 S.n20178 S.n20177 0.001
R53329 S.n21132 S.n21131 0.001
R53330 S.n22638 S.n22637 0.001
R53331 S.n22009 S.n22008 0.001
R53332 S.n21615 S.n21614 0.001
R53333 S.n21941 S.n21940 0.001
R53334 S.n20792 S.n20791 0.001
R53335 S.n22651 S.n22650 0.001
R53336 S.n21990 S.n21989 0.001
R53337 S.n21633 S.n21632 0.001
R53338 S.n21956 S.n21955 0.001
R53339 S.n20810 S.n20809 0.001
R53340 S.n19308 S.n19307 0.001
R53341 S.n19532 S.n19531 0.001
R53342 S.n22622 S.n22621 0.001
R53343 S.n22024 S.n22023 0.001
R53344 S.n21599 S.n21598 0.001
R53345 S.n21926 S.n21925 0.001
R53346 S.n20776 S.n20775 0.001
R53347 S.n21116 S.n21115 0.001
R53348 S.n20165 S.n20164 0.001
R53349 S.n18426 S.n18425 0.001
R53350 S.n18675 S.n18674 0.001
R53351 S.n22606 S.n22605 0.001
R53352 S.n22039 S.n22038 0.001
R53353 S.n21583 S.n21582 0.001
R53354 S.n21911 S.n21910 0.001
R53355 S.n20760 S.n20759 0.001
R53356 S.n21101 S.n21100 0.001
R53357 S.n20149 S.n20148 0.001
R53358 S.n19547 S.n19546 0.001
R53359 S.n19295 S.n19294 0.001
R53360 S.n17521 S.n17520 0.001
R53361 S.n17807 S.n17806 0.001
R53362 S.n22590 S.n22589 0.001
R53363 S.n22054 S.n22053 0.001
R53364 S.n21567 S.n21566 0.001
R53365 S.n21896 S.n21895 0.001
R53366 S.n20744 S.n20743 0.001
R53367 S.n21086 S.n21085 0.001
R53368 S.n20133 S.n20132 0.001
R53369 S.n19562 S.n19561 0.001
R53370 S.n19279 S.n19278 0.001
R53371 S.n18690 S.n18689 0.001
R53372 S.n18413 S.n18412 0.001
R53373 S.n16603 S.n16602 0.001
R53374 S.n16913 S.n16912 0.001
R53375 S.n22574 S.n22573 0.001
R53376 S.n22069 S.n22068 0.001
R53377 S.n21551 S.n21550 0.001
R53378 S.n21881 S.n21880 0.001
R53379 S.n20728 S.n20727 0.001
R53380 S.n21071 S.n21070 0.001
R53381 S.n20117 S.n20116 0.001
R53382 S.n19577 S.n19576 0.001
R53383 S.n19263 S.n19262 0.001
R53384 S.n18705 S.n18704 0.001
R53385 S.n18397 S.n18396 0.001
R53386 S.n17822 S.n17821 0.001
R53387 S.n17508 S.n17507 0.001
R53388 S.n15663 S.n15662 0.001
R53389 S.n16010 S.n16009 0.001
R53390 S.n22558 S.n22557 0.001
R53391 S.n22084 S.n22083 0.001
R53392 S.n21535 S.n21534 0.001
R53393 S.n21866 S.n21865 0.001
R53394 S.n20712 S.n20711 0.001
R53395 S.n21056 S.n21055 0.001
R53396 S.n20101 S.n20100 0.001
R53397 S.n19592 S.n19591 0.001
R53398 S.n19247 S.n19246 0.001
R53399 S.n18720 S.n18719 0.001
R53400 S.n18381 S.n18380 0.001
R53401 S.n17837 S.n17836 0.001
R53402 S.n17492 S.n17491 0.001
R53403 S.n16928 S.n16927 0.001
R53404 S.n16590 S.n16589 0.001
R53405 S.n14710 S.n14709 0.001
R53406 S.n15081 S.n15080 0.001
R53407 S.n22542 S.n22541 0.001
R53408 S.n22099 S.n22098 0.001
R53409 S.n21519 S.n21518 0.001
R53410 S.n21851 S.n21850 0.001
R53411 S.n20696 S.n20695 0.001
R53412 S.n21041 S.n21040 0.001
R53413 S.n20085 S.n20084 0.001
R53414 S.n19607 S.n19606 0.001
R53415 S.n19231 S.n19230 0.001
R53416 S.n18735 S.n18734 0.001
R53417 S.n18365 S.n18364 0.001
R53418 S.n17852 S.n17851 0.001
R53419 S.n17476 S.n17475 0.001
R53420 S.n16943 S.n16942 0.001
R53421 S.n16574 S.n16573 0.001
R53422 S.n16025 S.n16024 0.001
R53423 S.n15650 S.n15649 0.001
R53424 S.n13735 S.n13734 0.001
R53425 S.n14143 S.n14142 0.001
R53426 S.n22526 S.n22525 0.001
R53427 S.n22114 S.n22113 0.001
R53428 S.n21503 S.n21502 0.001
R53429 S.n21836 S.n21835 0.001
R53430 S.n20680 S.n20679 0.001
R53431 S.n21026 S.n21025 0.001
R53432 S.n20069 S.n20068 0.001
R53433 S.n19622 S.n19621 0.001
R53434 S.n19215 S.n19214 0.001
R53435 S.n18750 S.n18749 0.001
R53436 S.n18349 S.n18348 0.001
R53437 S.n17867 S.n17866 0.001
R53438 S.n17460 S.n17459 0.001
R53439 S.n16958 S.n16957 0.001
R53440 S.n16558 S.n16557 0.001
R53441 S.n16040 S.n16039 0.001
R53442 S.n15634 S.n15633 0.001
R53443 S.n15096 S.n15095 0.001
R53444 S.n14697 S.n14696 0.001
R53445 S.n12747 S.n12746 0.001
R53446 S.n13179 S.n13178 0.001
R53447 S.n22510 S.n22509 0.001
R53448 S.n22129 S.n22128 0.001
R53449 S.n21487 S.n21486 0.001
R53450 S.n21821 S.n21820 0.001
R53451 S.n20664 S.n20663 0.001
R53452 S.n21011 S.n21010 0.001
R53453 S.n20053 S.n20052 0.001
R53454 S.n19637 S.n19636 0.001
R53455 S.n19199 S.n19198 0.001
R53456 S.n18765 S.n18764 0.001
R53457 S.n18333 S.n18332 0.001
R53458 S.n17882 S.n17881 0.001
R53459 S.n17444 S.n17443 0.001
R53460 S.n16973 S.n16972 0.001
R53461 S.n16542 S.n16541 0.001
R53462 S.n16055 S.n16054 0.001
R53463 S.n15618 S.n15617 0.001
R53464 S.n15111 S.n15110 0.001
R53465 S.n14681 S.n14680 0.001
R53466 S.n14158 S.n14157 0.001
R53467 S.n13722 S.n13721 0.001
R53468 S.n11737 S.n11736 0.001
R53469 S.n12206 S.n12205 0.001
R53470 S.n22494 S.n22493 0.001
R53471 S.n22144 S.n22143 0.001
R53472 S.n21471 S.n21470 0.001
R53473 S.n21806 S.n21805 0.001
R53474 S.n20648 S.n20647 0.001
R53475 S.n20996 S.n20995 0.001
R53476 S.n20037 S.n20036 0.001
R53477 S.n19652 S.n19651 0.001
R53478 S.n19183 S.n19182 0.001
R53479 S.n18780 S.n18779 0.001
R53480 S.n18317 S.n18316 0.001
R53481 S.n17897 S.n17896 0.001
R53482 S.n17428 S.n17427 0.001
R53483 S.n16988 S.n16987 0.001
R53484 S.n16526 S.n16525 0.001
R53485 S.n16070 S.n16069 0.001
R53486 S.n15602 S.n15601 0.001
R53487 S.n15126 S.n15125 0.001
R53488 S.n14665 S.n14664 0.001
R53489 S.n14173 S.n14172 0.001
R53490 S.n13706 S.n13705 0.001
R53491 S.n13194 S.n13193 0.001
R53492 S.n12734 S.n12733 0.001
R53493 S.n10714 S.n10713 0.001
R53494 S.n11207 S.n11206 0.001
R53495 S.n22478 S.n22477 0.001
R53496 S.n22159 S.n22158 0.001
R53497 S.n21455 S.n21454 0.001
R53498 S.n21791 S.n21790 0.001
R53499 S.n20632 S.n20631 0.001
R53500 S.n20981 S.n20980 0.001
R53501 S.n20021 S.n20020 0.001
R53502 S.n19667 S.n19666 0.001
R53503 S.n19167 S.n19166 0.001
R53504 S.n18795 S.n18794 0.001
R53505 S.n18301 S.n18300 0.001
R53506 S.n17912 S.n17911 0.001
R53507 S.n17412 S.n17411 0.001
R53508 S.n17003 S.n17002 0.001
R53509 S.n16510 S.n16509 0.001
R53510 S.n16085 S.n16084 0.001
R53511 S.n15586 S.n15585 0.001
R53512 S.n15141 S.n15140 0.001
R53513 S.n14649 S.n14648 0.001
R53514 S.n14188 S.n14187 0.001
R53515 S.n13690 S.n13689 0.001
R53516 S.n13209 S.n13208 0.001
R53517 S.n12718 S.n12717 0.001
R53518 S.n12221 S.n12220 0.001
R53519 S.n11724 S.n11723 0.001
R53520 S.n9669 S.n9668 0.001
R53521 S.n10199 S.n10198 0.001
R53522 S.n22462 S.n22461 0.001
R53523 S.n22174 S.n22173 0.001
R53524 S.n21439 S.n21438 0.001
R53525 S.n21776 S.n21775 0.001
R53526 S.n20616 S.n20615 0.001
R53527 S.n20966 S.n20965 0.001
R53528 S.n20005 S.n20004 0.001
R53529 S.n19682 S.n19681 0.001
R53530 S.n19151 S.n19150 0.001
R53531 S.n18810 S.n18809 0.001
R53532 S.n18285 S.n18284 0.001
R53533 S.n17927 S.n17926 0.001
R53534 S.n17396 S.n17395 0.001
R53535 S.n17018 S.n17017 0.001
R53536 S.n16494 S.n16493 0.001
R53537 S.n16100 S.n16099 0.001
R53538 S.n15570 S.n15569 0.001
R53539 S.n15156 S.n15155 0.001
R53540 S.n14633 S.n14632 0.001
R53541 S.n14203 S.n14202 0.001
R53542 S.n13674 S.n13673 0.001
R53543 S.n13224 S.n13223 0.001
R53544 S.n12702 S.n12701 0.001
R53545 S.n12236 S.n12235 0.001
R53546 S.n11708 S.n11707 0.001
R53547 S.n11222 S.n11221 0.001
R53548 S.n10701 S.n10700 0.001
R53549 S.n8611 S.n8610 0.001
R53550 S.n9165 S.n9164 0.001
R53551 S.n22446 S.n22445 0.001
R53552 S.n22189 S.n22188 0.001
R53553 S.n21423 S.n21422 0.001
R53554 S.n21761 S.n21760 0.001
R53555 S.n20600 S.n20599 0.001
R53556 S.n20951 S.n20950 0.001
R53557 S.n19989 S.n19988 0.001
R53558 S.n19697 S.n19696 0.001
R53559 S.n19135 S.n19134 0.001
R53560 S.n18825 S.n18824 0.001
R53561 S.n18269 S.n18268 0.001
R53562 S.n17942 S.n17941 0.001
R53563 S.n17380 S.n17379 0.001
R53564 S.n17033 S.n17032 0.001
R53565 S.n16478 S.n16477 0.001
R53566 S.n16115 S.n16114 0.001
R53567 S.n15554 S.n15553 0.001
R53568 S.n15171 S.n15170 0.001
R53569 S.n14617 S.n14616 0.001
R53570 S.n14218 S.n14217 0.001
R53571 S.n13658 S.n13657 0.001
R53572 S.n13239 S.n13238 0.001
R53573 S.n12686 S.n12685 0.001
R53574 S.n12251 S.n12250 0.001
R53575 S.n11692 S.n11691 0.001
R53576 S.n11237 S.n11236 0.001
R53577 S.n10685 S.n10684 0.001
R53578 S.n10214 S.n10213 0.001
R53579 S.n9656 S.n9655 0.001
R53580 S.n7531 S.n7530 0.001
R53581 S.n8122 S.n8121 0.001
R53582 S.n22430 S.n22429 0.001
R53583 S.n22204 S.n22203 0.001
R53584 S.n21407 S.n21406 0.001
R53585 S.n21746 S.n21745 0.001
R53586 S.n20584 S.n20583 0.001
R53587 S.n20936 S.n20935 0.001
R53588 S.n19973 S.n19972 0.001
R53589 S.n19712 S.n19711 0.001
R53590 S.n19119 S.n19118 0.001
R53591 S.n18840 S.n18839 0.001
R53592 S.n18253 S.n18252 0.001
R53593 S.n17957 S.n17956 0.001
R53594 S.n17364 S.n17363 0.001
R53595 S.n17048 S.n17047 0.001
R53596 S.n16462 S.n16461 0.001
R53597 S.n16130 S.n16129 0.001
R53598 S.n15538 S.n15537 0.001
R53599 S.n15186 S.n15185 0.001
R53600 S.n14601 S.n14600 0.001
R53601 S.n14233 S.n14232 0.001
R53602 S.n13642 S.n13641 0.001
R53603 S.n13254 S.n13253 0.001
R53604 S.n12670 S.n12669 0.001
R53605 S.n12266 S.n12265 0.001
R53606 S.n11676 S.n11675 0.001
R53607 S.n11252 S.n11251 0.001
R53608 S.n10669 S.n10668 0.001
R53609 S.n10229 S.n10228 0.001
R53610 S.n9640 S.n9639 0.001
R53611 S.n9180 S.n9179 0.001
R53612 S.n8598 S.n8597 0.001
R53613 S.n6438 S.n6437 0.001
R53614 S.n7053 S.n7052 0.001
R53615 S.n22414 S.n22413 0.001
R53616 S.n22219 S.n22218 0.001
R53617 S.n21391 S.n21390 0.001
R53618 S.n21731 S.n21730 0.001
R53619 S.n20568 S.n20567 0.001
R53620 S.n20921 S.n20920 0.001
R53621 S.n19957 S.n19956 0.001
R53622 S.n19727 S.n19726 0.001
R53623 S.n19103 S.n19102 0.001
R53624 S.n18855 S.n18854 0.001
R53625 S.n18237 S.n18236 0.001
R53626 S.n17972 S.n17971 0.001
R53627 S.n17348 S.n17347 0.001
R53628 S.n17063 S.n17062 0.001
R53629 S.n16446 S.n16445 0.001
R53630 S.n16145 S.n16144 0.001
R53631 S.n15522 S.n15521 0.001
R53632 S.n15201 S.n15200 0.001
R53633 S.n14585 S.n14584 0.001
R53634 S.n14248 S.n14247 0.001
R53635 S.n13626 S.n13625 0.001
R53636 S.n13269 S.n13268 0.001
R53637 S.n12654 S.n12653 0.001
R53638 S.n12281 S.n12280 0.001
R53639 S.n11660 S.n11659 0.001
R53640 S.n11267 S.n11266 0.001
R53641 S.n10653 S.n10652 0.001
R53642 S.n10244 S.n10243 0.001
R53643 S.n9624 S.n9623 0.001
R53644 S.n9195 S.n9194 0.001
R53645 S.n8582 S.n8581 0.001
R53646 S.n8137 S.n8136 0.001
R53647 S.n7518 S.n7517 0.001
R53648 S.n5322 S.n5321 0.001
R53649 S.n5975 S.n5974 0.001
R53650 S.n22398 S.n22397 0.001
R53651 S.n22234 S.n22233 0.001
R53652 S.n21375 S.n21374 0.001
R53653 S.n21716 S.n21715 0.001
R53654 S.n20552 S.n20551 0.001
R53655 S.n20906 S.n20905 0.001
R53656 S.n19941 S.n19940 0.001
R53657 S.n19742 S.n19741 0.001
R53658 S.n19087 S.n19086 0.001
R53659 S.n18870 S.n18869 0.001
R53660 S.n18221 S.n18220 0.001
R53661 S.n17987 S.n17986 0.001
R53662 S.n17332 S.n17331 0.001
R53663 S.n17078 S.n17077 0.001
R53664 S.n16430 S.n16429 0.001
R53665 S.n16160 S.n16159 0.001
R53666 S.n15506 S.n15505 0.001
R53667 S.n15216 S.n15215 0.001
R53668 S.n14569 S.n14568 0.001
R53669 S.n14263 S.n14262 0.001
R53670 S.n13610 S.n13609 0.001
R53671 S.n13284 S.n13283 0.001
R53672 S.n12638 S.n12637 0.001
R53673 S.n12296 S.n12295 0.001
R53674 S.n11644 S.n11643 0.001
R53675 S.n11282 S.n11281 0.001
R53676 S.n10637 S.n10636 0.001
R53677 S.n10259 S.n10258 0.001
R53678 S.n9608 S.n9607 0.001
R53679 S.n9210 S.n9209 0.001
R53680 S.n8566 S.n8565 0.001
R53681 S.n8152 S.n8151 0.001
R53682 S.n7502 S.n7501 0.001
R53683 S.n7068 S.n7067 0.001
R53684 S.n6425 S.n6424 0.001
R53685 S.n4193 S.n4192 0.001
R53686 S.n4870 S.n4869 0.001
R53687 S.n22382 S.n22381 0.001
R53688 S.n22249 S.n22248 0.001
R53689 S.n21359 S.n21358 0.001
R53690 S.n21701 S.n21700 0.001
R53691 S.n20536 S.n20535 0.001
R53692 S.n20891 S.n20890 0.001
R53693 S.n19925 S.n19924 0.001
R53694 S.n19757 S.n19756 0.001
R53695 S.n19071 S.n19070 0.001
R53696 S.n18885 S.n18884 0.001
R53697 S.n18205 S.n18204 0.001
R53698 S.n18002 S.n18001 0.001
R53699 S.n17316 S.n17315 0.001
R53700 S.n17093 S.n17092 0.001
R53701 S.n16414 S.n16413 0.001
R53702 S.n16175 S.n16174 0.001
R53703 S.n15490 S.n15489 0.001
R53704 S.n15231 S.n15230 0.001
R53705 S.n14553 S.n14552 0.001
R53706 S.n14278 S.n14277 0.001
R53707 S.n13594 S.n13593 0.001
R53708 S.n13299 S.n13298 0.001
R53709 S.n12622 S.n12621 0.001
R53710 S.n12311 S.n12310 0.001
R53711 S.n11628 S.n11627 0.001
R53712 S.n11297 S.n11296 0.001
R53713 S.n10621 S.n10620 0.001
R53714 S.n10274 S.n10273 0.001
R53715 S.n9592 S.n9591 0.001
R53716 S.n9228 S.n9227 0.001
R53717 S.n8550 S.n8549 0.001
R53718 S.n8167 S.n8166 0.001
R53719 S.n7486 S.n7485 0.001
R53720 S.n7083 S.n7082 0.001
R53721 S.n6409 S.n6408 0.001
R53722 S.n5990 S.n5989 0.001
R53723 S.n5309 S.n5308 0.001
R53724 S.n3052 S.n3051 0.001
R53725 S.n3757 S.n3756 0.001
R53726 S.n22671 S.n22670 0.001
R53727 S.n22264 S.n22263 0.001
R53728 S.n21684 S.n21683 0.001
R53729 S.n21670 S.n21669 0.001
R53730 S.n20521 S.n20520 0.001
R53731 S.n20875 S.n20874 0.001
R53732 S.n19910 S.n19909 0.001
R53733 S.n19772 S.n19771 0.001
R53734 S.n19056 S.n19055 0.001
R53735 S.n18900 S.n18899 0.001
R53736 S.n18190 S.n18189 0.001
R53737 S.n18017 S.n18016 0.001
R53738 S.n17301 S.n17300 0.001
R53739 S.n17108 S.n17107 0.001
R53740 S.n16399 S.n16398 0.001
R53741 S.n16190 S.n16189 0.001
R53742 S.n15475 S.n15474 0.001
R53743 S.n15246 S.n15245 0.001
R53744 S.n14538 S.n14537 0.001
R53745 S.n14293 S.n14292 0.001
R53746 S.n13579 S.n13578 0.001
R53747 S.n13314 S.n13313 0.001
R53748 S.n12607 S.n12606 0.001
R53749 S.n12326 S.n12325 0.001
R53750 S.n11613 S.n11612 0.001
R53751 S.n11312 S.n11311 0.001
R53752 S.n10606 S.n10605 0.001
R53753 S.n10289 S.n10288 0.001
R53754 S.n9577 S.n9576 0.001
R53755 S.n9240 S.n9239 0.001
R53756 S.n8535 S.n8534 0.001
R53757 S.n8182 S.n8181 0.001
R53758 S.n7471 S.n7470 0.001
R53759 S.n7098 S.n7097 0.001
R53760 S.n6394 S.n6393 0.001
R53761 S.n6005 S.n6004 0.001
R53762 S.n5294 S.n5293 0.001
R53763 S.n4885 S.n4884 0.001
R53764 S.n4181 S.n4180 0.001
R53765 S.n1445 S.n1444 0.001
R53766 S.n2626 S.n2625 0.001
R53767 S.n22365 S.n22364 0.001
R53768 S.n22689 S.n22688 0.001
R53769 S.n21653 S.n21652 0.001
R53770 S.n21275 S.n21274 0.001
R53771 S.n20506 S.n20505 0.001
R53772 S.n20859 S.n20858 0.001
R53773 S.n19895 S.n19894 0.001
R53774 S.n19788 S.n19787 0.001
R53775 S.n19041 S.n19040 0.001
R53776 S.n18916 S.n18915 0.001
R53777 S.n18175 S.n18174 0.001
R53778 S.n18033 S.n18032 0.001
R53779 S.n17286 S.n17285 0.001
R53780 S.n17124 S.n17123 0.001
R53781 S.n16384 S.n16383 0.001
R53782 S.n16206 S.n16205 0.001
R53783 S.n15460 S.n15459 0.001
R53784 S.n15262 S.n15261 0.001
R53785 S.n14523 S.n14522 0.001
R53786 S.n14309 S.n14308 0.001
R53787 S.n13564 S.n13563 0.001
R53788 S.n13330 S.n13329 0.001
R53789 S.n12592 S.n12591 0.001
R53790 S.n12342 S.n12341 0.001
R53791 S.n11598 S.n11597 0.001
R53792 S.n11328 S.n11327 0.001
R53793 S.n10591 S.n10590 0.001
R53794 S.n10305 S.n10304 0.001
R53795 S.n9562 S.n9561 0.001
R53796 S.n9256 S.n9255 0.001
R53797 S.n8520 S.n8519 0.001
R53798 S.n8198 S.n8197 0.001
R53799 S.n7456 S.n7455 0.001
R53800 S.n7114 S.n7113 0.001
R53801 S.n6379 S.n6378 0.001
R53802 S.n6021 S.n6020 0.001
R53803 S.n5279 S.n5278 0.001
R53804 S.n4901 S.n4900 0.001
R53805 S.n4166 S.n4165 0.001
R53806 S.n3773 S.n3772 0.001
R53807 S.n3040 S.n3039 0.001
R53808 S.n896 S.n895 0.001
R53809 S.n1978 S.n1977 0.001
R53810 S.n22729 S.n22728 0.001
R53811 S.n21309 S.n21308 0.001
R53812 S.n21208 S.n21207 0.001
R53813 S.n20486 S.n20485 0.001
R53814 S.n20389 S.n20388 0.001
R53815 S.n19875 S.n19874 0.001
R53816 S.n20262 S.n20261 0.001
R53817 S.n19021 S.n19020 0.001
R53818 S.n19394 S.n19393 0.001
R53819 S.n18155 S.n18154 0.001
R53820 S.n18507 S.n18506 0.001
R53821 S.n17266 S.n17265 0.001
R53822 S.n17607 S.n17606 0.001
R53823 S.n16364 S.n16363 0.001
R53824 S.n16684 S.n16683 0.001
R53825 S.n15440 S.n15439 0.001
R53826 S.n15749 S.n15748 0.001
R53827 S.n14503 S.n14502 0.001
R53828 S.n14791 S.n14790 0.001
R53829 S.n13544 S.n13543 0.001
R53830 S.n13821 S.n13820 0.001
R53831 S.n12572 S.n12571 0.001
R53832 S.n12828 S.n12827 0.001
R53833 S.n11578 S.n11577 0.001
R53834 S.n11823 S.n11822 0.001
R53835 S.n10571 S.n10570 0.001
R53836 S.n10795 S.n10794 0.001
R53837 S.n9542 S.n9541 0.001
R53838 S.n9755 S.n9754 0.001
R53839 S.n8500 S.n8499 0.001
R53840 S.n8692 S.n8691 0.001
R53841 S.n7436 S.n7435 0.001
R53842 S.n7617 S.n7616 0.001
R53843 S.n6359 S.n6358 0.001
R53844 S.n6519 S.n6518 0.001
R53845 S.n5259 S.n5258 0.001
R53846 S.n5408 S.n5407 0.001
R53847 S.n4146 S.n4145 0.001
R53848 S.n4274 S.n4273 0.001
R53849 S.n3020 S.n3019 0.001
R53850 S.n3138 S.n3137 0.001
R53851 S.n1859 S.n1858 0.001
R53852 S.n874 S.n873 0.001
R53853 S.n798 S.n797 0.001
R53854 S.n22346 S.n22345 0.001
R53855 S.n22708 S.n22707 0.001
R53856 S.n21340 S.n21339 0.001
R53857 S.n21256 S.n21255 0.001
R53858 S.n20434 S.n20433 0.001
R53859 S.n20840 S.n20839 0.001
R53860 S.n19800 S.n19799 0.001
R53861 S.n20205 S.n20204 0.001
R53862 S.n18928 S.n18927 0.001
R53863 S.n19335 S.n19334 0.001
R53864 S.n18045 S.n18044 0.001
R53865 S.n18453 S.n18452 0.001
R53866 S.n17136 S.n17135 0.001
R53867 S.n17548 S.n17547 0.001
R53868 S.n16218 S.n16217 0.001
R53869 S.n16630 S.n16629 0.001
R53870 S.n15274 S.n15273 0.001
R53871 S.n15690 S.n15689 0.001
R53872 S.n14321 S.n14320 0.001
R53873 S.n14737 S.n14736 0.001
R53874 S.n13342 S.n13341 0.001
R53875 S.n13762 S.n13761 0.001
R53876 S.n12354 S.n12353 0.001
R53877 S.n12774 S.n12773 0.001
R53878 S.n11340 S.n11339 0.001
R53879 S.n11764 S.n11763 0.001
R53880 S.n10317 S.n10316 0.001
R53881 S.n10741 S.n10740 0.001
R53882 S.n9268 S.n9267 0.001
R53883 S.n9696 S.n9695 0.001
R53884 S.n8210 S.n8209 0.001
R53885 S.n8638 S.n8637 0.001
R53886 S.n7126 S.n7125 0.001
R53887 S.n7558 S.n7557 0.001
R53888 S.n6033 S.n6032 0.001
R53889 S.n6465 S.n6464 0.001
R53890 S.n4913 S.n4912 0.001
R53891 S.n5349 S.n5348 0.001
R53892 S.n3785 S.n3784 0.001
R53893 S.n4220 S.n4219 0.001
R53894 S.n2638 S.n2637 0.001
R53895 S.n3079 S.n3078 0.001
R53896 S.n1877 S.n1876 0.001
R53897 S.n1922 S.n1921 0.001
R53898 S.n401 S.n400 0.001
R53899 S.n2130 S.n2129 0.001
R53900 S.n18472 S.n18471 0.001
R53901 S.n17164 S.n17163 0.001
R53902 S.n17756 S.n17755 0.001
R53903 S.n16264 S.n16263 0.001
R53904 S.n16829 S.n16828 0.001
R53905 S.n15340 S.n15339 0.001
R53906 S.n15894 S.n15893 0.001
R53907 S.n14403 S.n14402 0.001
R53908 S.n14936 S.n14935 0.001
R53909 S.n13444 S.n13443 0.001
R53910 S.n13966 S.n13965 0.001
R53911 S.n12472 S.n12471 0.001
R53912 S.n12973 S.n12972 0.001
R53913 S.n11478 S.n11477 0.001
R53914 S.n11968 S.n11967 0.001
R53915 S.n10471 S.n10470 0.001
R53916 S.n10940 S.n10939 0.001
R53917 S.n9442 S.n9441 0.001
R53918 S.n9900 S.n9899 0.001
R53919 S.n8400 S.n8399 0.001
R53920 S.n8837 S.n8836 0.001
R53921 S.n7336 S.n7335 0.001
R53922 S.n7762 S.n7761 0.001
R53923 S.n6259 S.n6258 0.001
R53924 S.n6664 S.n6663 0.001
R53925 S.n5159 S.n5158 0.001
R53926 S.n5554 S.n5553 0.001
R53927 S.n4047 S.n4046 0.001
R53928 S.n4419 S.n4418 0.001
R53929 S.n2920 S.n2919 0.001
R53930 S.n3282 S.n3281 0.001
R53931 S.n1751 S.n1750 0.001
R53932 S.n13 S.n12 0.001
R53933 S.n19358 S.n19357 0.001
R53934 S.n18072 S.n18071 0.001
R53935 S.n18619 S.n18618 0.001
R53936 S.n17183 S.n17182 0.001
R53937 S.n17719 S.n17718 0.001
R53938 S.n16281 S.n16280 0.001
R53939 S.n16792 S.n16791 0.001
R53940 S.n15357 S.n15356 0.001
R53941 S.n15857 S.n15856 0.001
R53942 S.n14420 S.n14419 0.001
R53943 S.n14899 S.n14898 0.001
R53944 S.n13461 S.n13460 0.001
R53945 S.n13929 S.n13928 0.001
R53946 S.n12489 S.n12488 0.001
R53947 S.n12936 S.n12935 0.001
R53948 S.n11495 S.n11494 0.001
R53949 S.n11931 S.n11930 0.001
R53950 S.n10488 S.n10487 0.001
R53951 S.n10903 S.n10902 0.001
R53952 S.n9459 S.n9458 0.001
R53953 S.n9863 S.n9862 0.001
R53954 S.n8417 S.n8416 0.001
R53955 S.n8800 S.n8799 0.001
R53956 S.n7353 S.n7352 0.001
R53957 S.n7725 S.n7724 0.001
R53958 S.n6276 S.n6275 0.001
R53959 S.n6627 S.n6626 0.001
R53960 S.n5176 S.n5175 0.001
R53961 S.n5517 S.n5516 0.001
R53962 S.n4064 S.n4063 0.001
R53963 S.n4382 S.n4381 0.001
R53964 S.n2937 S.n2936 0.001
R53965 S.n3245 S.n3244 0.001
R53966 S.n1769 S.n1768 0.001
R53967 S.n1791 S.n1790 0.001
R53968 S.n2061 S.n2060 0.001
R53969 S.n416 S.n415 0.001
R53970 S.n829 S.n828 0.001
R53971 S.n3222 S.n3221 0.001
R53972 S.n4358 S.n4357 0.001
R53973 S.n5493 S.n5492 0.001
R53974 S.n6603 S.n6602 0.001
R53975 S.n7701 S.n7700 0.001
R53976 S.n8776 S.n8775 0.001
R53977 S.n9839 S.n9838 0.001
R53978 S.n10879 S.n10878 0.001
R53979 S.n11907 S.n11906 0.001
R53980 S.n12912 S.n12911 0.001
R53981 S.n13905 S.n13904 0.001
R53982 S.n14875 S.n14874 0.001
R53983 S.n15833 S.n15832 0.001
R53984 S.n16768 S.n16767 0.001
R53985 S.n17691 S.n17690 0.001
R53986 S.n18591 S.n18590 0.001
R53987 S.n19481 S.n19480 0.001
R53988 S.n20227 S.n20226 0.001
R53989 S.n18956 S.n18955 0.001
R53990 S.n18091 S.n18090 0.001
R53991 S.n17202 S.n17201 0.001
R53992 S.n16300 S.n16299 0.001
R53993 S.n15376 S.n15375 0.001
R53994 S.n14439 S.n14438 0.001
R53995 S.n13480 S.n13479 0.001
R53996 S.n12508 S.n12507 0.001
R53997 S.n11514 S.n11513 0.001
R53998 S.n10507 S.n10506 0.001
R53999 S.n9478 S.n9477 0.001
R54000 S.n8436 S.n8435 0.001
R54001 S.n7372 S.n7371 0.001
R54002 S.n6295 S.n6294 0.001
R54003 S.n5195 S.n5194 0.001
R54004 S.n4083 S.n4082 0.001
R54005 S.n2956 S.n2955 0.001
R54006 S.n2033 S.n2032 0.001
R54007 S.n754 S.n753 0.001
R54008 S.n1325 S.n1324 0.001
R54009 S.n20419 S.n20418 0.001
R54010 S.n19836 S.n19835 0.001
R54011 S.n20315 S.n20314 0.001
R54012 S.n18984 S.n18983 0.001
R54013 S.n19443 S.n19442 0.001
R54014 S.n18119 S.n18118 0.001
R54015 S.n18556 S.n18555 0.001
R54016 S.n17230 S.n17229 0.001
R54017 S.n17656 S.n17655 0.001
R54018 S.n16328 S.n16327 0.001
R54019 S.n16733 S.n16732 0.001
R54020 S.n15404 S.n15403 0.001
R54021 S.n15798 S.n15797 0.001
R54022 S.n14467 S.n14466 0.001
R54023 S.n14840 S.n14839 0.001
R54024 S.n13508 S.n13507 0.001
R54025 S.n13870 S.n13869 0.001
R54026 S.n12536 S.n12535 0.001
R54027 S.n12877 S.n12876 0.001
R54028 S.n11542 S.n11541 0.001
R54029 S.n11872 S.n11871 0.001
R54030 S.n10535 S.n10534 0.001
R54031 S.n10844 S.n10843 0.001
R54032 S.n9506 S.n9505 0.001
R54033 S.n9804 S.n9803 0.001
R54034 S.n8464 S.n8463 0.001
R54035 S.n8741 S.n8740 0.001
R54036 S.n7400 S.n7399 0.001
R54037 S.n7666 S.n7665 0.001
R54038 S.n6323 S.n6322 0.001
R54039 S.n6568 S.n6567 0.001
R54040 S.n5223 S.n5222 0.001
R54041 S.n5458 S.n5457 0.001
R54042 S.n4111 S.n4110 0.001
R54043 S.n4323 S.n4322 0.001
R54044 S.n2984 S.n2983 0.001
R54045 S.n3186 S.n3185 0.001
R54046 S.n1821 S.n1820 0.001
R54047 S.n2000 S.n1999 0.001
R54048 S.n778 S.n777 0.001
R54049 S.n1842 S.n1841 0.001
R54050 S.n3161 S.n3160 0.001
R54051 S.n2998 S.n2997 0.001
R54052 S.n4298 S.n4297 0.001
R54053 S.n4125 S.n4124 0.001
R54054 S.n5432 S.n5431 0.001
R54055 S.n5237 S.n5236 0.001
R54056 S.n6543 S.n6542 0.001
R54057 S.n6337 S.n6336 0.001
R54058 S.n7641 S.n7640 0.001
R54059 S.n7414 S.n7413 0.001
R54060 S.n8716 S.n8715 0.001
R54061 S.n8478 S.n8477 0.001
R54062 S.n9779 S.n9778 0.001
R54063 S.n9520 S.n9519 0.001
R54064 S.n10819 S.n10818 0.001
R54065 S.n10549 S.n10548 0.001
R54066 S.n11847 S.n11846 0.001
R54067 S.n11556 S.n11555 0.001
R54068 S.n12852 S.n12851 0.001
R54069 S.n12550 S.n12549 0.001
R54070 S.n13845 S.n13844 0.001
R54071 S.n13522 S.n13521 0.001
R54072 S.n14815 S.n14814 0.001
R54073 S.n14481 S.n14480 0.001
R54074 S.n15773 S.n15772 0.001
R54075 S.n15418 S.n15417 0.001
R54076 S.n16708 S.n16707 0.001
R54077 S.n16342 S.n16341 0.001
R54078 S.n17631 S.n17630 0.001
R54079 S.n17244 S.n17243 0.001
R54080 S.n18531 S.n18530 0.001
R54081 S.n18133 S.n18132 0.001
R54082 S.n19418 S.n19417 0.001
R54083 S.n18999 S.n18998 0.001
R54084 S.n20290 S.n20289 0.001
R54085 S.n19853 S.n19852 0.001
R54086 S.n20361 S.n20360 0.001
R54087 S.n20464 S.n20463 0.001
R54088 S.n21237 S.n21236 0.001
R54089 S.n853 S.n852 0.001
R54090 S.n2094 S.n2093 0.001
R54091 S.n738 S.n737 0.001
R54092 S.n721 S.n720 0.001
R54093 S.n369 S.n368 0.001
R54094 S.n2189 S.n2188 0.001
R54095 S.n16649 S.n16648 0.001
R54096 S.n15302 S.n15301 0.001
R54097 S.n15959 S.n15958 0.001
R54098 S.n14367 S.n14366 0.001
R54099 S.n14997 S.n14996 0.001
R54100 S.n13408 S.n13407 0.001
R54101 S.n14027 S.n14026 0.001
R54102 S.n12436 S.n12435 0.001
R54103 S.n13034 S.n13033 0.001
R54104 S.n11442 S.n11441 0.001
R54105 S.n12029 S.n12028 0.001
R54106 S.n10435 S.n10434 0.001
R54107 S.n11001 S.n11000 0.001
R54108 S.n9406 S.n9405 0.001
R54109 S.n9961 S.n9960 0.001
R54110 S.n8364 S.n8363 0.001
R54111 S.n8898 S.n8897 0.001
R54112 S.n7300 S.n7299 0.001
R54113 S.n7823 S.n7822 0.001
R54114 S.n6223 S.n6222 0.001
R54115 S.n6725 S.n6724 0.001
R54116 S.n5123 S.n5122 0.001
R54117 S.n5615 S.n5614 0.001
R54118 S.n4011 S.n4010 0.001
R54119 S.n4480 S.n4479 0.001
R54120 S.n2884 S.n2883 0.001
R54121 S.n3342 S.n3341 0.001
R54122 S.n1714 S.n1713 0.001
R54123 S.n60 S.n59 0.001
R54124 S.n17571 S.n17570 0.001
R54125 S.n16245 S.n16244 0.001
R54126 S.n16857 S.n16856 0.001
R54127 S.n15321 S.n15320 0.001
R54128 S.n15922 S.n15921 0.001
R54129 S.n14384 S.n14383 0.001
R54130 S.n14960 S.n14959 0.001
R54131 S.n13425 S.n13424 0.001
R54132 S.n13990 S.n13989 0.001
R54133 S.n12453 S.n12452 0.001
R54134 S.n12997 S.n12996 0.001
R54135 S.n11459 S.n11458 0.001
R54136 S.n11992 S.n11991 0.001
R54137 S.n10452 S.n10451 0.001
R54138 S.n10964 S.n10963 0.001
R54139 S.n9423 S.n9422 0.001
R54140 S.n9924 S.n9923 0.001
R54141 S.n8381 S.n8380 0.001
R54142 S.n8861 S.n8860 0.001
R54143 S.n7317 S.n7316 0.001
R54144 S.n7786 S.n7785 0.001
R54145 S.n6240 S.n6239 0.001
R54146 S.n6688 S.n6687 0.001
R54147 S.n5140 S.n5139 0.001
R54148 S.n5578 S.n5577 0.001
R54149 S.n4028 S.n4027 0.001
R54150 S.n4443 S.n4442 0.001
R54151 S.n2901 S.n2900 0.001
R54152 S.n3305 S.n3304 0.001
R54153 S.n1732 S.n1731 0.001
R54154 S.n2152 S.n2151 0.001
R54155 S.n703 S.n702 0.001
R54156 S.n686 S.n685 0.001
R54157 S.n337 S.n336 0.001
R54158 S.n2248 S.n2247 0.001
R54159 S.n14756 S.n14755 0.001
R54160 S.n13370 S.n13369 0.001
R54161 S.n14092 S.n14091 0.001
R54162 S.n12400 S.n12399 0.001
R54163 S.n13095 S.n13094 0.001
R54164 S.n11406 S.n11405 0.001
R54165 S.n12090 S.n12089 0.001
R54166 S.n10399 S.n10398 0.001
R54167 S.n11062 S.n11061 0.001
R54168 S.n9370 S.n9369 0.001
R54169 S.n10022 S.n10021 0.001
R54170 S.n8328 S.n8327 0.001
R54171 S.n8959 S.n8958 0.001
R54172 S.n7264 S.n7263 0.001
R54173 S.n7884 S.n7883 0.001
R54174 S.n6187 S.n6186 0.001
R54175 S.n6786 S.n6785 0.001
R54176 S.n5087 S.n5086 0.001
R54177 S.n5676 S.n5675 0.001
R54178 S.n3975 S.n3974 0.001
R54179 S.n4541 S.n4540 0.001
R54180 S.n2848 S.n2847 0.001
R54181 S.n3402 S.n3401 0.001
R54182 S.n1677 S.n1676 0.001
R54183 S.n92 S.n91 0.001
R54184 S.n15713 S.n15712 0.001
R54185 S.n14348 S.n14347 0.001
R54186 S.n15025 S.n15024 0.001
R54187 S.n13389 S.n13388 0.001
R54188 S.n14055 S.n14054 0.001
R54189 S.n12417 S.n12416 0.001
R54190 S.n13058 S.n13057 0.001
R54191 S.n11423 S.n11422 0.001
R54192 S.n12053 S.n12052 0.001
R54193 S.n10416 S.n10415 0.001
R54194 S.n11025 S.n11024 0.001
R54195 S.n9387 S.n9386 0.001
R54196 S.n9985 S.n9984 0.001
R54197 S.n8345 S.n8344 0.001
R54198 S.n8922 S.n8921 0.001
R54199 S.n7281 S.n7280 0.001
R54200 S.n7847 S.n7846 0.001
R54201 S.n6204 S.n6203 0.001
R54202 S.n6749 S.n6748 0.001
R54203 S.n5104 S.n5103 0.001
R54204 S.n5639 S.n5638 0.001
R54205 S.n3992 S.n3991 0.001
R54206 S.n4504 S.n4503 0.001
R54207 S.n2865 S.n2864 0.001
R54208 S.n3365 S.n3364 0.001
R54209 S.n1695 S.n1694 0.001
R54210 S.n2211 S.n2210 0.001
R54211 S.n668 S.n667 0.001
R54212 S.n651 S.n650 0.001
R54213 S.n305 S.n304 0.001
R54214 S.n2307 S.n2306 0.001
R54215 S.n12793 S.n12792 0.001
R54216 S.n11368 S.n11367 0.001
R54217 S.n12155 S.n12154 0.001
R54218 S.n10363 S.n10362 0.001
R54219 S.n11123 S.n11122 0.001
R54220 S.n9334 S.n9333 0.001
R54221 S.n10083 S.n10082 0.001
R54222 S.n8292 S.n8291 0.001
R54223 S.n9020 S.n9019 0.001
R54224 S.n7228 S.n7227 0.001
R54225 S.n7945 S.n7944 0.001
R54226 S.n6151 S.n6150 0.001
R54227 S.n6847 S.n6846 0.001
R54228 S.n5051 S.n5050 0.001
R54229 S.n5737 S.n5736 0.001
R54230 S.n3939 S.n3938 0.001
R54231 S.n4602 S.n4601 0.001
R54232 S.n2812 S.n2811 0.001
R54233 S.n3462 S.n3461 0.001
R54234 S.n1640 S.n1639 0.001
R54235 S.n124 S.n123 0.001
R54236 S.n13785 S.n13784 0.001
R54237 S.n12381 S.n12380 0.001
R54238 S.n13123 S.n13122 0.001
R54239 S.n11387 S.n11386 0.001
R54240 S.n12118 S.n12117 0.001
R54241 S.n10380 S.n10379 0.001
R54242 S.n11086 S.n11085 0.001
R54243 S.n9351 S.n9350 0.001
R54244 S.n10046 S.n10045 0.001
R54245 S.n8309 S.n8308 0.001
R54246 S.n8983 S.n8982 0.001
R54247 S.n7245 S.n7244 0.001
R54248 S.n7908 S.n7907 0.001
R54249 S.n6168 S.n6167 0.001
R54250 S.n6810 S.n6809 0.001
R54251 S.n5068 S.n5067 0.001
R54252 S.n5700 S.n5699 0.001
R54253 S.n3956 S.n3955 0.001
R54254 S.n4565 S.n4564 0.001
R54255 S.n2829 S.n2828 0.001
R54256 S.n3425 S.n3424 0.001
R54257 S.n1658 S.n1657 0.001
R54258 S.n2270 S.n2269 0.001
R54259 S.n633 S.n632 0.001
R54260 S.n616 S.n615 0.001
R54261 S.n273 S.n272 0.001
R54262 S.n2366 S.n2365 0.001
R54263 S.n10760 S.n10759 0.001
R54264 S.n9296 S.n9295 0.001
R54265 S.n10148 S.n10147 0.001
R54266 S.n8256 S.n8255 0.001
R54267 S.n9081 S.n9080 0.001
R54268 S.n7192 S.n7191 0.001
R54269 S.n8006 S.n8005 0.001
R54270 S.n6115 S.n6114 0.001
R54271 S.n6908 S.n6907 0.001
R54272 S.n5015 S.n5014 0.001
R54273 S.n5798 S.n5797 0.001
R54274 S.n3903 S.n3902 0.001
R54275 S.n4663 S.n4662 0.001
R54276 S.n2776 S.n2775 0.001
R54277 S.n3522 S.n3521 0.001
R54278 S.n1603 S.n1602 0.001
R54279 S.n1011 S.n1010 0.001
R54280 S.n11787 S.n11786 0.001
R54281 S.n10344 S.n10343 0.001
R54282 S.n11151 S.n11150 0.001
R54283 S.n9315 S.n9314 0.001
R54284 S.n10111 S.n10110 0.001
R54285 S.n8273 S.n8272 0.001
R54286 S.n9044 S.n9043 0.001
R54287 S.n7209 S.n7208 0.001
R54288 S.n7969 S.n7968 0.001
R54289 S.n6132 S.n6131 0.001
R54290 S.n6871 S.n6870 0.001
R54291 S.n5032 S.n5031 0.001
R54292 S.n5761 S.n5760 0.001
R54293 S.n3920 S.n3919 0.001
R54294 S.n4626 S.n4625 0.001
R54295 S.n2793 S.n2792 0.001
R54296 S.n3485 S.n3484 0.001
R54297 S.n1621 S.n1620 0.001
R54298 S.n2329 S.n2328 0.001
R54299 S.n598 S.n597 0.001
R54300 S.n581 S.n580 0.001
R54301 S.n244 S.n243 0.001
R54302 S.n2425 S.n2424 0.001
R54303 S.n8657 S.n8656 0.001
R54304 S.n7154 S.n7153 0.001
R54305 S.n8071 S.n8070 0.001
R54306 S.n6079 S.n6078 0.001
R54307 S.n6969 S.n6968 0.001
R54308 S.n4979 S.n4978 0.001
R54309 S.n5859 S.n5858 0.001
R54310 S.n3867 S.n3866 0.001
R54311 S.n4724 S.n4723 0.001
R54312 S.n2740 S.n2739 0.001
R54313 S.n3582 S.n3581 0.001
R54314 S.n1566 S.n1565 0.001
R54315 S.n1043 S.n1042 0.001
R54316 S.n9719 S.n9718 0.001
R54317 S.n8237 S.n8236 0.001
R54318 S.n9109 S.n9108 0.001
R54319 S.n7173 S.n7172 0.001
R54320 S.n8034 S.n8033 0.001
R54321 S.n6096 S.n6095 0.001
R54322 S.n6932 S.n6931 0.001
R54323 S.n4996 S.n4995 0.001
R54324 S.n5822 S.n5821 0.001
R54325 S.n3884 S.n3883 0.001
R54326 S.n4687 S.n4686 0.001
R54327 S.n2757 S.n2756 0.001
R54328 S.n3545 S.n3544 0.001
R54329 S.n1584 S.n1583 0.001
R54330 S.n2388 S.n2387 0.001
R54331 S.n563 S.n562 0.001
R54332 S.n546 S.n545 0.001
R54333 S.n209 S.n208 0.001
R54334 S.n2484 S.n2483 0.001
R54335 S.n6484 S.n6483 0.001
R54336 S.n4941 S.n4940 0.001
R54337 S.n5924 S.n5923 0.001
R54338 S.n3831 S.n3830 0.001
R54339 S.n4785 S.n4784 0.001
R54340 S.n2704 S.n2703 0.001
R54341 S.n3642 S.n3641 0.001
R54342 S.n1529 S.n1528 0.001
R54343 S.n1075 S.n1074 0.001
R54344 S.n7581 S.n7580 0.001
R54345 S.n6060 S.n6059 0.001
R54346 S.n6997 S.n6996 0.001
R54347 S.n4960 S.n4959 0.001
R54348 S.n5887 S.n5886 0.001
R54349 S.n3848 S.n3847 0.001
R54350 S.n4748 S.n4747 0.001
R54351 S.n2721 S.n2720 0.001
R54352 S.n3605 S.n3604 0.001
R54353 S.n1547 S.n1546 0.001
R54354 S.n2447 S.n2446 0.001
R54355 S.n528 S.n527 0.001
R54356 S.n511 S.n510 0.001
R54357 S.n177 S.n176 0.001
R54358 S.n2543 S.n2542 0.001
R54359 S.n4239 S.n4238 0.001
R54360 S.n2666 S.n2665 0.001
R54361 S.n3706 S.n3705 0.001
R54362 S.n1492 S.n1491 0.001
R54363 S.n1107 S.n1106 0.001
R54364 S.n5372 S.n5371 0.001
R54365 S.n3812 S.n3811 0.001
R54366 S.n4813 S.n4812 0.001
R54367 S.n2685 S.n2684 0.001
R54368 S.n3669 S.n3668 0.001
R54369 S.n1510 S.n1509 0.001
R54370 S.n2506 S.n2505 0.001
R54371 S.n493 S.n492 0.001
R54372 S.n476 S.n475 0.001
R54373 S.n145 S.n144 0.001
R54374 S.n1945 S.n1944 0.001
R54375 S.n1145 S.n1144 0.001
R54376 S.n3102 S.n3101 0.001
R54377 S.n1473 S.n1472 0.001
R54378 S.n2569 S.n2568 0.001
R54379 S.n458 S.n457 0.001
R54380 S.n442 S.n441 0.001
R54381 S.n932 S.n931 0.001
R54382 S.n22760 S.n22759 0.001
R54383 S.n21323 S.n21322 0.001
R54384 S.n44 S.n43 0.001
R54385 S.n43 S.n38 0.001
R54386 S.n22286 S.n22285 0.001
R54387 S.n21293 S.n21292 0.001
R54388 S.n20449 S.n20448 0.001
R54389 S.n19811 S.n19810 0.001
R54390 S.n18941 S.n18940 0.001
R54391 S.n18056 S.n18055 0.001
R54392 S.n17149 S.n17148 0.001
R54393 S.n16229 S.n16228 0.001
R54394 S.n15287 S.n15286 0.001
R54395 S.n14332 S.n14331 0.001
R54396 S.n13355 S.n13354 0.001
R54397 S.n12365 S.n12364 0.001
R54398 S.n11353 S.n11352 0.001
R54399 S.n10328 S.n10327 0.001
R54400 S.n9281 S.n9280 0.001
R54401 S.n8221 S.n8220 0.001
R54402 S.n7139 S.n7138 0.001
R54403 S.n6044 S.n6043 0.001
R54404 S.n4926 S.n4925 0.001
R54405 S.n3796 S.n3795 0.001
R54406 S.n2651 S.n2650 0.001
R54407 S.n1457 S.n1456 0.001
R54408 S.n429 S.n428 0.001
R54409 S.n20339 S.t262 0.001
R54410 S.t209 S.n20186 0.001
R54411 S.t209 S.n20189 0.001
R54412 S.t7 S.n21136 0.001
R54413 S.t7 S.n21139 0.001
R54414 S.t9 S.n22643 0.001
R54415 S.t9 S.n22646 0.001
R54416 S.t88 S.n22016 0.001
R54417 S.t88 S.n22013 0.001
R54418 S.n22013 S.n22010 0.001
R54419 S.t100 S.n21620 0.001
R54420 S.t100 S.n21623 0.001
R54421 S.t105 S.n21945 0.001
R54422 S.t105 S.n21948 0.001
R54423 S.t64 S.n20797 0.001
R54424 S.t64 S.n20800 0.001
R54425 S.n21142 S.t7 0.001
R54426 S.n21172 S.n21144 0.001
R54427 S.t9 S.n22659 0.001
R54428 S.t9 S.n22662 0.001
R54429 S.t88 S.n22001 0.001
R54430 S.t88 S.n21998 0.001
R54431 S.n21998 S.n21995 0.001
R54432 S.t100 S.n21641 0.001
R54433 S.t100 S.n21644 0.001
R54434 S.t105 S.n21965 0.001
R54435 S.t105 S.n21968 0.001
R54436 S.t64 S.n20821 0.001
R54437 S.t64 S.n20824 0.001
R54438 S.n20344 S.n20339 0.001
R54439 S.n19499 S.t21 0.001
R54440 S.t150 S.n19316 0.001
R54441 S.t150 S.n19319 0.001
R54442 S.t262 S.n19539 0.001
R54443 S.t262 S.n19536 0.001
R54444 S.n19536 S.n19533 0.001
R54445 S.t9 S.n22627 0.001
R54446 S.t9 S.n22630 0.001
R54447 S.t88 S.n22031 0.001
R54448 S.t88 S.n22028 0.001
R54449 S.n22028 S.n22025 0.001
R54450 S.t100 S.n21604 0.001
R54451 S.t100 S.n21607 0.001
R54452 S.t105 S.n21930 0.001
R54453 S.t105 S.n21933 0.001
R54454 S.t64 S.n20781 0.001
R54455 S.t64 S.n20784 0.001
R54456 S.t7 S.n21120 0.001
R54457 S.t7 S.n21123 0.001
R54458 S.t209 S.n20170 0.001
R54459 S.t209 S.n20173 0.001
R54460 S.n19504 S.n19499 0.001
R54461 S.n18642 S.t77 0.001
R54462 S.t79 S.n18434 0.001
R54463 S.t79 S.n18437 0.001
R54464 S.t21 S.n18682 0.001
R54465 S.t21 S.n18679 0.001
R54466 S.n18679 S.n18676 0.001
R54467 S.t9 S.n22611 0.001
R54468 S.t9 S.n22614 0.001
R54469 S.t88 S.n22046 0.001
R54470 S.t88 S.n22043 0.001
R54471 S.n22043 S.n22040 0.001
R54472 S.t100 S.n21588 0.001
R54473 S.t100 S.n21591 0.001
R54474 S.t105 S.n21915 0.001
R54475 S.t105 S.n21918 0.001
R54476 S.t64 S.n20765 0.001
R54477 S.t64 S.n20768 0.001
R54478 S.t7 S.n21105 0.001
R54479 S.t7 S.n21108 0.001
R54480 S.t209 S.n20154 0.001
R54481 S.t209 S.n20157 0.001
R54482 S.t262 S.n19554 0.001
R54483 S.t262 S.n19551 0.001
R54484 S.n19551 S.n19548 0.001
R54485 S.t150 S.n19300 0.001
R54486 S.t150 S.n19303 0.001
R54487 S.n18647 S.n18642 0.001
R54488 S.n17774 S.t169 0.001
R54489 S.t218 S.n17529 0.001
R54490 S.t218 S.n17532 0.001
R54491 S.t77 S.n17814 0.001
R54492 S.t77 S.n17811 0.001
R54493 S.n17811 S.n17808 0.001
R54494 S.t9 S.n22595 0.001
R54495 S.t9 S.n22598 0.001
R54496 S.t88 S.n22061 0.001
R54497 S.t88 S.n22058 0.001
R54498 S.n22058 S.n22055 0.001
R54499 S.t100 S.n21572 0.001
R54500 S.t100 S.n21575 0.001
R54501 S.t105 S.n21900 0.001
R54502 S.t105 S.n21903 0.001
R54503 S.t64 S.n20749 0.001
R54504 S.t64 S.n20752 0.001
R54505 S.t7 S.n21090 0.001
R54506 S.t7 S.n21093 0.001
R54507 S.t209 S.n20138 0.001
R54508 S.t209 S.n20141 0.001
R54509 S.t262 S.n19569 0.001
R54510 S.t262 S.n19566 0.001
R54511 S.n19566 S.n19563 0.001
R54512 S.t150 S.n19284 0.001
R54513 S.t150 S.n19287 0.001
R54514 S.t21 S.n18697 0.001
R54515 S.t21 S.n18694 0.001
R54516 S.n18694 S.n18691 0.001
R54517 S.t79 S.n18418 0.001
R54518 S.t79 S.n18421 0.001
R54519 S.n17779 S.n17774 0.001
R54520 S.n16880 S.t187 0.001
R54521 S.t167 S.n16611 0.001
R54522 S.t167 S.n16614 0.001
R54523 S.t169 S.n16920 0.001
R54524 S.t169 S.n16917 0.001
R54525 S.n16917 S.n16914 0.001
R54526 S.t9 S.n22579 0.001
R54527 S.t9 S.n22582 0.001
R54528 S.t88 S.n22076 0.001
R54529 S.t88 S.n22073 0.001
R54530 S.n22073 S.n22070 0.001
R54531 S.t100 S.n21556 0.001
R54532 S.t100 S.n21559 0.001
R54533 S.t105 S.n21885 0.001
R54534 S.t105 S.n21888 0.001
R54535 S.t64 S.n20733 0.001
R54536 S.t64 S.n20736 0.001
R54537 S.t7 S.n21075 0.001
R54538 S.t7 S.n21078 0.001
R54539 S.t209 S.n20122 0.001
R54540 S.t209 S.n20125 0.001
R54541 S.t262 S.n19584 0.001
R54542 S.t262 S.n19581 0.001
R54543 S.n19581 S.n19578 0.001
R54544 S.t150 S.n19268 0.001
R54545 S.t150 S.n19271 0.001
R54546 S.t21 S.n18712 0.001
R54547 S.t21 S.n18709 0.001
R54548 S.n18709 S.n18706 0.001
R54549 S.t79 S.n18402 0.001
R54550 S.t79 S.n18405 0.001
R54551 S.t77 S.n17829 0.001
R54552 S.t77 S.n17826 0.001
R54553 S.n17826 S.n17823 0.001
R54554 S.t218 S.n17513 0.001
R54555 S.t218 S.n17516 0.001
R54556 S.n16885 S.n16880 0.001
R54557 S.n15977 S.t29 0.001
R54558 S.t60 S.n15671 0.001
R54559 S.t60 S.n15674 0.001
R54560 S.t187 S.n16017 0.001
R54561 S.t187 S.n16014 0.001
R54562 S.n16014 S.n16011 0.001
R54563 S.t9 S.n22563 0.001
R54564 S.t9 S.n22566 0.001
R54565 S.t88 S.n22091 0.001
R54566 S.t88 S.n22088 0.001
R54567 S.n22088 S.n22085 0.001
R54568 S.t100 S.n21540 0.001
R54569 S.t100 S.n21543 0.001
R54570 S.t105 S.n21870 0.001
R54571 S.t105 S.n21873 0.001
R54572 S.t64 S.n20717 0.001
R54573 S.t64 S.n20720 0.001
R54574 S.t7 S.n21060 0.001
R54575 S.t7 S.n21063 0.001
R54576 S.t209 S.n20106 0.001
R54577 S.t209 S.n20109 0.001
R54578 S.t262 S.n19599 0.001
R54579 S.t262 S.n19596 0.001
R54580 S.n19596 S.n19593 0.001
R54581 S.t150 S.n19252 0.001
R54582 S.t150 S.n19255 0.001
R54583 S.t21 S.n18727 0.001
R54584 S.t21 S.n18724 0.001
R54585 S.n18724 S.n18721 0.001
R54586 S.t79 S.n18386 0.001
R54587 S.t79 S.n18389 0.001
R54588 S.t77 S.n17844 0.001
R54589 S.t77 S.n17841 0.001
R54590 S.n17841 S.n17838 0.001
R54591 S.t218 S.n17497 0.001
R54592 S.t218 S.n17500 0.001
R54593 S.t169 S.n16935 0.001
R54594 S.t169 S.n16932 0.001
R54595 S.n16932 S.n16929 0.001
R54596 S.t167 S.n16595 0.001
R54597 S.t167 S.n16598 0.001
R54598 S.n15982 S.n15977 0.001
R54599 S.n15048 S.t102 0.001
R54600 S.t0 S.n14718 0.001
R54601 S.t0 S.n14721 0.001
R54602 S.t29 S.n15088 0.001
R54603 S.t29 S.n15085 0.001
R54604 S.n15085 S.n15082 0.001
R54605 S.t9 S.n22547 0.001
R54606 S.t9 S.n22550 0.001
R54607 S.t88 S.n22106 0.001
R54608 S.t88 S.n22103 0.001
R54609 S.n22103 S.n22100 0.001
R54610 S.t100 S.n21524 0.001
R54611 S.t100 S.n21527 0.001
R54612 S.t105 S.n21855 0.001
R54613 S.t105 S.n21858 0.001
R54614 S.t64 S.n20701 0.001
R54615 S.t64 S.n20704 0.001
R54616 S.t7 S.n21045 0.001
R54617 S.t7 S.n21048 0.001
R54618 S.t209 S.n20090 0.001
R54619 S.t209 S.n20093 0.001
R54620 S.t262 S.n19614 0.001
R54621 S.t262 S.n19611 0.001
R54622 S.n19611 S.n19608 0.001
R54623 S.t150 S.n19236 0.001
R54624 S.t150 S.n19239 0.001
R54625 S.t21 S.n18742 0.001
R54626 S.t21 S.n18739 0.001
R54627 S.n18739 S.n18736 0.001
R54628 S.t79 S.n18370 0.001
R54629 S.t79 S.n18373 0.001
R54630 S.t77 S.n17859 0.001
R54631 S.t77 S.n17856 0.001
R54632 S.n17856 S.n17853 0.001
R54633 S.t218 S.n17481 0.001
R54634 S.t218 S.n17484 0.001
R54635 S.t169 S.n16950 0.001
R54636 S.t169 S.n16947 0.001
R54637 S.n16947 S.n16944 0.001
R54638 S.t167 S.n16579 0.001
R54639 S.t167 S.n16582 0.001
R54640 S.t187 S.n16032 0.001
R54641 S.t187 S.n16029 0.001
R54642 S.n16029 S.n16026 0.001
R54643 S.t60 S.n15655 0.001
R54644 S.t60 S.n15658 0.001
R54645 S.n15053 S.n15048 0.001
R54646 S.n14110 S.t538 0.001
R54647 S.t73 S.n13743 0.001
R54648 S.t73 S.n13746 0.001
R54649 S.t102 S.n14150 0.001
R54650 S.t102 S.n14147 0.001
R54651 S.n14147 S.n14144 0.001
R54652 S.t9 S.n22531 0.001
R54653 S.t9 S.n22534 0.001
R54654 S.t88 S.n22121 0.001
R54655 S.t88 S.n22118 0.001
R54656 S.n22118 S.n22115 0.001
R54657 S.t100 S.n21508 0.001
R54658 S.t100 S.n21511 0.001
R54659 S.t105 S.n21840 0.001
R54660 S.t105 S.n21843 0.001
R54661 S.t64 S.n20685 0.001
R54662 S.t64 S.n20688 0.001
R54663 S.t7 S.n21030 0.001
R54664 S.t7 S.n21033 0.001
R54665 S.t209 S.n20074 0.001
R54666 S.t209 S.n20077 0.001
R54667 S.t262 S.n19629 0.001
R54668 S.t262 S.n19626 0.001
R54669 S.n19626 S.n19623 0.001
R54670 S.t150 S.n19220 0.001
R54671 S.t150 S.n19223 0.001
R54672 S.t21 S.n18757 0.001
R54673 S.t21 S.n18754 0.001
R54674 S.n18754 S.n18751 0.001
R54675 S.t79 S.n18354 0.001
R54676 S.t79 S.n18357 0.001
R54677 S.t77 S.n17874 0.001
R54678 S.t77 S.n17871 0.001
R54679 S.n17871 S.n17868 0.001
R54680 S.t218 S.n17465 0.001
R54681 S.t218 S.n17468 0.001
R54682 S.t169 S.n16965 0.001
R54683 S.t169 S.n16962 0.001
R54684 S.n16962 S.n16959 0.001
R54685 S.t167 S.n16563 0.001
R54686 S.t167 S.n16566 0.001
R54687 S.t187 S.n16047 0.001
R54688 S.t187 S.n16044 0.001
R54689 S.n16044 S.n16041 0.001
R54690 S.t60 S.n15639 0.001
R54691 S.t60 S.n15642 0.001
R54692 S.t29 S.n15103 0.001
R54693 S.t29 S.n15100 0.001
R54694 S.n15100 S.n15097 0.001
R54695 S.t0 S.n14702 0.001
R54696 S.t0 S.n14705 0.001
R54697 S.n14115 S.n14110 0.001
R54698 S.n13146 S.t443 0.001
R54699 S.t357 S.n12755 0.001
R54700 S.t357 S.n12758 0.001
R54701 S.t538 S.n13186 0.001
R54702 S.t538 S.n13183 0.001
R54703 S.n13183 S.n13180 0.001
R54704 S.t9 S.n22515 0.001
R54705 S.t9 S.n22518 0.001
R54706 S.t88 S.n22136 0.001
R54707 S.t88 S.n22133 0.001
R54708 S.n22133 S.n22130 0.001
R54709 S.t100 S.n21492 0.001
R54710 S.t100 S.n21495 0.001
R54711 S.t105 S.n21825 0.001
R54712 S.t105 S.n21828 0.001
R54713 S.t64 S.n20669 0.001
R54714 S.t64 S.n20672 0.001
R54715 S.t7 S.n21015 0.001
R54716 S.t7 S.n21018 0.001
R54717 S.t209 S.n20058 0.001
R54718 S.t209 S.n20061 0.001
R54719 S.t262 S.n19644 0.001
R54720 S.t262 S.n19641 0.001
R54721 S.n19641 S.n19638 0.001
R54722 S.t150 S.n19204 0.001
R54723 S.t150 S.n19207 0.001
R54724 S.t21 S.n18772 0.001
R54725 S.t21 S.n18769 0.001
R54726 S.n18769 S.n18766 0.001
R54727 S.t79 S.n18338 0.001
R54728 S.t79 S.n18341 0.001
R54729 S.t77 S.n17889 0.001
R54730 S.t77 S.n17886 0.001
R54731 S.n17886 S.n17883 0.001
R54732 S.t218 S.n17449 0.001
R54733 S.t218 S.n17452 0.001
R54734 S.t169 S.n16980 0.001
R54735 S.t169 S.n16977 0.001
R54736 S.n16977 S.n16974 0.001
R54737 S.t167 S.n16547 0.001
R54738 S.t167 S.n16550 0.001
R54739 S.t187 S.n16062 0.001
R54740 S.t187 S.n16059 0.001
R54741 S.n16059 S.n16056 0.001
R54742 S.t60 S.n15623 0.001
R54743 S.t60 S.n15626 0.001
R54744 S.t29 S.n15118 0.001
R54745 S.t29 S.n15115 0.001
R54746 S.n15115 S.n15112 0.001
R54747 S.t0 S.n14686 0.001
R54748 S.t0 S.n14689 0.001
R54749 S.t102 S.n14165 0.001
R54750 S.t102 S.n14162 0.001
R54751 S.n14162 S.n14159 0.001
R54752 S.t73 S.n13727 0.001
R54753 S.t73 S.n13730 0.001
R54754 S.n13151 S.n13146 0.001
R54755 S.n12173 S.t67 0.001
R54756 S.t54 S.n11745 0.001
R54757 S.t54 S.n11748 0.001
R54758 S.t443 S.n12213 0.001
R54759 S.t443 S.n12210 0.001
R54760 S.n12210 S.n12207 0.001
R54761 S.t9 S.n22499 0.001
R54762 S.t9 S.n22502 0.001
R54763 S.t88 S.n22151 0.001
R54764 S.t88 S.n22148 0.001
R54765 S.n22148 S.n22145 0.001
R54766 S.t100 S.n21476 0.001
R54767 S.t100 S.n21479 0.001
R54768 S.t105 S.n21810 0.001
R54769 S.t105 S.n21813 0.001
R54770 S.t64 S.n20653 0.001
R54771 S.t64 S.n20656 0.001
R54772 S.t7 S.n21000 0.001
R54773 S.t7 S.n21003 0.001
R54774 S.t209 S.n20042 0.001
R54775 S.t209 S.n20045 0.001
R54776 S.t262 S.n19659 0.001
R54777 S.t262 S.n19656 0.001
R54778 S.n19656 S.n19653 0.001
R54779 S.t150 S.n19188 0.001
R54780 S.t150 S.n19191 0.001
R54781 S.t21 S.n18787 0.001
R54782 S.t21 S.n18784 0.001
R54783 S.n18784 S.n18781 0.001
R54784 S.t79 S.n18322 0.001
R54785 S.t79 S.n18325 0.001
R54786 S.t77 S.n17904 0.001
R54787 S.t77 S.n17901 0.001
R54788 S.n17901 S.n17898 0.001
R54789 S.t218 S.n17433 0.001
R54790 S.t218 S.n17436 0.001
R54791 S.t169 S.n16995 0.001
R54792 S.t169 S.n16992 0.001
R54793 S.n16992 S.n16989 0.001
R54794 S.t167 S.n16531 0.001
R54795 S.t167 S.n16534 0.001
R54796 S.t187 S.n16077 0.001
R54797 S.t187 S.n16074 0.001
R54798 S.n16074 S.n16071 0.001
R54799 S.t60 S.n15607 0.001
R54800 S.t60 S.n15610 0.001
R54801 S.t29 S.n15133 0.001
R54802 S.t29 S.n15130 0.001
R54803 S.n15130 S.n15127 0.001
R54804 S.t0 S.n14670 0.001
R54805 S.t0 S.n14673 0.001
R54806 S.t102 S.n14180 0.001
R54807 S.t102 S.n14177 0.001
R54808 S.n14177 S.n14174 0.001
R54809 S.t73 S.n13711 0.001
R54810 S.t73 S.n13714 0.001
R54811 S.t538 S.n13201 0.001
R54812 S.t538 S.n13198 0.001
R54813 S.n13198 S.n13195 0.001
R54814 S.t357 S.n12739 0.001
R54815 S.t357 S.n12742 0.001
R54816 S.n12178 S.n12173 0.001
R54817 S.n11174 S.t172 0.001
R54818 S.t31 S.n10722 0.001
R54819 S.t31 S.n10725 0.001
R54820 S.t67 S.n11214 0.001
R54821 S.t67 S.n11211 0.001
R54822 S.n11211 S.n11208 0.001
R54823 S.t9 S.n22483 0.001
R54824 S.t9 S.n22486 0.001
R54825 S.t88 S.n22166 0.001
R54826 S.t88 S.n22163 0.001
R54827 S.n22163 S.n22160 0.001
R54828 S.t100 S.n21460 0.001
R54829 S.t100 S.n21463 0.001
R54830 S.t105 S.n21795 0.001
R54831 S.t105 S.n21798 0.001
R54832 S.t64 S.n20637 0.001
R54833 S.t64 S.n20640 0.001
R54834 S.t7 S.n20985 0.001
R54835 S.t7 S.n20988 0.001
R54836 S.t209 S.n20026 0.001
R54837 S.t209 S.n20029 0.001
R54838 S.t262 S.n19674 0.001
R54839 S.t262 S.n19671 0.001
R54840 S.n19671 S.n19668 0.001
R54841 S.t150 S.n19172 0.001
R54842 S.t150 S.n19175 0.001
R54843 S.t21 S.n18802 0.001
R54844 S.t21 S.n18799 0.001
R54845 S.n18799 S.n18796 0.001
R54846 S.t79 S.n18306 0.001
R54847 S.t79 S.n18309 0.001
R54848 S.t77 S.n17919 0.001
R54849 S.t77 S.n17916 0.001
R54850 S.n17916 S.n17913 0.001
R54851 S.t218 S.n17417 0.001
R54852 S.t218 S.n17420 0.001
R54853 S.t169 S.n17010 0.001
R54854 S.t169 S.n17007 0.001
R54855 S.n17007 S.n17004 0.001
R54856 S.t167 S.n16515 0.001
R54857 S.t167 S.n16518 0.001
R54858 S.t187 S.n16092 0.001
R54859 S.t187 S.n16089 0.001
R54860 S.n16089 S.n16086 0.001
R54861 S.t60 S.n15591 0.001
R54862 S.t60 S.n15594 0.001
R54863 S.t29 S.n15148 0.001
R54864 S.t29 S.n15145 0.001
R54865 S.n15145 S.n15142 0.001
R54866 S.t0 S.n14654 0.001
R54867 S.t0 S.n14657 0.001
R54868 S.t102 S.n14195 0.001
R54869 S.t102 S.n14192 0.001
R54870 S.n14192 S.n14189 0.001
R54871 S.t73 S.n13695 0.001
R54872 S.t73 S.n13698 0.001
R54873 S.t538 S.n13216 0.001
R54874 S.t538 S.n13213 0.001
R54875 S.n13213 S.n13210 0.001
R54876 S.t357 S.n12723 0.001
R54877 S.t357 S.n12726 0.001
R54878 S.t443 S.n12228 0.001
R54879 S.t443 S.n12225 0.001
R54880 S.n12225 S.n12222 0.001
R54881 S.t54 S.n11729 0.001
R54882 S.t54 S.n11732 0.001
R54883 S.n11179 S.n11174 0.001
R54884 S.n10166 S.t160 0.001
R54885 S.t366 S.n9677 0.001
R54886 S.t366 S.n9680 0.001
R54887 S.t172 S.n10206 0.001
R54888 S.t172 S.n10203 0.001
R54889 S.n10203 S.n10200 0.001
R54890 S.t9 S.n22467 0.001
R54891 S.t9 S.n22470 0.001
R54892 S.t88 S.n22181 0.001
R54893 S.t88 S.n22178 0.001
R54894 S.n22178 S.n22175 0.001
R54895 S.t100 S.n21444 0.001
R54896 S.t100 S.n21447 0.001
R54897 S.t105 S.n21780 0.001
R54898 S.t105 S.n21783 0.001
R54899 S.t64 S.n20621 0.001
R54900 S.t64 S.n20624 0.001
R54901 S.t7 S.n20970 0.001
R54902 S.t7 S.n20973 0.001
R54903 S.t209 S.n20010 0.001
R54904 S.t209 S.n20013 0.001
R54905 S.t262 S.n19689 0.001
R54906 S.t262 S.n19686 0.001
R54907 S.n19686 S.n19683 0.001
R54908 S.t150 S.n19156 0.001
R54909 S.t150 S.n19159 0.001
R54910 S.t21 S.n18817 0.001
R54911 S.t21 S.n18814 0.001
R54912 S.n18814 S.n18811 0.001
R54913 S.t79 S.n18290 0.001
R54914 S.t79 S.n18293 0.001
R54915 S.t77 S.n17934 0.001
R54916 S.t77 S.n17931 0.001
R54917 S.n17931 S.n17928 0.001
R54918 S.t218 S.n17401 0.001
R54919 S.t218 S.n17404 0.001
R54920 S.t169 S.n17025 0.001
R54921 S.t169 S.n17022 0.001
R54922 S.n17022 S.n17019 0.001
R54923 S.t167 S.n16499 0.001
R54924 S.t167 S.n16502 0.001
R54925 S.t187 S.n16107 0.001
R54926 S.t187 S.n16104 0.001
R54927 S.n16104 S.n16101 0.001
R54928 S.t60 S.n15575 0.001
R54929 S.t60 S.n15578 0.001
R54930 S.t29 S.n15163 0.001
R54931 S.t29 S.n15160 0.001
R54932 S.n15160 S.n15157 0.001
R54933 S.t0 S.n14638 0.001
R54934 S.t0 S.n14641 0.001
R54935 S.t102 S.n14210 0.001
R54936 S.t102 S.n14207 0.001
R54937 S.n14207 S.n14204 0.001
R54938 S.t73 S.n13679 0.001
R54939 S.t73 S.n13682 0.001
R54940 S.t538 S.n13231 0.001
R54941 S.t538 S.n13228 0.001
R54942 S.n13228 S.n13225 0.001
R54943 S.t357 S.n12707 0.001
R54944 S.t357 S.n12710 0.001
R54945 S.t443 S.n12243 0.001
R54946 S.t443 S.n12240 0.001
R54947 S.n12240 S.n12237 0.001
R54948 S.t54 S.n11713 0.001
R54949 S.t54 S.n11716 0.001
R54950 S.t67 S.n11229 0.001
R54951 S.t67 S.n11226 0.001
R54952 S.n11226 S.n11223 0.001
R54953 S.t31 S.n10706 0.001
R54954 S.t31 S.n10709 0.001
R54955 S.n10171 S.n10166 0.001
R54956 S.n9132 S.t141 0.001
R54957 S.t19 S.n8619 0.001
R54958 S.t19 S.n8622 0.001
R54959 S.t160 S.n9172 0.001
R54960 S.t160 S.n9169 0.001
R54961 S.n9169 S.n9166 0.001
R54962 S.t9 S.n22451 0.001
R54963 S.t9 S.n22454 0.001
R54964 S.t88 S.n22196 0.001
R54965 S.t88 S.n22193 0.001
R54966 S.n22193 S.n22190 0.001
R54967 S.t100 S.n21428 0.001
R54968 S.t100 S.n21431 0.001
R54969 S.t105 S.n21765 0.001
R54970 S.t105 S.n21768 0.001
R54971 S.t64 S.n20605 0.001
R54972 S.t64 S.n20608 0.001
R54973 S.t7 S.n20955 0.001
R54974 S.t7 S.n20958 0.001
R54975 S.t209 S.n19994 0.001
R54976 S.t209 S.n19997 0.001
R54977 S.t262 S.n19704 0.001
R54978 S.t262 S.n19701 0.001
R54979 S.n19701 S.n19698 0.001
R54980 S.t150 S.n19140 0.001
R54981 S.t150 S.n19143 0.001
R54982 S.t21 S.n18832 0.001
R54983 S.t21 S.n18829 0.001
R54984 S.n18829 S.n18826 0.001
R54985 S.t79 S.n18274 0.001
R54986 S.t79 S.n18277 0.001
R54987 S.t77 S.n17949 0.001
R54988 S.t77 S.n17946 0.001
R54989 S.n17946 S.n17943 0.001
R54990 S.t218 S.n17385 0.001
R54991 S.t218 S.n17388 0.001
R54992 S.t169 S.n17040 0.001
R54993 S.t169 S.n17037 0.001
R54994 S.n17037 S.n17034 0.001
R54995 S.t167 S.n16483 0.001
R54996 S.t167 S.n16486 0.001
R54997 S.t187 S.n16122 0.001
R54998 S.t187 S.n16119 0.001
R54999 S.n16119 S.n16116 0.001
R55000 S.t60 S.n15559 0.001
R55001 S.t60 S.n15562 0.001
R55002 S.t29 S.n15178 0.001
R55003 S.t29 S.n15175 0.001
R55004 S.n15175 S.n15172 0.001
R55005 S.t0 S.n14622 0.001
R55006 S.t0 S.n14625 0.001
R55007 S.t102 S.n14225 0.001
R55008 S.t102 S.n14222 0.001
R55009 S.n14222 S.n14219 0.001
R55010 S.t73 S.n13663 0.001
R55011 S.t73 S.n13666 0.001
R55012 S.t538 S.n13246 0.001
R55013 S.t538 S.n13243 0.001
R55014 S.n13243 S.n13240 0.001
R55015 S.t357 S.n12691 0.001
R55016 S.t357 S.n12694 0.001
R55017 S.t443 S.n12258 0.001
R55018 S.t443 S.n12255 0.001
R55019 S.n12255 S.n12252 0.001
R55020 S.t54 S.n11697 0.001
R55021 S.t54 S.n11700 0.001
R55022 S.t67 S.n11244 0.001
R55023 S.t67 S.n11241 0.001
R55024 S.n11241 S.n11238 0.001
R55025 S.t31 S.n10690 0.001
R55026 S.t31 S.n10693 0.001
R55027 S.t172 S.n10221 0.001
R55028 S.t172 S.n10218 0.001
R55029 S.n10218 S.n10215 0.001
R55030 S.t366 S.n9661 0.001
R55031 S.t366 S.n9664 0.001
R55032 S.n9137 S.n9132 0.001
R55033 S.n8089 S.t406 0.001
R55034 S.t47 S.n7539 0.001
R55035 S.t47 S.n7542 0.001
R55036 S.t141 S.n8129 0.001
R55037 S.t141 S.n8126 0.001
R55038 S.n8126 S.n8123 0.001
R55039 S.t9 S.n22435 0.001
R55040 S.t9 S.n22438 0.001
R55041 S.t88 S.n22211 0.001
R55042 S.t88 S.n22208 0.001
R55043 S.n22208 S.n22205 0.001
R55044 S.t100 S.n21412 0.001
R55045 S.t100 S.n21415 0.001
R55046 S.t105 S.n21750 0.001
R55047 S.t105 S.n21753 0.001
R55048 S.t64 S.n20589 0.001
R55049 S.t64 S.n20592 0.001
R55050 S.t7 S.n20940 0.001
R55051 S.t7 S.n20943 0.001
R55052 S.t209 S.n19978 0.001
R55053 S.t209 S.n19981 0.001
R55054 S.t262 S.n19719 0.001
R55055 S.t262 S.n19716 0.001
R55056 S.n19716 S.n19713 0.001
R55057 S.t150 S.n19124 0.001
R55058 S.t150 S.n19127 0.001
R55059 S.t21 S.n18847 0.001
R55060 S.t21 S.n18844 0.001
R55061 S.n18844 S.n18841 0.001
R55062 S.t79 S.n18258 0.001
R55063 S.t79 S.n18261 0.001
R55064 S.t77 S.n17964 0.001
R55065 S.t77 S.n17961 0.001
R55066 S.n17961 S.n17958 0.001
R55067 S.t218 S.n17369 0.001
R55068 S.t218 S.n17372 0.001
R55069 S.t169 S.n17055 0.001
R55070 S.t169 S.n17052 0.001
R55071 S.n17052 S.n17049 0.001
R55072 S.t167 S.n16467 0.001
R55073 S.t167 S.n16470 0.001
R55074 S.t187 S.n16137 0.001
R55075 S.t187 S.n16134 0.001
R55076 S.n16134 S.n16131 0.001
R55077 S.t60 S.n15543 0.001
R55078 S.t60 S.n15546 0.001
R55079 S.t29 S.n15193 0.001
R55080 S.t29 S.n15190 0.001
R55081 S.n15190 S.n15187 0.001
R55082 S.t0 S.n14606 0.001
R55083 S.t0 S.n14609 0.001
R55084 S.t102 S.n14240 0.001
R55085 S.t102 S.n14237 0.001
R55086 S.n14237 S.n14234 0.001
R55087 S.t73 S.n13647 0.001
R55088 S.t73 S.n13650 0.001
R55089 S.t538 S.n13261 0.001
R55090 S.t538 S.n13258 0.001
R55091 S.n13258 S.n13255 0.001
R55092 S.t357 S.n12675 0.001
R55093 S.t357 S.n12678 0.001
R55094 S.t443 S.n12273 0.001
R55095 S.t443 S.n12270 0.001
R55096 S.n12270 S.n12267 0.001
R55097 S.t54 S.n11681 0.001
R55098 S.t54 S.n11684 0.001
R55099 S.t67 S.n11259 0.001
R55100 S.t67 S.n11256 0.001
R55101 S.n11256 S.n11253 0.001
R55102 S.t31 S.n10674 0.001
R55103 S.t31 S.n10677 0.001
R55104 S.t172 S.n10236 0.001
R55105 S.t172 S.n10233 0.001
R55106 S.n10233 S.n10230 0.001
R55107 S.t366 S.n9645 0.001
R55108 S.t366 S.n9648 0.001
R55109 S.t160 S.n9187 0.001
R55110 S.t160 S.n9184 0.001
R55111 S.n9184 S.n9181 0.001
R55112 S.t19 S.n8603 0.001
R55113 S.t19 S.n8606 0.001
R55114 S.n8094 S.n8089 0.001
R55115 S.n7020 S.t130 0.001
R55116 S.t83 S.n6446 0.001
R55117 S.t83 S.n6449 0.001
R55118 S.t406 S.n7060 0.001
R55119 S.t406 S.n7057 0.001
R55120 S.n7057 S.n7054 0.001
R55121 S.t9 S.n22419 0.001
R55122 S.t9 S.n22422 0.001
R55123 S.t88 S.n22226 0.001
R55124 S.t88 S.n22223 0.001
R55125 S.n22223 S.n22220 0.001
R55126 S.t100 S.n21396 0.001
R55127 S.t100 S.n21399 0.001
R55128 S.t105 S.n21735 0.001
R55129 S.t105 S.n21738 0.001
R55130 S.t64 S.n20573 0.001
R55131 S.t64 S.n20576 0.001
R55132 S.t7 S.n20925 0.001
R55133 S.t7 S.n20928 0.001
R55134 S.t209 S.n19962 0.001
R55135 S.t209 S.n19965 0.001
R55136 S.t262 S.n19734 0.001
R55137 S.t262 S.n19731 0.001
R55138 S.n19731 S.n19728 0.001
R55139 S.t150 S.n19108 0.001
R55140 S.t150 S.n19111 0.001
R55141 S.t21 S.n18862 0.001
R55142 S.t21 S.n18859 0.001
R55143 S.n18859 S.n18856 0.001
R55144 S.t79 S.n18242 0.001
R55145 S.t79 S.n18245 0.001
R55146 S.t77 S.n17979 0.001
R55147 S.t77 S.n17976 0.001
R55148 S.n17976 S.n17973 0.001
R55149 S.t218 S.n17353 0.001
R55150 S.t218 S.n17356 0.001
R55151 S.t169 S.n17070 0.001
R55152 S.t169 S.n17067 0.001
R55153 S.n17067 S.n17064 0.001
R55154 S.t167 S.n16451 0.001
R55155 S.t167 S.n16454 0.001
R55156 S.t187 S.n16152 0.001
R55157 S.t187 S.n16149 0.001
R55158 S.n16149 S.n16146 0.001
R55159 S.t60 S.n15527 0.001
R55160 S.t60 S.n15530 0.001
R55161 S.t29 S.n15208 0.001
R55162 S.t29 S.n15205 0.001
R55163 S.n15205 S.n15202 0.001
R55164 S.t0 S.n14590 0.001
R55165 S.t0 S.n14593 0.001
R55166 S.t102 S.n14255 0.001
R55167 S.t102 S.n14252 0.001
R55168 S.n14252 S.n14249 0.001
R55169 S.t73 S.n13631 0.001
R55170 S.t73 S.n13634 0.001
R55171 S.t538 S.n13276 0.001
R55172 S.t538 S.n13273 0.001
R55173 S.n13273 S.n13270 0.001
R55174 S.t357 S.n12659 0.001
R55175 S.t357 S.n12662 0.001
R55176 S.t443 S.n12288 0.001
R55177 S.t443 S.n12285 0.001
R55178 S.n12285 S.n12282 0.001
R55179 S.t54 S.n11665 0.001
R55180 S.t54 S.n11668 0.001
R55181 S.t67 S.n11274 0.001
R55182 S.t67 S.n11271 0.001
R55183 S.n11271 S.n11268 0.001
R55184 S.t31 S.n10658 0.001
R55185 S.t31 S.n10661 0.001
R55186 S.t172 S.n10251 0.001
R55187 S.t172 S.n10248 0.001
R55188 S.n10248 S.n10245 0.001
R55189 S.t366 S.n9629 0.001
R55190 S.t366 S.n9632 0.001
R55191 S.t160 S.n9202 0.001
R55192 S.t160 S.n9199 0.001
R55193 S.n9199 S.n9196 0.001
R55194 S.t19 S.n8587 0.001
R55195 S.t19 S.n8590 0.001
R55196 S.t141 S.n8144 0.001
R55197 S.t141 S.n8141 0.001
R55198 S.n8141 S.n8138 0.001
R55199 S.t47 S.n7523 0.001
R55200 S.t47 S.n7526 0.001
R55201 S.n7025 S.n7020 0.001
R55202 S.n5942 S.t288 0.001
R55203 S.t214 S.n5330 0.001
R55204 S.t214 S.n5333 0.001
R55205 S.t130 S.n5982 0.001
R55206 S.t130 S.n5979 0.001
R55207 S.n5979 S.n5976 0.001
R55208 S.t9 S.n22403 0.001
R55209 S.t9 S.n22406 0.001
R55210 S.t88 S.n22241 0.001
R55211 S.t88 S.n22238 0.001
R55212 S.n22238 S.n22235 0.001
R55213 S.t100 S.n21380 0.001
R55214 S.t100 S.n21383 0.001
R55215 S.t105 S.n21720 0.001
R55216 S.t105 S.n21723 0.001
R55217 S.t64 S.n20557 0.001
R55218 S.t64 S.n20560 0.001
R55219 S.t7 S.n20910 0.001
R55220 S.t7 S.n20913 0.001
R55221 S.t209 S.n19946 0.001
R55222 S.t209 S.n19949 0.001
R55223 S.t262 S.n19749 0.001
R55224 S.t262 S.n19746 0.001
R55225 S.n19746 S.n19743 0.001
R55226 S.t150 S.n19092 0.001
R55227 S.t150 S.n19095 0.001
R55228 S.t21 S.n18877 0.001
R55229 S.t21 S.n18874 0.001
R55230 S.n18874 S.n18871 0.001
R55231 S.t79 S.n18226 0.001
R55232 S.t79 S.n18229 0.001
R55233 S.t77 S.n17994 0.001
R55234 S.t77 S.n17991 0.001
R55235 S.n17991 S.n17988 0.001
R55236 S.t218 S.n17337 0.001
R55237 S.t218 S.n17340 0.001
R55238 S.t169 S.n17085 0.001
R55239 S.t169 S.n17082 0.001
R55240 S.n17082 S.n17079 0.001
R55241 S.t167 S.n16435 0.001
R55242 S.t167 S.n16438 0.001
R55243 S.t187 S.n16167 0.001
R55244 S.t187 S.n16164 0.001
R55245 S.n16164 S.n16161 0.001
R55246 S.t60 S.n15511 0.001
R55247 S.t60 S.n15514 0.001
R55248 S.t29 S.n15223 0.001
R55249 S.t29 S.n15220 0.001
R55250 S.n15220 S.n15217 0.001
R55251 S.t0 S.n14574 0.001
R55252 S.t0 S.n14577 0.001
R55253 S.t102 S.n14270 0.001
R55254 S.t102 S.n14267 0.001
R55255 S.n14267 S.n14264 0.001
R55256 S.t73 S.n13615 0.001
R55257 S.t73 S.n13618 0.001
R55258 S.t538 S.n13291 0.001
R55259 S.t538 S.n13288 0.001
R55260 S.n13288 S.n13285 0.001
R55261 S.t357 S.n12643 0.001
R55262 S.t357 S.n12646 0.001
R55263 S.t443 S.n12303 0.001
R55264 S.t443 S.n12300 0.001
R55265 S.n12300 S.n12297 0.001
R55266 S.t54 S.n11649 0.001
R55267 S.t54 S.n11652 0.001
R55268 S.t67 S.n11289 0.001
R55269 S.t67 S.n11286 0.001
R55270 S.n11286 S.n11283 0.001
R55271 S.t31 S.n10642 0.001
R55272 S.t31 S.n10645 0.001
R55273 S.t172 S.n10266 0.001
R55274 S.t172 S.n10263 0.001
R55275 S.n10263 S.n10260 0.001
R55276 S.t366 S.n9613 0.001
R55277 S.t366 S.n9616 0.001
R55278 S.t160 S.n9217 0.001
R55279 S.t160 S.n9214 0.001
R55280 S.n9214 S.n9211 0.001
R55281 S.t19 S.n8571 0.001
R55282 S.t19 S.n8574 0.001
R55283 S.t141 S.n8159 0.001
R55284 S.t141 S.n8156 0.001
R55285 S.n8156 S.n8153 0.001
R55286 S.t47 S.n7507 0.001
R55287 S.t47 S.n7510 0.001
R55288 S.t406 S.n7075 0.001
R55289 S.t406 S.n7072 0.001
R55290 S.n7072 S.n7069 0.001
R55291 S.t83 S.n6430 0.001
R55292 S.t83 S.n6433 0.001
R55293 S.n5947 S.n5942 0.001
R55294 S.n4836 S.t134 0.001
R55295 S.t176 S.n4201 0.001
R55296 S.t176 S.n4204 0.001
R55297 S.t288 S.n4877 0.001
R55298 S.t288 S.n4874 0.001
R55299 S.n4874 S.n4871 0.001
R55300 S.t9 S.n22387 0.001
R55301 S.t9 S.n22390 0.001
R55302 S.t88 S.n22256 0.001
R55303 S.t88 S.n22253 0.001
R55304 S.n22253 S.n22250 0.001
R55305 S.t100 S.n21364 0.001
R55306 S.t100 S.n21367 0.001
R55307 S.t105 S.n21705 0.001
R55308 S.t105 S.n21708 0.001
R55309 S.t64 S.n20541 0.001
R55310 S.t64 S.n20544 0.001
R55311 S.t7 S.n20895 0.001
R55312 S.t7 S.n20898 0.001
R55313 S.t209 S.n19930 0.001
R55314 S.t209 S.n19933 0.001
R55315 S.t262 S.n19764 0.001
R55316 S.t262 S.n19761 0.001
R55317 S.n19761 S.n19758 0.001
R55318 S.t150 S.n19076 0.001
R55319 S.t150 S.n19079 0.001
R55320 S.t21 S.n18892 0.001
R55321 S.t21 S.n18889 0.001
R55322 S.n18889 S.n18886 0.001
R55323 S.t79 S.n18210 0.001
R55324 S.t79 S.n18213 0.001
R55325 S.t77 S.n18009 0.001
R55326 S.t77 S.n18006 0.001
R55327 S.n18006 S.n18003 0.001
R55328 S.t218 S.n17321 0.001
R55329 S.t218 S.n17324 0.001
R55330 S.t169 S.n17100 0.001
R55331 S.t169 S.n17097 0.001
R55332 S.n17097 S.n17094 0.001
R55333 S.t167 S.n16419 0.001
R55334 S.t167 S.n16422 0.001
R55335 S.t187 S.n16182 0.001
R55336 S.t187 S.n16179 0.001
R55337 S.n16179 S.n16176 0.001
R55338 S.t60 S.n15495 0.001
R55339 S.t60 S.n15498 0.001
R55340 S.t29 S.n15238 0.001
R55341 S.t29 S.n15235 0.001
R55342 S.n15235 S.n15232 0.001
R55343 S.t0 S.n14558 0.001
R55344 S.t0 S.n14561 0.001
R55345 S.t102 S.n14285 0.001
R55346 S.t102 S.n14282 0.001
R55347 S.n14282 S.n14279 0.001
R55348 S.t73 S.n13599 0.001
R55349 S.t73 S.n13602 0.001
R55350 S.t538 S.n13306 0.001
R55351 S.t538 S.n13303 0.001
R55352 S.n13303 S.n13300 0.001
R55353 S.t357 S.n12627 0.001
R55354 S.t357 S.n12630 0.001
R55355 S.t443 S.n12318 0.001
R55356 S.t443 S.n12315 0.001
R55357 S.n12315 S.n12312 0.001
R55358 S.t54 S.n11633 0.001
R55359 S.t54 S.n11636 0.001
R55360 S.t67 S.n11304 0.001
R55361 S.t67 S.n11301 0.001
R55362 S.n11301 S.n11298 0.001
R55363 S.t31 S.n10626 0.001
R55364 S.t31 S.n10629 0.001
R55365 S.t172 S.n10281 0.001
R55366 S.t172 S.n10278 0.001
R55367 S.n10278 S.n10275 0.001
R55368 S.t366 S.n9597 0.001
R55369 S.t366 S.n9600 0.001
R55370 S.t160 S.n9232 0.001
R55371 S.t160 S.n9220 0.001
R55372 S.t19 S.n8555 0.001
R55373 S.t19 S.n8558 0.001
R55374 S.t141 S.n8174 0.001
R55375 S.t141 S.n8171 0.001
R55376 S.n8171 S.n8168 0.001
R55377 S.t47 S.n7491 0.001
R55378 S.t47 S.n7494 0.001
R55379 S.t406 S.n7090 0.001
R55380 S.t406 S.n7087 0.001
R55381 S.n7087 S.n7084 0.001
R55382 S.t83 S.n6414 0.001
R55383 S.t83 S.n6417 0.001
R55384 S.t130 S.n5997 0.001
R55385 S.t130 S.n5994 0.001
R55386 S.n5994 S.n5991 0.001
R55387 S.t214 S.n5314 0.001
R55388 S.t214 S.n5317 0.001
R55389 S.n4841 S.n4836 0.001
R55390 S.n3723 S.t163 0.001
R55391 S.t14 S.n3060 0.001
R55392 S.t14 S.n3063 0.001
R55393 S.t134 S.n3765 0.001
R55394 S.t134 S.n3762 0.001
R55395 S.n3762 S.n3759 0.001
R55396 S.n22665 S.t9 0.001
R55397 S.n22672 S.n22665 0.001
R55398 S.t88 S.n22681 0.001
R55399 S.t88 S.n22678 0.001
R55400 S.n22678 S.n22675 0.001
R55401 S.n21685 S.n21678 0.001
R55402 S.t105 S.n21690 0.001
R55403 S.t105 S.n21693 0.001
R55404 S.t64 S.n20525 0.001
R55405 S.t64 S.n20528 0.001
R55406 S.t7 S.n20880 0.001
R55407 S.t7 S.n20883 0.001
R55408 S.t209 S.n19914 0.001
R55409 S.t209 S.n19917 0.001
R55410 S.t262 S.n19780 0.001
R55411 S.t262 S.n19777 0.001
R55412 S.n19777 S.n19774 0.001
R55413 S.t150 S.n19060 0.001
R55414 S.t150 S.n19063 0.001
R55415 S.t21 S.n18908 0.001
R55416 S.t21 S.n18905 0.001
R55417 S.n18905 S.n18902 0.001
R55418 S.t79 S.n18194 0.001
R55419 S.t79 S.n18197 0.001
R55420 S.t77 S.n18025 0.001
R55421 S.t77 S.n18022 0.001
R55422 S.n18022 S.n18019 0.001
R55423 S.t218 S.n17305 0.001
R55424 S.t218 S.n17308 0.001
R55425 S.t169 S.n17116 0.001
R55426 S.t169 S.n17113 0.001
R55427 S.n17113 S.n17110 0.001
R55428 S.t167 S.n16403 0.001
R55429 S.t167 S.n16406 0.001
R55430 S.t187 S.n16198 0.001
R55431 S.t187 S.n16195 0.001
R55432 S.n16195 S.n16192 0.001
R55433 S.t60 S.n15479 0.001
R55434 S.t60 S.n15482 0.001
R55435 S.t29 S.n15254 0.001
R55436 S.t29 S.n15251 0.001
R55437 S.n15251 S.n15248 0.001
R55438 S.t0 S.n14542 0.001
R55439 S.t0 S.n14545 0.001
R55440 S.t102 S.n14301 0.001
R55441 S.t102 S.n14298 0.001
R55442 S.n14298 S.n14295 0.001
R55443 S.t73 S.n13583 0.001
R55444 S.t73 S.n13586 0.001
R55445 S.t538 S.n13322 0.001
R55446 S.t538 S.n13319 0.001
R55447 S.n13319 S.n13316 0.001
R55448 S.t357 S.n12611 0.001
R55449 S.t357 S.n12614 0.001
R55450 S.t443 S.n12334 0.001
R55451 S.t443 S.n12331 0.001
R55452 S.n12331 S.n12328 0.001
R55453 S.t54 S.n11617 0.001
R55454 S.t54 S.n11620 0.001
R55455 S.t67 S.n11320 0.001
R55456 S.t67 S.n11317 0.001
R55457 S.n11317 S.n11314 0.001
R55458 S.t31 S.n10610 0.001
R55459 S.t31 S.n10613 0.001
R55460 S.t172 S.n10297 0.001
R55461 S.t172 S.n10294 0.001
R55462 S.n10294 S.n10291 0.001
R55463 S.t366 S.n9581 0.001
R55464 S.t366 S.n9584 0.001
R55465 S.t160 S.n9248 0.001
R55466 S.t160 S.n9245 0.001
R55467 S.n9245 S.n9242 0.001
R55468 S.t19 S.n8539 0.001
R55469 S.t19 S.n8542 0.001
R55470 S.t141 S.n8190 0.001
R55471 S.t141 S.n8187 0.001
R55472 S.n8187 S.n8184 0.001
R55473 S.t47 S.n7475 0.001
R55474 S.t47 S.n7478 0.001
R55475 S.t406 S.n7106 0.001
R55476 S.t406 S.n7103 0.001
R55477 S.n7103 S.n7100 0.001
R55478 S.t83 S.n6398 0.001
R55479 S.t83 S.n6401 0.001
R55480 S.t130 S.n6013 0.001
R55481 S.t130 S.n6010 0.001
R55482 S.n6010 S.n6007 0.001
R55483 S.t214 S.n5298 0.001
R55484 S.t214 S.n5301 0.001
R55485 S.t288 S.n4893 0.001
R55486 S.t288 S.n4890 0.001
R55487 S.n4890 S.n4887 0.001
R55488 S.t176 S.n4185 0.001
R55489 S.t176 S.n4188 0.001
R55490 S.n3728 S.n3723 0.001
R55491 S.n2592 S.t270 0.001
R55492 S.n1891 S.t75 0.001
R55493 S.n1899 S.n1894 0.001
R55494 S.t163 S.n2634 0.001
R55495 S.t163 S.n2631 0.001
R55496 S.n2631 S.n2628 0.001
R55497 S.t9 S.n22371 0.001
R55498 S.t9 S.n22374 0.001
R55499 S.t88 S.n22700 0.001
R55500 S.t88 S.n22697 0.001
R55501 S.n22697 S.n22694 0.001
R55502 S.n21647 S.t100 0.001
R55503 S.n21654 S.n21647 0.001
R55504 S.t105 S.n21659 0.001
R55505 S.t105 S.n21662 0.001
R55506 S.t64 S.n20510 0.001
R55507 S.t64 S.n20513 0.001
R55508 S.t7 S.n20864 0.001
R55509 S.t7 S.n20867 0.001
R55510 S.t209 S.n19899 0.001
R55511 S.t209 S.n19902 0.001
R55512 S.t262 S.n19796 0.001
R55513 S.t262 S.n19793 0.001
R55514 S.n19793 S.n19790 0.001
R55515 S.t150 S.n19045 0.001
R55516 S.t150 S.n19048 0.001
R55517 S.t21 S.n18924 0.001
R55518 S.t21 S.n18921 0.001
R55519 S.n18921 S.n18918 0.001
R55520 S.t79 S.n18179 0.001
R55521 S.t79 S.n18182 0.001
R55522 S.t77 S.n18041 0.001
R55523 S.t77 S.n18038 0.001
R55524 S.n18038 S.n18035 0.001
R55525 S.t218 S.n17290 0.001
R55526 S.t218 S.n17293 0.001
R55527 S.t169 S.n17132 0.001
R55528 S.t169 S.n17129 0.001
R55529 S.n17129 S.n17126 0.001
R55530 S.t167 S.n16388 0.001
R55531 S.t167 S.n16391 0.001
R55532 S.t187 S.n16214 0.001
R55533 S.t187 S.n16211 0.001
R55534 S.n16211 S.n16208 0.001
R55535 S.t60 S.n15464 0.001
R55536 S.t60 S.n15467 0.001
R55537 S.t29 S.n15270 0.001
R55538 S.t29 S.n15267 0.001
R55539 S.n15267 S.n15264 0.001
R55540 S.t0 S.n14527 0.001
R55541 S.t0 S.n14530 0.001
R55542 S.t102 S.n14317 0.001
R55543 S.t102 S.n14314 0.001
R55544 S.n14314 S.n14311 0.001
R55545 S.t73 S.n13568 0.001
R55546 S.t73 S.n13571 0.001
R55547 S.t538 S.n13338 0.001
R55548 S.t538 S.n13335 0.001
R55549 S.n13335 S.n13332 0.001
R55550 S.t357 S.n12596 0.001
R55551 S.t357 S.n12599 0.001
R55552 S.t443 S.n12350 0.001
R55553 S.t443 S.n12347 0.001
R55554 S.n12347 S.n12344 0.001
R55555 S.t54 S.n11602 0.001
R55556 S.t54 S.n11605 0.001
R55557 S.t67 S.n11336 0.001
R55558 S.t67 S.n11333 0.001
R55559 S.n11333 S.n11330 0.001
R55560 S.t31 S.n10595 0.001
R55561 S.t31 S.n10598 0.001
R55562 S.t172 S.n10313 0.001
R55563 S.t172 S.n10310 0.001
R55564 S.n10310 S.n10307 0.001
R55565 S.t366 S.n9566 0.001
R55566 S.t366 S.n9569 0.001
R55567 S.t160 S.n9264 0.001
R55568 S.t160 S.n9261 0.001
R55569 S.n9261 S.n9258 0.001
R55570 S.t19 S.n8524 0.001
R55571 S.t19 S.n8527 0.001
R55572 S.t141 S.n8206 0.001
R55573 S.t141 S.n8203 0.001
R55574 S.n8203 S.n8200 0.001
R55575 S.t47 S.n7460 0.001
R55576 S.t47 S.n7463 0.001
R55577 S.t406 S.n7122 0.001
R55578 S.t406 S.n7119 0.001
R55579 S.n7119 S.n7116 0.001
R55580 S.t83 S.n6383 0.001
R55581 S.t83 S.n6386 0.001
R55582 S.t130 S.n6029 0.001
R55583 S.t130 S.n6026 0.001
R55584 S.n6026 S.n6023 0.001
R55585 S.t214 S.n5283 0.001
R55586 S.t214 S.n5286 0.001
R55587 S.t288 S.n4909 0.001
R55588 S.t288 S.n4906 0.001
R55589 S.n4906 S.n4903 0.001
R55590 S.t176 S.n4170 0.001
R55591 S.t176 S.n4173 0.001
R55592 S.t134 S.n3781 0.001
R55593 S.t134 S.n3778 0.001
R55594 S.n3778 S.n3775 0.001
R55595 S.t14 S.n3044 0.001
R55596 S.t14 S.n3047 0.001
R55597 S.n2597 S.n2592 0.001
R55598 S.n1432 S.n1422 0.001
R55599 S.t109 S.n920 0.001
R55600 S.t109 S.n917 0.001
R55601 S.n917 S.n914 0.001
R55602 S.t270 S.n1988 0.001
R55603 S.t270 S.n1991 0.001
R55604 S.t88 S.n22747 0.001
R55605 S.t88 S.n22744 0.001
R55606 S.n22744 S.n22741 0.001
R55607 S.t100 S.n21320 0.001
R55608 S.t100 S.n21317 0.001
R55609 S.n21317 S.n21314 0.001
R55610 S.t105 S.n21223 0.001
R55611 S.t105 S.n21220 0.001
R55612 S.n21220 S.n21217 0.001
R55613 S.t64 S.n20497 0.001
R55614 S.t64 S.n20494 0.001
R55615 S.n20494 S.n20491 0.001
R55616 S.t7 S.n20404 0.001
R55617 S.t7 S.n20401 0.001
R55618 S.n20401 S.n20398 0.001
R55619 S.t209 S.n19886 0.001
R55620 S.t209 S.n19883 0.001
R55621 S.n19883 S.n19880 0.001
R55622 S.t262 S.n20274 0.001
R55623 S.t262 S.n20277 0.001
R55624 S.t150 S.n19032 0.001
R55625 S.t150 S.n19029 0.001
R55626 S.n19029 S.n19026 0.001
R55627 S.t21 S.n19406 0.001
R55628 S.t21 S.n19409 0.001
R55629 S.t79 S.n18166 0.001
R55630 S.t79 S.n18163 0.001
R55631 S.n18163 S.n18160 0.001
R55632 S.t77 S.n18519 0.001
R55633 S.t77 S.n18522 0.001
R55634 S.t218 S.n17277 0.001
R55635 S.t218 S.n17274 0.001
R55636 S.n17274 S.n17271 0.001
R55637 S.t169 S.n17619 0.001
R55638 S.t169 S.n17622 0.001
R55639 S.t167 S.n16375 0.001
R55640 S.t167 S.n16372 0.001
R55641 S.n16372 S.n16369 0.001
R55642 S.t187 S.n16696 0.001
R55643 S.t187 S.n16699 0.001
R55644 S.t60 S.n15451 0.001
R55645 S.t60 S.n15448 0.001
R55646 S.n15448 S.n15445 0.001
R55647 S.t29 S.n15761 0.001
R55648 S.t29 S.n15764 0.001
R55649 S.t0 S.n14514 0.001
R55650 S.t0 S.n14511 0.001
R55651 S.n14511 S.n14508 0.001
R55652 S.t102 S.n14803 0.001
R55653 S.t102 S.n14806 0.001
R55654 S.t73 S.n13555 0.001
R55655 S.t73 S.n13552 0.001
R55656 S.n13552 S.n13549 0.001
R55657 S.t538 S.n13833 0.001
R55658 S.t538 S.n13836 0.001
R55659 S.t357 S.n12583 0.001
R55660 S.t357 S.n12580 0.001
R55661 S.n12580 S.n12577 0.001
R55662 S.t443 S.n12840 0.001
R55663 S.t443 S.n12843 0.001
R55664 S.t54 S.n11589 0.001
R55665 S.t54 S.n11586 0.001
R55666 S.n11586 S.n11583 0.001
R55667 S.t67 S.n11835 0.001
R55668 S.t67 S.n11838 0.001
R55669 S.t31 S.n10582 0.001
R55670 S.t31 S.n10579 0.001
R55671 S.n10579 S.n10576 0.001
R55672 S.t172 S.n10807 0.001
R55673 S.t172 S.n10810 0.001
R55674 S.t366 S.n9553 0.001
R55675 S.t366 S.n9550 0.001
R55676 S.n9550 S.n9547 0.001
R55677 S.t160 S.n9767 0.001
R55678 S.t160 S.n9770 0.001
R55679 S.t19 S.n8511 0.001
R55680 S.t19 S.n8508 0.001
R55681 S.n8508 S.n8505 0.001
R55682 S.t141 S.n8704 0.001
R55683 S.t141 S.n8707 0.001
R55684 S.t47 S.n7447 0.001
R55685 S.t47 S.n7444 0.001
R55686 S.n7444 S.n7441 0.001
R55687 S.t406 S.n7629 0.001
R55688 S.t406 S.n7632 0.001
R55689 S.t83 S.n6370 0.001
R55690 S.t83 S.n6367 0.001
R55691 S.n6367 S.n6364 0.001
R55692 S.t130 S.n6531 0.001
R55693 S.t130 S.n6534 0.001
R55694 S.t214 S.n5270 0.001
R55695 S.t214 S.n5267 0.001
R55696 S.n5267 S.n5264 0.001
R55697 S.t288 S.n5420 0.001
R55698 S.t288 S.n5423 0.001
R55699 S.t176 S.n4157 0.001
R55700 S.t176 S.n4154 0.001
R55701 S.n4154 S.n4151 0.001
R55702 S.t134 S.n4286 0.001
R55703 S.t134 S.n4289 0.001
R55704 S.t14 S.n3031 0.001
R55705 S.t14 S.n3028 0.001
R55706 S.n3028 S.n3025 0.001
R55707 S.t163 S.n3149 0.001
R55708 S.t163 S.n3152 0.001
R55709 S.t75 S.n1871 0.001
R55710 S.t75 S.n1868 0.001
R55711 S.n1868 S.n1865 0.001
R55712 S.n890 S.n880 0.001
R55713 S.t137 S.n809 0.001
R55714 S.t137 S.n812 0.001
R55715 S.t109 S.n977 0.001
R55716 S.t109 S.n979 0.001
R55717 S.t9 S.n22354 0.001
R55718 S.t9 S.n22357 0.001
R55719 S.t88 S.n22719 0.001
R55720 S.t88 S.n22716 0.001
R55721 S.n22716 S.n22713 0.001
R55722 S.t100 S.n21348 0.001
R55723 S.t100 S.n21351 0.001
R55724 S.t105 S.n21264 0.001
R55725 S.t105 S.n21267 0.001
R55726 S.n20827 S.t64 0.001
R55727 S.n20835 S.n20830 0.001
R55728 S.t7 S.n20848 0.001
R55729 S.t7 S.n20851 0.001
R55730 S.n20192 S.t209 0.001
R55731 S.n20200 S.n20195 0.001
R55732 S.t262 S.n20216 0.001
R55733 S.t262 S.n20213 0.001
R55734 S.n20213 S.n20210 0.001
R55735 S.n19322 S.t150 0.001
R55736 S.n19330 S.n19325 0.001
R55737 S.t21 S.n19346 0.001
R55738 S.t21 S.n19343 0.001
R55739 S.n19343 S.n19340 0.001
R55740 S.n18440 S.t79 0.001
R55741 S.n18448 S.n18443 0.001
R55742 S.t77 S.n18464 0.001
R55743 S.t77 S.n18461 0.001
R55744 S.n18461 S.n18458 0.001
R55745 S.n17535 S.t218 0.001
R55746 S.n17543 S.n17538 0.001
R55747 S.t169 S.n17559 0.001
R55748 S.t169 S.n17556 0.001
R55749 S.n17556 S.n17553 0.001
R55750 S.n16617 S.t167 0.001
R55751 S.n16625 S.n16620 0.001
R55752 S.t187 S.n16641 0.001
R55753 S.t187 S.n16638 0.001
R55754 S.n16638 S.n16635 0.001
R55755 S.n15677 S.t60 0.001
R55756 S.n15685 S.n15680 0.001
R55757 S.t29 S.n15701 0.001
R55758 S.t29 S.n15698 0.001
R55759 S.n15698 S.n15695 0.001
R55760 S.n14724 S.t0 0.001
R55761 S.n14732 S.n14727 0.001
R55762 S.t102 S.n14748 0.001
R55763 S.t102 S.n14745 0.001
R55764 S.n14745 S.n14742 0.001
R55765 S.n13749 S.t73 0.001
R55766 S.n13757 S.n13752 0.001
R55767 S.t538 S.n13773 0.001
R55768 S.t538 S.n13770 0.001
R55769 S.n13770 S.n13767 0.001
R55770 S.n12761 S.t357 0.001
R55771 S.n12769 S.n12764 0.001
R55772 S.t443 S.n12785 0.001
R55773 S.t443 S.n12782 0.001
R55774 S.n12782 S.n12779 0.001
R55775 S.n11751 S.t54 0.001
R55776 S.n11759 S.n11754 0.001
R55777 S.t67 S.n11775 0.001
R55778 S.t67 S.n11772 0.001
R55779 S.n11772 S.n11769 0.001
R55780 S.n10728 S.t31 0.001
R55781 S.n10736 S.n10731 0.001
R55782 S.t172 S.n10752 0.001
R55783 S.t172 S.n10749 0.001
R55784 S.n10749 S.n10746 0.001
R55785 S.n9683 S.t366 0.001
R55786 S.n9691 S.n9686 0.001
R55787 S.t160 S.n9707 0.001
R55788 S.t160 S.n9704 0.001
R55789 S.n9704 S.n9701 0.001
R55790 S.n8625 S.t19 0.001
R55791 S.n8633 S.n8628 0.001
R55792 S.t141 S.n8649 0.001
R55793 S.t141 S.n8646 0.001
R55794 S.n8646 S.n8643 0.001
R55795 S.n7545 S.t47 0.001
R55796 S.n7553 S.n7548 0.001
R55797 S.t406 S.n7569 0.001
R55798 S.t406 S.n7566 0.001
R55799 S.n7566 S.n7563 0.001
R55800 S.n6452 S.t83 0.001
R55801 S.n6460 S.n6455 0.001
R55802 S.t130 S.n6476 0.001
R55803 S.t130 S.n6473 0.001
R55804 S.n6473 S.n6470 0.001
R55805 S.n5336 S.t214 0.001
R55806 S.n5344 S.n5339 0.001
R55807 S.t288 S.n5360 0.001
R55808 S.t288 S.n5357 0.001
R55809 S.n5357 S.n5354 0.001
R55810 S.n4207 S.t176 0.001
R55811 S.n4215 S.n4210 0.001
R55812 S.t134 S.n4231 0.001
R55813 S.t134 S.n4228 0.001
R55814 S.n4228 S.n4225 0.001
R55815 S.n3066 S.t14 0.001
R55816 S.n3074 S.n3069 0.001
R55817 S.t163 S.n3090 0.001
R55818 S.t163 S.n3087 0.001
R55819 S.n3087 S.n3084 0.001
R55820 S.t75 S.n1885 0.001
R55821 S.t75 S.n1888 0.001
R55822 S.t270 S.n1937 0.001
R55823 S.t270 S.n1934 0.001
R55824 S.n1934 S.n1931 0.001
R55825 S.t109 S.n412 0.001
R55826 S.t109 S.n409 0.001
R55827 S.n409 S.n406 0.001
R55828 S.t270 S.n2140 0.001
R55829 S.t270 S.n2143 0.001
R55830 S.t77 S.n18489 0.001
R55831 S.t77 S.n18486 0.001
R55832 S.n18486 S.n18483 0.001
R55833 S.t218 S.n17175 0.001
R55834 S.t218 S.n17172 0.001
R55835 S.n17172 S.n17169 0.001
R55836 S.t169 S.n17768 0.001
R55837 S.t169 S.n17771 0.001
R55838 S.t167 S.n16275 0.001
R55839 S.t167 S.n16272 0.001
R55840 S.n16272 S.n16269 0.001
R55841 S.t187 S.n16841 0.001
R55842 S.t187 S.n16844 0.001
R55843 S.t60 S.n15351 0.001
R55844 S.t60 S.n15348 0.001
R55845 S.n15348 S.n15345 0.001
R55846 S.t29 S.n15906 0.001
R55847 S.t29 S.n15909 0.001
R55848 S.t0 S.n14414 0.001
R55849 S.t0 S.n14411 0.001
R55850 S.n14411 S.n14408 0.001
R55851 S.t102 S.n14948 0.001
R55852 S.t102 S.n14951 0.001
R55853 S.t73 S.n13455 0.001
R55854 S.t73 S.n13452 0.001
R55855 S.n13452 S.n13449 0.001
R55856 S.t538 S.n13978 0.001
R55857 S.t538 S.n13981 0.001
R55858 S.t357 S.n12483 0.001
R55859 S.t357 S.n12480 0.001
R55860 S.n12480 S.n12477 0.001
R55861 S.t443 S.n12985 0.001
R55862 S.t443 S.n12988 0.001
R55863 S.t54 S.n11489 0.001
R55864 S.t54 S.n11486 0.001
R55865 S.n11486 S.n11483 0.001
R55866 S.t67 S.n11980 0.001
R55867 S.t67 S.n11983 0.001
R55868 S.t31 S.n10482 0.001
R55869 S.t31 S.n10479 0.001
R55870 S.n10479 S.n10476 0.001
R55871 S.t172 S.n10952 0.001
R55872 S.t172 S.n10955 0.001
R55873 S.t366 S.n9453 0.001
R55874 S.t366 S.n9450 0.001
R55875 S.n9450 S.n9447 0.001
R55876 S.t160 S.n9912 0.001
R55877 S.t160 S.n9915 0.001
R55878 S.t19 S.n8411 0.001
R55879 S.t19 S.n8408 0.001
R55880 S.n8408 S.n8405 0.001
R55881 S.t141 S.n8849 0.001
R55882 S.t141 S.n8852 0.001
R55883 S.t47 S.n7347 0.001
R55884 S.t47 S.n7344 0.001
R55885 S.n7344 S.n7341 0.001
R55886 S.t406 S.n7774 0.001
R55887 S.t406 S.n7777 0.001
R55888 S.t83 S.n6270 0.001
R55889 S.t83 S.n6267 0.001
R55890 S.n6267 S.n6264 0.001
R55891 S.t130 S.n6676 0.001
R55892 S.t130 S.n6679 0.001
R55893 S.t214 S.n5170 0.001
R55894 S.t214 S.n5167 0.001
R55895 S.n5167 S.n5164 0.001
R55896 S.t288 S.n5566 0.001
R55897 S.t288 S.n5569 0.001
R55898 S.t176 S.n4058 0.001
R55899 S.t176 S.n4055 0.001
R55900 S.n4055 S.n4052 0.001
R55901 S.t134 S.n4431 0.001
R55902 S.t134 S.n4434 0.001
R55903 S.t14 S.n2931 0.001
R55904 S.t14 S.n2928 0.001
R55905 S.n2928 S.n2925 0.001
R55906 S.t163 S.n3293 0.001
R55907 S.t163 S.n3296 0.001
R55908 S.t75 S.n1763 0.001
R55909 S.t75 S.n1760 0.001
R55910 S.n1760 S.n1757 0.001
R55911 S.n24 S.n19 0.001
R55912 S.t21 S.n19376 0.001
R55913 S.t21 S.n19373 0.001
R55914 S.n19373 S.n19370 0.001
R55915 S.t79 S.n18083 0.001
R55916 S.t79 S.n18080 0.001
R55917 S.n18080 S.n18077 0.001
R55918 S.t77 S.n18636 0.001
R55919 S.t77 S.n18639 0.001
R55920 S.t218 S.n17194 0.001
R55921 S.t218 S.n17191 0.001
R55922 S.n17191 S.n17188 0.001
R55923 S.t169 S.n17736 0.001
R55924 S.t169 S.n17739 0.001
R55925 S.t167 S.n16292 0.001
R55926 S.t167 S.n16289 0.001
R55927 S.n16289 S.n16286 0.001
R55928 S.t187 S.n16809 0.001
R55929 S.t187 S.n16812 0.001
R55930 S.t60 S.n15368 0.001
R55931 S.t60 S.n15365 0.001
R55932 S.n15365 S.n15362 0.001
R55933 S.t29 S.n15874 0.001
R55934 S.t29 S.n15877 0.001
R55935 S.t0 S.n14431 0.001
R55936 S.t0 S.n14428 0.001
R55937 S.n14428 S.n14425 0.001
R55938 S.t102 S.n14916 0.001
R55939 S.t102 S.n14919 0.001
R55940 S.t73 S.n13472 0.001
R55941 S.t73 S.n13469 0.001
R55942 S.n13469 S.n13466 0.001
R55943 S.t538 S.n13946 0.001
R55944 S.t538 S.n13949 0.001
R55945 S.t357 S.n12500 0.001
R55946 S.t357 S.n12497 0.001
R55947 S.n12497 S.n12494 0.001
R55948 S.t443 S.n12953 0.001
R55949 S.t443 S.n12956 0.001
R55950 S.t54 S.n11506 0.001
R55951 S.t54 S.n11503 0.001
R55952 S.n11503 S.n11500 0.001
R55953 S.t67 S.n11948 0.001
R55954 S.t67 S.n11951 0.001
R55955 S.t31 S.n10499 0.001
R55956 S.t31 S.n10496 0.001
R55957 S.n10496 S.n10493 0.001
R55958 S.t172 S.n10920 0.001
R55959 S.t172 S.n10923 0.001
R55960 S.t366 S.n9470 0.001
R55961 S.t366 S.n9467 0.001
R55962 S.n9467 S.n9464 0.001
R55963 S.t160 S.n9880 0.001
R55964 S.t160 S.n9883 0.001
R55965 S.t19 S.n8428 0.001
R55966 S.t19 S.n8425 0.001
R55967 S.n8425 S.n8422 0.001
R55968 S.t141 S.n8817 0.001
R55969 S.t141 S.n8820 0.001
R55970 S.t47 S.n7364 0.001
R55971 S.t47 S.n7361 0.001
R55972 S.n7361 S.n7358 0.001
R55973 S.t406 S.n7742 0.001
R55974 S.t406 S.n7745 0.001
R55975 S.t83 S.n6287 0.001
R55976 S.t83 S.n6284 0.001
R55977 S.n6284 S.n6281 0.001
R55978 S.t130 S.n6644 0.001
R55979 S.t130 S.n6647 0.001
R55980 S.t214 S.n5187 0.001
R55981 S.t214 S.n5184 0.001
R55982 S.n5184 S.n5181 0.001
R55983 S.t288 S.n5534 0.001
R55984 S.t288 S.n5537 0.001
R55985 S.t176 S.n4075 0.001
R55986 S.t176 S.n4072 0.001
R55987 S.n4072 S.n4069 0.001
R55988 S.t134 S.n4399 0.001
R55989 S.t134 S.n4402 0.001
R55990 S.t14 S.n2948 0.001
R55991 S.t14 S.n2945 0.001
R55992 S.n2945 S.n2942 0.001
R55993 S.t163 S.n3262 0.001
R55994 S.t163 S.n3265 0.001
R55995 S.t75 S.n1782 0.001
R55996 S.t75 S.n1779 0.001
R55997 S.n1779 S.n1776 0.001
R55998 S.t75 S.n1805 0.001
R55999 S.t75 S.n1802 0.001
R56000 S.n1802 S.n1799 0.001
R56001 S.t270 S.n2082 0.001
R56002 S.t270 S.n2085 0.001
R56003 S.n815 S.t137 0.001
R56004 S.n823 S.n818 0.001
R56005 S.t109 S.n844 0.001
R56006 S.t109 S.n841 0.001
R56007 S.n841 S.n838 0.001
R56008 S.t163 S.n3233 0.001
R56009 S.t163 S.n3236 0.001
R56010 S.t134 S.n4370 0.001
R56011 S.t134 S.n4373 0.001
R56012 S.t288 S.n5505 0.001
R56013 S.t288 S.n5508 0.001
R56014 S.t130 S.n6615 0.001
R56015 S.t130 S.n6618 0.001
R56016 S.t406 S.n7713 0.001
R56017 S.t406 S.n7716 0.001
R56018 S.t141 S.n8788 0.001
R56019 S.t141 S.n8791 0.001
R56020 S.t160 S.n9851 0.001
R56021 S.t160 S.n9854 0.001
R56022 S.t172 S.n10891 0.001
R56023 S.t172 S.n10894 0.001
R56024 S.t67 S.n11919 0.001
R56025 S.t67 S.n11922 0.001
R56026 S.t443 S.n12924 0.001
R56027 S.t443 S.n12927 0.001
R56028 S.t538 S.n13917 0.001
R56029 S.t538 S.n13920 0.001
R56030 S.t102 S.n14887 0.001
R56031 S.t102 S.n14890 0.001
R56032 S.t29 S.n15845 0.001
R56033 S.t29 S.n15848 0.001
R56034 S.t187 S.n16780 0.001
R56035 S.t187 S.n16783 0.001
R56036 S.t169 S.n17703 0.001
R56037 S.t169 S.n17706 0.001
R56038 S.t77 S.n18603 0.001
R56039 S.t77 S.n18606 0.001
R56040 S.t21 S.n19493 0.001
R56041 S.t21 S.n19496 0.001
R56042 S.t262 S.n20244 0.001
R56043 S.t262 S.n20241 0.001
R56044 S.n20241 S.n20238 0.001
R56045 S.t150 S.n18967 0.001
R56046 S.t150 S.n18964 0.001
R56047 S.n18964 S.n18961 0.001
R56048 S.t79 S.n18102 0.001
R56049 S.t79 S.n18099 0.001
R56050 S.n18099 S.n18096 0.001
R56051 S.t218 S.n17213 0.001
R56052 S.t218 S.n17210 0.001
R56053 S.n17210 S.n17207 0.001
R56054 S.t167 S.n16311 0.001
R56055 S.t167 S.n16308 0.001
R56056 S.n16308 S.n16305 0.001
R56057 S.t60 S.n15387 0.001
R56058 S.t60 S.n15384 0.001
R56059 S.n15384 S.n15381 0.001
R56060 S.t0 S.n14450 0.001
R56061 S.t0 S.n14447 0.001
R56062 S.n14447 S.n14444 0.001
R56063 S.t73 S.n13491 0.001
R56064 S.t73 S.n13488 0.001
R56065 S.n13488 S.n13485 0.001
R56066 S.t357 S.n12519 0.001
R56067 S.t357 S.n12516 0.001
R56068 S.n12516 S.n12513 0.001
R56069 S.t54 S.n11525 0.001
R56070 S.t54 S.n11522 0.001
R56071 S.n11522 S.n11519 0.001
R56072 S.t31 S.n10518 0.001
R56073 S.t31 S.n10515 0.001
R56074 S.n10515 S.n10512 0.001
R56075 S.t366 S.n9489 0.001
R56076 S.t366 S.n9486 0.001
R56077 S.n9486 S.n9483 0.001
R56078 S.t19 S.n8447 0.001
R56079 S.t19 S.n8444 0.001
R56080 S.n8444 S.n8441 0.001
R56081 S.t47 S.n7383 0.001
R56082 S.t47 S.n7380 0.001
R56083 S.n7380 S.n7377 0.001
R56084 S.t83 S.n6306 0.001
R56085 S.t83 S.n6303 0.001
R56086 S.n6303 S.n6300 0.001
R56087 S.t214 S.n5206 0.001
R56088 S.t214 S.n5203 0.001
R56089 S.n5203 S.n5200 0.001
R56090 S.t176 S.n4094 0.001
R56091 S.t176 S.n4091 0.001
R56092 S.n4091 S.n4088 0.001
R56093 S.t14 S.n2967 0.001
R56094 S.t14 S.n2964 0.001
R56095 S.n2964 S.n2961 0.001
R56096 S.t270 S.n2048 0.001
R56097 S.t270 S.n2051 0.001
R56098 S.t137 S.n773 0.001
R56099 S.t137 S.n770 0.001
R56100 S.n770 S.n767 0.001
R56101 S.n1337 S.n1331 0.001
R56102 S.t7 S.n20427 0.001
R56103 S.t7 S.n20430 0.001
R56104 S.t209 S.n19845 0.001
R56105 S.t209 S.n19842 0.001
R56106 S.n19842 S.n19839 0.001
R56107 S.t262 S.n20333 0.001
R56108 S.t262 S.n20336 0.001
R56109 S.t150 S.n18993 0.001
R56110 S.t150 S.n18990 0.001
R56111 S.n18990 S.n18987 0.001
R56112 S.t21 S.n19461 0.001
R56113 S.t21 S.n19464 0.001
R56114 S.t79 S.n18127 0.001
R56115 S.t79 S.n18124 0.001
R56116 S.n18124 S.n18121 0.001
R56117 S.t77 S.n18571 0.001
R56118 S.t77 S.n18574 0.001
R56119 S.t218 S.n17238 0.001
R56120 S.t218 S.n17235 0.001
R56121 S.n17235 S.n17232 0.001
R56122 S.t169 S.n17671 0.001
R56123 S.t169 S.n17674 0.001
R56124 S.t167 S.n16336 0.001
R56125 S.t167 S.n16333 0.001
R56126 S.n16333 S.n16330 0.001
R56127 S.t187 S.n16748 0.001
R56128 S.t187 S.n16751 0.001
R56129 S.t60 S.n15412 0.001
R56130 S.t60 S.n15409 0.001
R56131 S.n15409 S.n15406 0.001
R56132 S.t29 S.n15813 0.001
R56133 S.t29 S.n15816 0.001
R56134 S.t0 S.n14475 0.001
R56135 S.t0 S.n14472 0.001
R56136 S.n14472 S.n14469 0.001
R56137 S.t102 S.n14855 0.001
R56138 S.t102 S.n14858 0.001
R56139 S.t73 S.n13516 0.001
R56140 S.t73 S.n13513 0.001
R56141 S.n13513 S.n13510 0.001
R56142 S.t538 S.n13885 0.001
R56143 S.t538 S.n13888 0.001
R56144 S.t357 S.n12544 0.001
R56145 S.t357 S.n12541 0.001
R56146 S.n12541 S.n12538 0.001
R56147 S.t443 S.n12892 0.001
R56148 S.t443 S.n12895 0.001
R56149 S.t54 S.n11550 0.001
R56150 S.t54 S.n11547 0.001
R56151 S.n11547 S.n11544 0.001
R56152 S.t67 S.n11887 0.001
R56153 S.t67 S.n11890 0.001
R56154 S.t31 S.n10543 0.001
R56155 S.t31 S.n10540 0.001
R56156 S.n10540 S.n10537 0.001
R56157 S.t172 S.n10859 0.001
R56158 S.t172 S.n10862 0.001
R56159 S.t366 S.n9514 0.001
R56160 S.t366 S.n9511 0.001
R56161 S.n9511 S.n9508 0.001
R56162 S.t160 S.n9819 0.001
R56163 S.t160 S.n9822 0.001
R56164 S.t19 S.n8472 0.001
R56165 S.t19 S.n8469 0.001
R56166 S.n8469 S.n8466 0.001
R56167 S.t141 S.n8756 0.001
R56168 S.t141 S.n8759 0.001
R56169 S.t47 S.n7408 0.001
R56170 S.t47 S.n7405 0.001
R56171 S.n7405 S.n7402 0.001
R56172 S.t406 S.n7681 0.001
R56173 S.t406 S.n7684 0.001
R56174 S.t83 S.n6331 0.001
R56175 S.t83 S.n6328 0.001
R56176 S.n6328 S.n6325 0.001
R56177 S.t130 S.n6583 0.001
R56178 S.t130 S.n6586 0.001
R56179 S.t214 S.n5231 0.001
R56180 S.t214 S.n5228 0.001
R56181 S.n5228 S.n5225 0.001
R56182 S.t288 S.n5473 0.001
R56183 S.t288 S.n5476 0.001
R56184 S.t176 S.n4119 0.001
R56185 S.t176 S.n4116 0.001
R56186 S.n4116 S.n4113 0.001
R56187 S.t134 S.n4338 0.001
R56188 S.t134 S.n4341 0.001
R56189 S.t14 S.n2992 0.001
R56190 S.t14 S.n2989 0.001
R56191 S.n2989 S.n2986 0.001
R56192 S.t163 S.n3201 0.001
R56193 S.t163 S.n3204 0.001
R56194 S.t75 S.n1829 0.001
R56195 S.t75 S.n1826 0.001
R56196 S.n1826 S.n1823 0.001
R56197 S.t270 S.n2015 0.001
R56198 S.t270 S.n2018 0.001
R56199 S.t137 S.n792 0.001
R56200 S.t137 S.n789 0.001
R56201 S.n789 S.n786 0.001
R56202 S.t75 S.n1851 0.001
R56203 S.t75 S.n1848 0.001
R56204 S.n1848 S.n1845 0.001
R56205 S.t163 S.n3169 0.001
R56206 S.t163 S.n3172 0.001
R56207 S.t14 S.n3012 0.001
R56208 S.t14 S.n3009 0.001
R56209 S.n3009 S.n3006 0.001
R56210 S.t134 S.n4306 0.001
R56211 S.t134 S.n4309 0.001
R56212 S.t176 S.n4138 0.001
R56213 S.t176 S.n4135 0.001
R56214 S.n4135 S.n4132 0.001
R56215 S.t288 S.n5441 0.001
R56216 S.t288 S.n5444 0.001
R56217 S.t214 S.n5251 0.001
R56218 S.t214 S.n5248 0.001
R56219 S.n5248 S.n5245 0.001
R56220 S.t130 S.n6551 0.001
R56221 S.t130 S.n6554 0.001
R56222 S.t83 S.n6351 0.001
R56223 S.t83 S.n6348 0.001
R56224 S.n6348 S.n6345 0.001
R56225 S.t406 S.n7649 0.001
R56226 S.t406 S.n7652 0.001
R56227 S.t47 S.n7428 0.001
R56228 S.t47 S.n7425 0.001
R56229 S.n7425 S.n7422 0.001
R56230 S.t141 S.n8724 0.001
R56231 S.t141 S.n8727 0.001
R56232 S.t19 S.n8492 0.001
R56233 S.t19 S.n8489 0.001
R56234 S.n8489 S.n8486 0.001
R56235 S.t160 S.n9787 0.001
R56236 S.t160 S.n9790 0.001
R56237 S.t366 S.n9534 0.001
R56238 S.t366 S.n9531 0.001
R56239 S.n9531 S.n9528 0.001
R56240 S.t172 S.n10827 0.001
R56241 S.t172 S.n10830 0.001
R56242 S.t31 S.n10563 0.001
R56243 S.t31 S.n10560 0.001
R56244 S.n10560 S.n10557 0.001
R56245 S.t67 S.n11855 0.001
R56246 S.t67 S.n11858 0.001
R56247 S.t54 S.n11570 0.001
R56248 S.t54 S.n11567 0.001
R56249 S.n11567 S.n11564 0.001
R56250 S.t443 S.n12860 0.001
R56251 S.t443 S.n12863 0.001
R56252 S.t357 S.n12564 0.001
R56253 S.t357 S.n12561 0.001
R56254 S.n12561 S.n12558 0.001
R56255 S.t538 S.n13853 0.001
R56256 S.t538 S.n13856 0.001
R56257 S.t73 S.n13536 0.001
R56258 S.t73 S.n13533 0.001
R56259 S.n13533 S.n13530 0.001
R56260 S.t102 S.n14823 0.001
R56261 S.t102 S.n14826 0.001
R56262 S.t0 S.n14495 0.001
R56263 S.t0 S.n14492 0.001
R56264 S.n14492 S.n14489 0.001
R56265 S.t29 S.n15781 0.001
R56266 S.t29 S.n15784 0.001
R56267 S.t60 S.n15432 0.001
R56268 S.t60 S.n15429 0.001
R56269 S.n15429 S.n15426 0.001
R56270 S.t187 S.n16716 0.001
R56271 S.t187 S.n16719 0.001
R56272 S.t167 S.n16356 0.001
R56273 S.t167 S.n16353 0.001
R56274 S.n16353 S.n16350 0.001
R56275 S.t169 S.n17639 0.001
R56276 S.t169 S.n17642 0.001
R56277 S.t218 S.n17258 0.001
R56278 S.t218 S.n17255 0.001
R56279 S.n17255 S.n17252 0.001
R56280 S.t77 S.n18539 0.001
R56281 S.t77 S.n18542 0.001
R56282 S.t79 S.n18147 0.001
R56283 S.t79 S.n18144 0.001
R56284 S.n18144 S.n18141 0.001
R56285 S.t21 S.n19426 0.001
R56286 S.t21 S.n19429 0.001
R56287 S.t150 S.n19013 0.001
R56288 S.t150 S.n19010 0.001
R56289 S.n19010 S.n19007 0.001
R56290 S.t262 S.n20298 0.001
R56291 S.t262 S.n20301 0.001
R56292 S.t209 S.n19867 0.001
R56293 S.t209 S.n19864 0.001
R56294 S.n19864 S.n19861 0.001
R56295 S.t7 S.n20372 0.001
R56296 S.t7 S.n20369 0.001
R56297 S.n20369 S.n20366 0.001
R56298 S.t64 S.n20478 0.001
R56299 S.t64 S.n20475 0.001
R56300 S.n20475 S.n20472 0.001
R56301 S.t105 S.n21245 0.001
R56302 S.t105 S.n21248 0.001
R56303 S.t109 S.n870 0.001
R56304 S.t109 S.n867 0.001
R56305 S.n867 S.n864 0.001
R56306 S.t270 S.n2110 0.001
R56307 S.t270 S.n2113 0.001
R56308 S.t137 S.n749 0.001
R56309 S.t137 S.n746 0.001
R56310 S.n746 S.n743 0.001
R56311 S.t137 S.n732 0.001
R56312 S.t137 S.n729 0.001
R56313 S.n729 S.n726 0.001
R56314 S.t109 S.n380 0.001
R56315 S.t109 S.n377 0.001
R56316 S.n377 S.n374 0.001
R56317 S.t270 S.n2199 0.001
R56318 S.t270 S.n2202 0.001
R56319 S.t187 S.n16666 0.001
R56320 S.t187 S.n16663 0.001
R56321 S.n16663 S.n16660 0.001
R56322 S.t60 S.n15313 0.001
R56323 S.t60 S.n15310 0.001
R56324 S.n15310 S.n15307 0.001
R56325 S.t29 S.n15971 0.001
R56326 S.t29 S.n15974 0.001
R56327 S.t0 S.n14378 0.001
R56328 S.t0 S.n14375 0.001
R56329 S.n14375 S.n14372 0.001
R56330 S.t102 S.n15009 0.001
R56331 S.t102 S.n15012 0.001
R56332 S.t73 S.n13419 0.001
R56333 S.t73 S.n13416 0.001
R56334 S.n13416 S.n13413 0.001
R56335 S.t538 S.n14039 0.001
R56336 S.t538 S.n14042 0.001
R56337 S.t357 S.n12447 0.001
R56338 S.t357 S.n12444 0.001
R56339 S.n12444 S.n12441 0.001
R56340 S.t443 S.n13046 0.001
R56341 S.t443 S.n13049 0.001
R56342 S.t54 S.n11453 0.001
R56343 S.t54 S.n11450 0.001
R56344 S.n11450 S.n11447 0.001
R56345 S.t67 S.n12041 0.001
R56346 S.t67 S.n12044 0.001
R56347 S.t31 S.n10446 0.001
R56348 S.t31 S.n10443 0.001
R56349 S.n10443 S.n10440 0.001
R56350 S.t172 S.n11013 0.001
R56351 S.t172 S.n11016 0.001
R56352 S.t366 S.n9417 0.001
R56353 S.t366 S.n9414 0.001
R56354 S.n9414 S.n9411 0.001
R56355 S.t160 S.n9973 0.001
R56356 S.t160 S.n9976 0.001
R56357 S.t19 S.n8375 0.001
R56358 S.t19 S.n8372 0.001
R56359 S.n8372 S.n8369 0.001
R56360 S.t141 S.n8910 0.001
R56361 S.t141 S.n8913 0.001
R56362 S.t47 S.n7311 0.001
R56363 S.t47 S.n7308 0.001
R56364 S.n7308 S.n7305 0.001
R56365 S.t406 S.n7835 0.001
R56366 S.t406 S.n7838 0.001
R56367 S.t83 S.n6234 0.001
R56368 S.t83 S.n6231 0.001
R56369 S.n6231 S.n6228 0.001
R56370 S.t130 S.n6737 0.001
R56371 S.t130 S.n6740 0.001
R56372 S.t214 S.n5134 0.001
R56373 S.t214 S.n5131 0.001
R56374 S.n5131 S.n5128 0.001
R56375 S.t288 S.n5627 0.001
R56376 S.t288 S.n5630 0.001
R56377 S.t176 S.n4022 0.001
R56378 S.t176 S.n4019 0.001
R56379 S.n4019 S.n4016 0.001
R56380 S.t134 S.n4492 0.001
R56381 S.t134 S.n4495 0.001
R56382 S.t14 S.n2895 0.001
R56383 S.t14 S.n2892 0.001
R56384 S.n2892 S.n2889 0.001
R56385 S.t163 S.n3353 0.001
R56386 S.t163 S.n3356 0.001
R56387 S.t75 S.n1726 0.001
R56388 S.t75 S.n1723 0.001
R56389 S.n1723 S.n1720 0.001
R56390 S.n71 S.n66 0.001
R56391 S.t169 S.n17589 0.001
R56392 S.t169 S.n17586 0.001
R56393 S.n17586 S.n17583 0.001
R56394 S.t167 S.n16256 0.001
R56395 S.t167 S.n16253 0.001
R56396 S.n16253 S.n16250 0.001
R56397 S.t187 S.n16874 0.001
R56398 S.t187 S.n16877 0.001
R56399 S.t60 S.n15332 0.001
R56400 S.t60 S.n15329 0.001
R56401 S.n15329 S.n15326 0.001
R56402 S.t29 S.n15939 0.001
R56403 S.t29 S.n15942 0.001
R56404 S.t0 S.n14395 0.001
R56405 S.t0 S.n14392 0.001
R56406 S.n14392 S.n14389 0.001
R56407 S.t102 S.n14977 0.001
R56408 S.t102 S.n14980 0.001
R56409 S.t73 S.n13436 0.001
R56410 S.t73 S.n13433 0.001
R56411 S.n13433 S.n13430 0.001
R56412 S.t538 S.n14007 0.001
R56413 S.t538 S.n14010 0.001
R56414 S.t357 S.n12464 0.001
R56415 S.t357 S.n12461 0.001
R56416 S.n12461 S.n12458 0.001
R56417 S.t443 S.n13014 0.001
R56418 S.t443 S.n13017 0.001
R56419 S.t54 S.n11470 0.001
R56420 S.t54 S.n11467 0.001
R56421 S.n11467 S.n11464 0.001
R56422 S.t67 S.n12009 0.001
R56423 S.t67 S.n12012 0.001
R56424 S.t31 S.n10463 0.001
R56425 S.t31 S.n10460 0.001
R56426 S.n10460 S.n10457 0.001
R56427 S.t172 S.n10981 0.001
R56428 S.t172 S.n10984 0.001
R56429 S.t366 S.n9434 0.001
R56430 S.t366 S.n9431 0.001
R56431 S.n9431 S.n9428 0.001
R56432 S.t160 S.n9941 0.001
R56433 S.t160 S.n9944 0.001
R56434 S.t19 S.n8392 0.001
R56435 S.t19 S.n8389 0.001
R56436 S.n8389 S.n8386 0.001
R56437 S.t141 S.n8878 0.001
R56438 S.t141 S.n8881 0.001
R56439 S.t47 S.n7328 0.001
R56440 S.t47 S.n7325 0.001
R56441 S.n7325 S.n7322 0.001
R56442 S.t406 S.n7803 0.001
R56443 S.t406 S.n7806 0.001
R56444 S.t83 S.n6251 0.001
R56445 S.t83 S.n6248 0.001
R56446 S.n6248 S.n6245 0.001
R56447 S.t130 S.n6705 0.001
R56448 S.t130 S.n6708 0.001
R56449 S.t214 S.n5151 0.001
R56450 S.t214 S.n5148 0.001
R56451 S.n5148 S.n5145 0.001
R56452 S.t288 S.n5595 0.001
R56453 S.t288 S.n5598 0.001
R56454 S.t176 S.n4039 0.001
R56455 S.t176 S.n4036 0.001
R56456 S.n4036 S.n4033 0.001
R56457 S.t134 S.n4460 0.001
R56458 S.t134 S.n4463 0.001
R56459 S.t14 S.n2912 0.001
R56460 S.t14 S.n2909 0.001
R56461 S.n2909 S.n2906 0.001
R56462 S.t163 S.n3322 0.001
R56463 S.t163 S.n3325 0.001
R56464 S.t75 S.n1743 0.001
R56465 S.t75 S.n1740 0.001
R56466 S.n1740 S.n1737 0.001
R56467 S.t270 S.n2169 0.001
R56468 S.t270 S.n2172 0.001
R56469 S.t137 S.n714 0.001
R56470 S.t137 S.n711 0.001
R56471 S.n711 S.n708 0.001
R56472 S.t137 S.n697 0.001
R56473 S.t137 S.n694 0.001
R56474 S.n694 S.n691 0.001
R56475 S.t109 S.n348 0.001
R56476 S.t109 S.n345 0.001
R56477 S.n345 S.n342 0.001
R56478 S.t270 S.n2258 0.001
R56479 S.t270 S.n2261 0.001
R56480 S.t102 S.n14773 0.001
R56481 S.t102 S.n14770 0.001
R56482 S.n14770 S.n14767 0.001
R56483 S.t73 S.n13381 0.001
R56484 S.t73 S.n13378 0.001
R56485 S.n13378 S.n13375 0.001
R56486 S.t538 S.n14104 0.001
R56487 S.t538 S.n14107 0.001
R56488 S.t357 S.n12411 0.001
R56489 S.t357 S.n12408 0.001
R56490 S.n12408 S.n12405 0.001
R56491 S.t443 S.n13107 0.001
R56492 S.t443 S.n13110 0.001
R56493 S.t54 S.n11417 0.001
R56494 S.t54 S.n11414 0.001
R56495 S.n11414 S.n11411 0.001
R56496 S.t67 S.n12102 0.001
R56497 S.t67 S.n12105 0.001
R56498 S.t31 S.n10410 0.001
R56499 S.t31 S.n10407 0.001
R56500 S.n10407 S.n10404 0.001
R56501 S.t172 S.n11074 0.001
R56502 S.t172 S.n11077 0.001
R56503 S.t366 S.n9381 0.001
R56504 S.t366 S.n9378 0.001
R56505 S.n9378 S.n9375 0.001
R56506 S.t160 S.n10034 0.001
R56507 S.t160 S.n10037 0.001
R56508 S.t19 S.n8339 0.001
R56509 S.t19 S.n8336 0.001
R56510 S.n8336 S.n8333 0.001
R56511 S.t141 S.n8971 0.001
R56512 S.t141 S.n8974 0.001
R56513 S.t47 S.n7275 0.001
R56514 S.t47 S.n7272 0.001
R56515 S.n7272 S.n7269 0.001
R56516 S.t406 S.n7896 0.001
R56517 S.t406 S.n7899 0.001
R56518 S.t83 S.n6198 0.001
R56519 S.t83 S.n6195 0.001
R56520 S.n6195 S.n6192 0.001
R56521 S.t130 S.n6798 0.001
R56522 S.t130 S.n6801 0.001
R56523 S.t214 S.n5098 0.001
R56524 S.t214 S.n5095 0.001
R56525 S.n5095 S.n5092 0.001
R56526 S.t288 S.n5688 0.001
R56527 S.t288 S.n5691 0.001
R56528 S.t176 S.n3986 0.001
R56529 S.t176 S.n3983 0.001
R56530 S.n3983 S.n3980 0.001
R56531 S.t134 S.n4553 0.001
R56532 S.t134 S.n4556 0.001
R56533 S.t14 S.n2859 0.001
R56534 S.t14 S.n2856 0.001
R56535 S.n2856 S.n2853 0.001
R56536 S.t163 S.n3413 0.001
R56537 S.t163 S.n3416 0.001
R56538 S.t75 S.n1689 0.001
R56539 S.t75 S.n1686 0.001
R56540 S.n1686 S.n1683 0.001
R56541 S.n103 S.n98 0.001
R56542 S.t29 S.n15731 0.001
R56543 S.t29 S.n15728 0.001
R56544 S.n15728 S.n15725 0.001
R56545 S.t0 S.n14359 0.001
R56546 S.t0 S.n14356 0.001
R56547 S.n14356 S.n14353 0.001
R56548 S.t102 S.n15042 0.001
R56549 S.t102 S.n15045 0.001
R56550 S.t73 S.n13400 0.001
R56551 S.t73 S.n13397 0.001
R56552 S.n13397 S.n13394 0.001
R56553 S.t538 S.n14072 0.001
R56554 S.t538 S.n14075 0.001
R56555 S.t357 S.n12428 0.001
R56556 S.t357 S.n12425 0.001
R56557 S.n12425 S.n12422 0.001
R56558 S.t443 S.n13075 0.001
R56559 S.t443 S.n13078 0.001
R56560 S.t54 S.n11434 0.001
R56561 S.t54 S.n11431 0.001
R56562 S.n11431 S.n11428 0.001
R56563 S.t67 S.n12070 0.001
R56564 S.t67 S.n12073 0.001
R56565 S.t31 S.n10427 0.001
R56566 S.t31 S.n10424 0.001
R56567 S.n10424 S.n10421 0.001
R56568 S.t172 S.n11042 0.001
R56569 S.t172 S.n11045 0.001
R56570 S.t366 S.n9398 0.001
R56571 S.t366 S.n9395 0.001
R56572 S.n9395 S.n9392 0.001
R56573 S.t160 S.n10002 0.001
R56574 S.t160 S.n10005 0.001
R56575 S.t19 S.n8356 0.001
R56576 S.t19 S.n8353 0.001
R56577 S.n8353 S.n8350 0.001
R56578 S.t141 S.n8939 0.001
R56579 S.t141 S.n8942 0.001
R56580 S.t47 S.n7292 0.001
R56581 S.t47 S.n7289 0.001
R56582 S.n7289 S.n7286 0.001
R56583 S.t406 S.n7864 0.001
R56584 S.t406 S.n7867 0.001
R56585 S.t83 S.n6215 0.001
R56586 S.t83 S.n6212 0.001
R56587 S.n6212 S.n6209 0.001
R56588 S.t130 S.n6766 0.001
R56589 S.t130 S.n6769 0.001
R56590 S.t214 S.n5115 0.001
R56591 S.t214 S.n5112 0.001
R56592 S.n5112 S.n5109 0.001
R56593 S.t288 S.n5656 0.001
R56594 S.t288 S.n5659 0.001
R56595 S.t176 S.n4003 0.001
R56596 S.t176 S.n4000 0.001
R56597 S.n4000 S.n3997 0.001
R56598 S.t134 S.n4521 0.001
R56599 S.t134 S.n4524 0.001
R56600 S.t14 S.n2876 0.001
R56601 S.t14 S.n2873 0.001
R56602 S.n2873 S.n2870 0.001
R56603 S.t163 S.n3382 0.001
R56604 S.t163 S.n3385 0.001
R56605 S.t75 S.n1706 0.001
R56606 S.t75 S.n1703 0.001
R56607 S.n1703 S.n1700 0.001
R56608 S.t270 S.n2228 0.001
R56609 S.t270 S.n2231 0.001
R56610 S.t137 S.n679 0.001
R56611 S.t137 S.n676 0.001
R56612 S.n676 S.n673 0.001
R56613 S.t137 S.n662 0.001
R56614 S.t137 S.n659 0.001
R56615 S.n659 S.n656 0.001
R56616 S.t109 S.n316 0.001
R56617 S.t109 S.n313 0.001
R56618 S.n313 S.n310 0.001
R56619 S.t270 S.n2317 0.001
R56620 S.t270 S.n2320 0.001
R56621 S.t443 S.n12810 0.001
R56622 S.t443 S.n12807 0.001
R56623 S.n12807 S.n12804 0.001
R56624 S.t54 S.n11379 0.001
R56625 S.t54 S.n11376 0.001
R56626 S.n11376 S.n11373 0.001
R56627 S.t67 S.n12167 0.001
R56628 S.t67 S.n12170 0.001
R56629 S.t31 S.n10374 0.001
R56630 S.t31 S.n10371 0.001
R56631 S.n10371 S.n10368 0.001
R56632 S.t172 S.n11135 0.001
R56633 S.t172 S.n11138 0.001
R56634 S.t366 S.n9345 0.001
R56635 S.t366 S.n9342 0.001
R56636 S.n9342 S.n9339 0.001
R56637 S.t160 S.n10095 0.001
R56638 S.t160 S.n10098 0.001
R56639 S.t19 S.n8303 0.001
R56640 S.t19 S.n8300 0.001
R56641 S.n8300 S.n8297 0.001
R56642 S.t141 S.n9032 0.001
R56643 S.t141 S.n9035 0.001
R56644 S.t47 S.n7239 0.001
R56645 S.t47 S.n7236 0.001
R56646 S.n7236 S.n7233 0.001
R56647 S.t406 S.n7957 0.001
R56648 S.t406 S.n7960 0.001
R56649 S.t83 S.n6162 0.001
R56650 S.t83 S.n6159 0.001
R56651 S.n6159 S.n6156 0.001
R56652 S.t130 S.n6859 0.001
R56653 S.t130 S.n6862 0.001
R56654 S.t214 S.n5062 0.001
R56655 S.t214 S.n5059 0.001
R56656 S.n5059 S.n5056 0.001
R56657 S.t288 S.n5749 0.001
R56658 S.t288 S.n5752 0.001
R56659 S.t176 S.n3950 0.001
R56660 S.t176 S.n3947 0.001
R56661 S.n3947 S.n3944 0.001
R56662 S.t134 S.n4614 0.001
R56663 S.t134 S.n4617 0.001
R56664 S.t14 S.n2823 0.001
R56665 S.t14 S.n2820 0.001
R56666 S.n2820 S.n2817 0.001
R56667 S.t163 S.n3473 0.001
R56668 S.t163 S.n3476 0.001
R56669 S.t75 S.n1652 0.001
R56670 S.t75 S.n1649 0.001
R56671 S.n1649 S.n1646 0.001
R56672 S.n982 S.t109 0.001
R56673 S.n990 S.n985 0.001
R56674 S.t538 S.n13803 0.001
R56675 S.t538 S.n13800 0.001
R56676 S.n13800 S.n13797 0.001
R56677 S.t357 S.n12392 0.001
R56678 S.t357 S.n12389 0.001
R56679 S.n12389 S.n12386 0.001
R56680 S.t443 S.n13140 0.001
R56681 S.t443 S.n13143 0.001
R56682 S.t54 S.n11398 0.001
R56683 S.t54 S.n11395 0.001
R56684 S.n11395 S.n11392 0.001
R56685 S.t67 S.n12135 0.001
R56686 S.t67 S.n12138 0.001
R56687 S.t31 S.n10391 0.001
R56688 S.t31 S.n10388 0.001
R56689 S.n10388 S.n10385 0.001
R56690 S.t172 S.n11103 0.001
R56691 S.t172 S.n11106 0.001
R56692 S.t366 S.n9362 0.001
R56693 S.t366 S.n9359 0.001
R56694 S.n9359 S.n9356 0.001
R56695 S.t160 S.n10063 0.001
R56696 S.t160 S.n10066 0.001
R56697 S.t19 S.n8320 0.001
R56698 S.t19 S.n8317 0.001
R56699 S.n8317 S.n8314 0.001
R56700 S.t141 S.n9000 0.001
R56701 S.t141 S.n9003 0.001
R56702 S.t47 S.n7256 0.001
R56703 S.t47 S.n7253 0.001
R56704 S.n7253 S.n7250 0.001
R56705 S.t406 S.n7925 0.001
R56706 S.t406 S.n7928 0.001
R56707 S.t83 S.n6179 0.001
R56708 S.t83 S.n6176 0.001
R56709 S.n6176 S.n6173 0.001
R56710 S.t130 S.n6827 0.001
R56711 S.t130 S.n6830 0.001
R56712 S.t214 S.n5079 0.001
R56713 S.t214 S.n5076 0.001
R56714 S.n5076 S.n5073 0.001
R56715 S.t288 S.n5717 0.001
R56716 S.t288 S.n5720 0.001
R56717 S.t176 S.n3967 0.001
R56718 S.t176 S.n3964 0.001
R56719 S.n3964 S.n3961 0.001
R56720 S.t134 S.n4582 0.001
R56721 S.t134 S.n4585 0.001
R56722 S.t14 S.n2840 0.001
R56723 S.t14 S.n2837 0.001
R56724 S.n2837 S.n2834 0.001
R56725 S.t163 S.n3442 0.001
R56726 S.t163 S.n3445 0.001
R56727 S.t75 S.n1669 0.001
R56728 S.t75 S.n1666 0.001
R56729 S.n1666 S.n1663 0.001
R56730 S.t270 S.n2287 0.001
R56731 S.t270 S.n2290 0.001
R56732 S.t137 S.n644 0.001
R56733 S.t137 S.n641 0.001
R56734 S.n641 S.n638 0.001
R56735 S.t137 S.n627 0.001
R56736 S.t137 S.n624 0.001
R56737 S.n624 S.n621 0.001
R56738 S.t109 S.n284 0.001
R56739 S.t109 S.n281 0.001
R56740 S.n281 S.n278 0.001
R56741 S.t270 S.n2376 0.001
R56742 S.t270 S.n2379 0.001
R56743 S.t172 S.n10777 0.001
R56744 S.t172 S.n10774 0.001
R56745 S.n10774 S.n10771 0.001
R56746 S.t366 S.n9307 0.001
R56747 S.t366 S.n9304 0.001
R56748 S.n9304 S.n9301 0.001
R56749 S.t160 S.n10160 0.001
R56750 S.t160 S.n10163 0.001
R56751 S.t19 S.n8267 0.001
R56752 S.t19 S.n8264 0.001
R56753 S.n8264 S.n8261 0.001
R56754 S.t141 S.n9093 0.001
R56755 S.t141 S.n9096 0.001
R56756 S.t47 S.n7203 0.001
R56757 S.t47 S.n7200 0.001
R56758 S.n7200 S.n7197 0.001
R56759 S.t406 S.n8018 0.001
R56760 S.t406 S.n8021 0.001
R56761 S.t83 S.n6126 0.001
R56762 S.t83 S.n6123 0.001
R56763 S.n6123 S.n6120 0.001
R56764 S.t130 S.n6920 0.001
R56765 S.t130 S.n6923 0.001
R56766 S.t214 S.n5026 0.001
R56767 S.t214 S.n5023 0.001
R56768 S.n5023 S.n5020 0.001
R56769 S.t288 S.n5810 0.001
R56770 S.t288 S.n5813 0.001
R56771 S.t176 S.n3914 0.001
R56772 S.t176 S.n3911 0.001
R56773 S.n3911 S.n3908 0.001
R56774 S.t134 S.n4675 0.001
R56775 S.t134 S.n4678 0.001
R56776 S.t14 S.n2787 0.001
R56777 S.t14 S.n2784 0.001
R56778 S.n2784 S.n2781 0.001
R56779 S.t163 S.n3533 0.001
R56780 S.t163 S.n3536 0.001
R56781 S.t75 S.n1615 0.001
R56782 S.t75 S.n1612 0.001
R56783 S.n1612 S.n1609 0.001
R56784 S.n1022 S.n1017 0.001
R56785 S.t67 S.n11805 0.001
R56786 S.t67 S.n11802 0.001
R56787 S.n11802 S.n11799 0.001
R56788 S.t31 S.n10355 0.001
R56789 S.t31 S.n10352 0.001
R56790 S.n10352 S.n10349 0.001
R56791 S.t172 S.n11168 0.001
R56792 S.t172 S.n11171 0.001
R56793 S.t366 S.n9326 0.001
R56794 S.t366 S.n9323 0.001
R56795 S.n9323 S.n9320 0.001
R56796 S.t160 S.n10128 0.001
R56797 S.t160 S.n10131 0.001
R56798 S.t19 S.n8284 0.001
R56799 S.t19 S.n8281 0.001
R56800 S.n8281 S.n8278 0.001
R56801 S.t141 S.n9061 0.001
R56802 S.t141 S.n9064 0.001
R56803 S.t47 S.n7220 0.001
R56804 S.t47 S.n7217 0.001
R56805 S.n7217 S.n7214 0.001
R56806 S.t406 S.n7986 0.001
R56807 S.t406 S.n7989 0.001
R56808 S.t83 S.n6143 0.001
R56809 S.t83 S.n6140 0.001
R56810 S.n6140 S.n6137 0.001
R56811 S.t130 S.n6888 0.001
R56812 S.t130 S.n6891 0.001
R56813 S.t214 S.n5043 0.001
R56814 S.t214 S.n5040 0.001
R56815 S.n5040 S.n5037 0.001
R56816 S.t288 S.n5778 0.001
R56817 S.t288 S.n5781 0.001
R56818 S.t176 S.n3931 0.001
R56819 S.t176 S.n3928 0.001
R56820 S.n3928 S.n3925 0.001
R56821 S.t134 S.n4643 0.001
R56822 S.t134 S.n4646 0.001
R56823 S.t14 S.n2804 0.001
R56824 S.t14 S.n2801 0.001
R56825 S.n2801 S.n2798 0.001
R56826 S.t163 S.n3502 0.001
R56827 S.t163 S.n3505 0.001
R56828 S.t75 S.n1632 0.001
R56829 S.t75 S.n1629 0.001
R56830 S.n1629 S.n1626 0.001
R56831 S.t270 S.n2346 0.001
R56832 S.t270 S.n2349 0.001
R56833 S.t137 S.n609 0.001
R56834 S.t137 S.n606 0.001
R56835 S.n606 S.n603 0.001
R56836 S.t137 S.n592 0.001
R56837 S.t137 S.n589 0.001
R56838 S.n589 S.n586 0.001
R56839 S.t109 S.n252 0.001
R56840 S.t109 S.n223 0.001
R56841 S.t270 S.n2435 0.001
R56842 S.t270 S.n2438 0.001
R56843 S.t141 S.n8674 0.001
R56844 S.t141 S.n8671 0.001
R56845 S.n8671 S.n8668 0.001
R56846 S.t47 S.n7165 0.001
R56847 S.t47 S.n7162 0.001
R56848 S.n7162 S.n7159 0.001
R56849 S.t406 S.n8083 0.001
R56850 S.t406 S.n8086 0.001
R56851 S.t83 S.n6090 0.001
R56852 S.t83 S.n6087 0.001
R56853 S.n6087 S.n6084 0.001
R56854 S.t130 S.n6981 0.001
R56855 S.t130 S.n6984 0.001
R56856 S.t214 S.n4990 0.001
R56857 S.t214 S.n4987 0.001
R56858 S.n4987 S.n4984 0.001
R56859 S.t288 S.n5871 0.001
R56860 S.t288 S.n5874 0.001
R56861 S.t176 S.n3878 0.001
R56862 S.t176 S.n3875 0.001
R56863 S.n3875 S.n3872 0.001
R56864 S.t134 S.n4736 0.001
R56865 S.t134 S.n4739 0.001
R56866 S.t14 S.n2751 0.001
R56867 S.t14 S.n2748 0.001
R56868 S.n2748 S.n2745 0.001
R56869 S.t163 S.n3593 0.001
R56870 S.t163 S.n3596 0.001
R56871 S.t75 S.n1578 0.001
R56872 S.t75 S.n1575 0.001
R56873 S.n1575 S.n1572 0.001
R56874 S.n1054 S.n1049 0.001
R56875 S.t160 S.n9737 0.001
R56876 S.t160 S.n9734 0.001
R56877 S.n9734 S.n9731 0.001
R56878 S.t19 S.n8248 0.001
R56879 S.t19 S.n8245 0.001
R56880 S.n8245 S.n8242 0.001
R56881 S.t141 S.n9126 0.001
R56882 S.t141 S.n9129 0.001
R56883 S.t47 S.n7184 0.001
R56884 S.t47 S.n7181 0.001
R56885 S.n7181 S.n7178 0.001
R56886 S.t406 S.n8051 0.001
R56887 S.t406 S.n8054 0.001
R56888 S.t83 S.n6107 0.001
R56889 S.t83 S.n6104 0.001
R56890 S.n6104 S.n6101 0.001
R56891 S.t130 S.n6949 0.001
R56892 S.t130 S.n6952 0.001
R56893 S.t214 S.n5007 0.001
R56894 S.t214 S.n5004 0.001
R56895 S.n5004 S.n5001 0.001
R56896 S.t288 S.n5839 0.001
R56897 S.t288 S.n5842 0.001
R56898 S.t176 S.n3895 0.001
R56899 S.t176 S.n3892 0.001
R56900 S.n3892 S.n3889 0.001
R56901 S.t134 S.n4704 0.001
R56902 S.t134 S.n4707 0.001
R56903 S.t14 S.n2768 0.001
R56904 S.t14 S.n2765 0.001
R56905 S.n2765 S.n2762 0.001
R56906 S.t163 S.n3562 0.001
R56907 S.t163 S.n3565 0.001
R56908 S.t75 S.n1595 0.001
R56909 S.t75 S.n1592 0.001
R56910 S.n1592 S.n1589 0.001
R56911 S.t270 S.n2405 0.001
R56912 S.t270 S.n2408 0.001
R56913 S.t137 S.n574 0.001
R56914 S.t137 S.n571 0.001
R56915 S.n571 S.n568 0.001
R56916 S.t137 S.n557 0.001
R56917 S.t137 S.n554 0.001
R56918 S.n554 S.n551 0.001
R56919 S.t109 S.n220 0.001
R56920 S.t109 S.n217 0.001
R56921 S.n217 S.n214 0.001
R56922 S.t270 S.n2494 0.001
R56923 S.t270 S.n2497 0.001
R56924 S.t130 S.n6501 0.001
R56925 S.t130 S.n6498 0.001
R56926 S.n6498 S.n6495 0.001
R56927 S.t214 S.n4952 0.001
R56928 S.t214 S.n4949 0.001
R56929 S.n4949 S.n4946 0.001
R56930 S.t288 S.n5936 0.001
R56931 S.t288 S.n5939 0.001
R56932 S.t176 S.n3842 0.001
R56933 S.t176 S.n3839 0.001
R56934 S.n3839 S.n3836 0.001
R56935 S.t134 S.n4797 0.001
R56936 S.t134 S.n4800 0.001
R56937 S.t14 S.n2715 0.001
R56938 S.t14 S.n2712 0.001
R56939 S.n2712 S.n2709 0.001
R56940 S.t163 S.n3653 0.001
R56941 S.t163 S.n3656 0.001
R56942 S.t75 S.n1541 0.001
R56943 S.t75 S.n1538 0.001
R56944 S.n1538 S.n1535 0.001
R56945 S.n1086 S.n1081 0.001
R56946 S.t406 S.n7599 0.001
R56947 S.t406 S.n7596 0.001
R56948 S.n7596 S.n7593 0.001
R56949 S.t83 S.n6071 0.001
R56950 S.t83 S.n6068 0.001
R56951 S.n6068 S.n6065 0.001
R56952 S.t130 S.n7014 0.001
R56953 S.t130 S.n7017 0.001
R56954 S.t214 S.n4971 0.001
R56955 S.t214 S.n4968 0.001
R56956 S.n4968 S.n4965 0.001
R56957 S.t288 S.n5904 0.001
R56958 S.t288 S.n5907 0.001
R56959 S.t176 S.n3859 0.001
R56960 S.t176 S.n3856 0.001
R56961 S.n3856 S.n3853 0.001
R56962 S.t134 S.n4765 0.001
R56963 S.t134 S.n4768 0.001
R56964 S.t14 S.n2732 0.001
R56965 S.t14 S.n2729 0.001
R56966 S.n2729 S.n2726 0.001
R56967 S.t163 S.n3622 0.001
R56968 S.t163 S.n3625 0.001
R56969 S.t75 S.n1558 0.001
R56970 S.t75 S.n1555 0.001
R56971 S.n1555 S.n1552 0.001
R56972 S.t270 S.n2464 0.001
R56973 S.t270 S.n2467 0.001
R56974 S.t137 S.n539 0.001
R56975 S.t137 S.n536 0.001
R56976 S.n536 S.n533 0.001
R56977 S.t137 S.n522 0.001
R56978 S.t137 S.n519 0.001
R56979 S.n519 S.n516 0.001
R56980 S.t109 S.n188 0.001
R56981 S.t109 S.n185 0.001
R56982 S.n185 S.n182 0.001
R56983 S.t270 S.n2553 0.001
R56984 S.t270 S.n2556 0.001
R56985 S.t134 S.n4256 0.001
R56986 S.t134 S.n4253 0.001
R56987 S.n4253 S.n4250 0.001
R56988 S.t14 S.n2677 0.001
R56989 S.t14 S.n2674 0.001
R56990 S.n2674 S.n2671 0.001
R56991 S.t163 S.n3717 0.001
R56992 S.t163 S.n3720 0.001
R56993 S.t75 S.n1504 0.001
R56994 S.t75 S.n1501 0.001
R56995 S.n1501 S.n1498 0.001
R56996 S.n1118 S.n1113 0.001
R56997 S.t288 S.n5390 0.001
R56998 S.t288 S.n5387 0.001
R56999 S.n5387 S.n5384 0.001
R57000 S.t176 S.n3823 0.001
R57001 S.t176 S.n3820 0.001
R57002 S.n3820 S.n3817 0.001
R57003 S.t134 S.n4830 0.001
R57004 S.t134 S.n4833 0.001
R57005 S.t14 S.n2696 0.001
R57006 S.t14 S.n2693 0.001
R57007 S.n2693 S.n2690 0.001
R57008 S.t163 S.n3686 0.001
R57009 S.t163 S.n3689 0.001
R57010 S.t75 S.n1521 0.001
R57011 S.t75 S.n1518 0.001
R57012 S.n1518 S.n1515 0.001
R57013 S.t270 S.n2523 0.001
R57014 S.t270 S.n2526 0.001
R57015 S.t137 S.n504 0.001
R57016 S.t137 S.n501 0.001
R57017 S.n501 S.n498 0.001
R57018 S.t137 S.n487 0.001
R57019 S.t137 S.n484 0.001
R57020 S.n484 S.n481 0.001
R57021 S.t109 S.n156 0.001
R57022 S.t109 S.n153 0.001
R57023 S.n153 S.n150 0.001
R57024 S.t270 S.n1960 0.001
R57025 S.t270 S.n1957 0.001
R57026 S.n1957 S.n1954 0.001
R57027 S.n1156 S.n1151 0.001
R57028 S.t163 S.n3120 0.001
R57029 S.t163 S.n3117 0.001
R57030 S.n3117 S.n3114 0.001
R57031 S.t75 S.n1484 0.001
R57032 S.t75 S.n1481 0.001
R57033 S.n1481 S.n1478 0.001
R57034 S.t270 S.n2586 0.001
R57035 S.t270 S.n2589 0.001
R57036 S.t137 S.n469 0.001
R57037 S.t137 S.n466 0.001
R57038 S.n466 S.n463 0.001
R57039 S.t137 S.n453 0.001
R57040 S.t137 S.n450 0.001
R57041 S.n450 S.n447 0.001
R57042 S.t109 S.n945 0.001
R57043 S.t109 S.n948 0.001
R57044 S.n22310 S.n22307 0.001
R57045 S.t9 S.n22313 0.001
R57046 S.n21971 S.t105 0.001
R57047 S.n21980 S.n21973 0.001
R57048 S.t88 S.n22768 0.001
R57049 S.t88 S.n22771 0.001
R57050 S.t100 S.n21334 0.001
R57051 S.t100 S.n21331 0.001
R57052 S.n21331 S.n21328 0.001
R57053 S.t9 S.n22339 0.001
R57054 S.n22333 S.n22332 0.001
R57055 S.t9 S.n22310 0.001
R57056 S.n22768 S.n22765 0.001
R57057 S.n21980 S.n21971 0.001
R57058 S.n1422 S.t158 0.001
R57059 S.n890 S.n877 0.001
R57060 S.n1988 S.n1985 0.001
R57061 S.n3149 S.n3146 0.001
R57062 S.n4286 S.n4283 0.001
R57063 S.n5420 S.n5417 0.001
R57064 S.n6531 S.n6528 0.001
R57065 S.n7629 S.n7626 0.001
R57066 S.n8704 S.n8701 0.001
R57067 S.n9767 S.n9764 0.001
R57068 S.n10807 S.n10804 0.001
R57069 S.n11835 S.n11832 0.001
R57070 S.n12840 S.n12837 0.001
R57071 S.n13833 S.n13830 0.001
R57072 S.n14803 S.n14800 0.001
R57073 S.n15761 S.n15758 0.001
R57074 S.n16696 S.n16693 0.001
R57075 S.n17619 S.n17616 0.001
R57076 S.n18519 S.n18516 0.001
R57077 S.n19406 S.n19403 0.001
R57078 S.n20274 S.n20271 0.001
R57079 S.n21245 S.n21242 0.001
R57080 S.n20298 S.n20295 0.001
R57081 S.n19426 S.n19423 0.001
R57082 S.n18539 S.n18536 0.001
R57083 S.n17639 S.n17636 0.001
R57084 S.n16716 S.n16713 0.001
R57085 S.n15781 S.n15778 0.001
R57086 S.n14823 S.n14820 0.001
R57087 S.n13853 S.n13850 0.001
R57088 S.n12860 S.n12857 0.001
R57089 S.n11855 S.n11852 0.001
R57090 S.n10827 S.n10824 0.001
R57091 S.n9787 S.n9784 0.001
R57092 S.n8724 S.n8721 0.001
R57093 S.n7649 S.n7646 0.001
R57094 S.n6551 S.n6548 0.001
R57095 S.n5441 S.n5438 0.001
R57096 S.n4306 S.n4303 0.001
R57097 S.n3169 S.n3166 0.001
R57098 S.n2015 S.n2012 0.001
R57099 S.n20427 S.n20424 0.001
R57100 S.n20333 S.n20330 0.001
R57101 S.n19461 S.n19458 0.001
R57102 S.n18571 S.n18568 0.001
R57103 S.n17671 S.n17668 0.001
R57104 S.n16748 S.n16745 0.001
R57105 S.n15813 S.n15810 0.001
R57106 S.n14855 S.n14852 0.001
R57107 S.n13885 S.n13882 0.001
R57108 S.n12892 S.n12889 0.001
R57109 S.n11887 S.n11884 0.001
R57110 S.n10859 S.n10856 0.001
R57111 S.n9819 S.n9816 0.001
R57112 S.n8756 S.n8753 0.001
R57113 S.n7681 S.n7678 0.001
R57114 S.n6583 S.n6580 0.001
R57115 S.n5473 S.n5470 0.001
R57116 S.n4338 S.n4335 0.001
R57117 S.n3201 S.n3198 0.001
R57118 S.n2048 S.n2045 0.001
R57119 S.n1337 S.n1328 0.001
R57120 S.n823 S.n815 0.001
R57121 S.n2082 S.n2079 0.001
R57122 S.n3233 S.n3230 0.001
R57123 S.n4370 S.n4367 0.001
R57124 S.n5505 S.n5502 0.001
R57125 S.n6615 S.n6612 0.001
R57126 S.n7713 S.n7710 0.001
R57127 S.n8788 S.n8785 0.001
R57128 S.n9851 S.n9848 0.001
R57129 S.n10891 S.n10888 0.001
R57130 S.n11919 S.n11916 0.001
R57131 S.n12924 S.n12921 0.001
R57132 S.n13917 S.n13914 0.001
R57133 S.n14887 S.n14884 0.001
R57134 S.n15845 S.n15842 0.001
R57135 S.n16780 S.n16777 0.001
R57136 S.n17703 S.n17700 0.001
R57137 S.n18603 S.n18600 0.001
R57138 S.n19493 S.n19490 0.001
R57139 S.n18636 S.n18633 0.001
R57140 S.n17736 S.n17733 0.001
R57141 S.n16809 S.n16806 0.001
R57142 S.n15874 S.n15871 0.001
R57143 S.n14916 S.n14913 0.001
R57144 S.n13946 S.n13943 0.001
R57145 S.n12953 S.n12950 0.001
R57146 S.n11948 S.n11945 0.001
R57147 S.n10920 S.n10917 0.001
R57148 S.n9880 S.n9877 0.001
R57149 S.n8817 S.n8814 0.001
R57150 S.n7742 S.n7739 0.001
R57151 S.n6644 S.n6641 0.001
R57152 S.n5534 S.n5531 0.001
R57153 S.n4399 S.n4396 0.001
R57154 S.n3262 S.n3259 0.001
R57155 S.n2110 S.n2107 0.001
R57156 S.n24 S.n16 0.001
R57157 S.n2140 S.n2137 0.001
R57158 S.n3293 S.n3290 0.001
R57159 S.n4431 S.n4428 0.001
R57160 S.n5566 S.n5563 0.001
R57161 S.n6676 S.n6673 0.001
R57162 S.n7774 S.n7771 0.001
R57163 S.n8849 S.n8846 0.001
R57164 S.n9912 S.n9909 0.001
R57165 S.n10952 S.n10949 0.001
R57166 S.n11980 S.n11977 0.001
R57167 S.n12985 S.n12982 0.001
R57168 S.n13978 S.n13975 0.001
R57169 S.n14948 S.n14945 0.001
R57170 S.n15906 S.n15903 0.001
R57171 S.n16841 S.n16838 0.001
R57172 S.n17768 S.n17765 0.001
R57173 S.n16874 S.n16871 0.001
R57174 S.n15939 S.n15936 0.001
R57175 S.n14977 S.n14974 0.001
R57176 S.n14007 S.n14004 0.001
R57177 S.n13014 S.n13011 0.001
R57178 S.n12009 S.n12006 0.001
R57179 S.n10981 S.n10978 0.001
R57180 S.n9941 S.n9938 0.001
R57181 S.n8878 S.n8875 0.001
R57182 S.n7803 S.n7800 0.001
R57183 S.n6705 S.n6702 0.001
R57184 S.n5595 S.n5592 0.001
R57185 S.n4460 S.n4457 0.001
R57186 S.n3322 S.n3319 0.001
R57187 S.n2169 S.n2166 0.001
R57188 S.n71 S.n63 0.001
R57189 S.n2199 S.n2196 0.001
R57190 S.n3353 S.n3350 0.001
R57191 S.n4492 S.n4489 0.001
R57192 S.n5627 S.n5624 0.001
R57193 S.n6737 S.n6734 0.001
R57194 S.n7835 S.n7832 0.001
R57195 S.n8910 S.n8907 0.001
R57196 S.n9973 S.n9970 0.001
R57197 S.n11013 S.n11010 0.001
R57198 S.n12041 S.n12038 0.001
R57199 S.n13046 S.n13043 0.001
R57200 S.n14039 S.n14036 0.001
R57201 S.n15009 S.n15006 0.001
R57202 S.n15971 S.n15968 0.001
R57203 S.n15042 S.n15039 0.001
R57204 S.n14072 S.n14069 0.001
R57205 S.n13075 S.n13072 0.001
R57206 S.n12070 S.n12067 0.001
R57207 S.n11042 S.n11039 0.001
R57208 S.n10002 S.n9999 0.001
R57209 S.n8939 S.n8936 0.001
R57210 S.n7864 S.n7861 0.001
R57211 S.n6766 S.n6763 0.001
R57212 S.n5656 S.n5653 0.001
R57213 S.n4521 S.n4518 0.001
R57214 S.n3382 S.n3379 0.001
R57215 S.n2228 S.n2225 0.001
R57216 S.n103 S.n95 0.001
R57217 S.n2258 S.n2255 0.001
R57218 S.n3413 S.n3410 0.001
R57219 S.n4553 S.n4550 0.001
R57220 S.n5688 S.n5685 0.001
R57221 S.n6798 S.n6795 0.001
R57222 S.n7896 S.n7893 0.001
R57223 S.n8971 S.n8968 0.001
R57224 S.n10034 S.n10031 0.001
R57225 S.n11074 S.n11071 0.001
R57226 S.n12102 S.n12099 0.001
R57227 S.n13107 S.n13104 0.001
R57228 S.n14104 S.n14101 0.001
R57229 S.n13140 S.n13137 0.001
R57230 S.n12135 S.n12132 0.001
R57231 S.n11103 S.n11100 0.001
R57232 S.n10063 S.n10060 0.001
R57233 S.n9000 S.n8997 0.001
R57234 S.n7925 S.n7922 0.001
R57235 S.n6827 S.n6824 0.001
R57236 S.n5717 S.n5714 0.001
R57237 S.n4582 S.n4579 0.001
R57238 S.n3442 S.n3439 0.001
R57239 S.n2287 S.n2284 0.001
R57240 S.n990 S.n982 0.001
R57241 S.n2317 S.n2314 0.001
R57242 S.n3473 S.n3470 0.001
R57243 S.n4614 S.n4611 0.001
R57244 S.n5749 S.n5746 0.001
R57245 S.n6859 S.n6856 0.001
R57246 S.n7957 S.n7954 0.001
R57247 S.n9032 S.n9029 0.001
R57248 S.n10095 S.n10092 0.001
R57249 S.n11135 S.n11132 0.001
R57250 S.n12167 S.n12164 0.001
R57251 S.n11168 S.n11165 0.001
R57252 S.n10128 S.n10125 0.001
R57253 S.n9061 S.n9058 0.001
R57254 S.n7986 S.n7983 0.001
R57255 S.n6888 S.n6885 0.001
R57256 S.n5778 S.n5775 0.001
R57257 S.n4643 S.n4640 0.001
R57258 S.n3502 S.n3499 0.001
R57259 S.n2346 S.n2343 0.001
R57260 S.n1022 S.n1014 0.001
R57261 S.n2376 S.n2373 0.001
R57262 S.n3533 S.n3530 0.001
R57263 S.n4675 S.n4672 0.001
R57264 S.n5810 S.n5807 0.001
R57265 S.n6920 S.n6917 0.001
R57266 S.n8018 S.n8015 0.001
R57267 S.n9093 S.n9090 0.001
R57268 S.n10160 S.n10157 0.001
R57269 S.n9126 S.n9123 0.001
R57270 S.n8051 S.n8048 0.001
R57271 S.n6949 S.n6946 0.001
R57272 S.n5839 S.n5836 0.001
R57273 S.n4704 S.n4701 0.001
R57274 S.n3562 S.n3559 0.001
R57275 S.n2405 S.n2402 0.001
R57276 S.n1054 S.n1046 0.001
R57277 S.n252 S.n249 0.001
R57278 S.n2435 S.n2432 0.001
R57279 S.n3593 S.n3590 0.001
R57280 S.n4736 S.n4733 0.001
R57281 S.n5871 S.n5868 0.001
R57282 S.n6981 S.n6978 0.001
R57283 S.n8083 S.n8080 0.001
R57284 S.n7014 S.n7011 0.001
R57285 S.n5904 S.n5901 0.001
R57286 S.n4765 S.n4762 0.001
R57287 S.n3622 S.n3619 0.001
R57288 S.n2464 S.n2461 0.001
R57289 S.n1086 S.n1078 0.001
R57290 S.n2494 S.n2491 0.001
R57291 S.n3653 S.n3650 0.001
R57292 S.n4797 S.n4794 0.001
R57293 S.n5936 S.n5933 0.001
R57294 S.n4830 S.n4827 0.001
R57295 S.n3686 S.n3683 0.001
R57296 S.n2523 S.n2520 0.001
R57297 S.n1118 S.n1110 0.001
R57298 S.n2553 S.n2550 0.001
R57299 S.n3717 S.n3714 0.001
R57300 S.n2586 S.n2583 0.001
R57301 S.n1156 S.n1148 0.001
R57302 S.n945 S.n942 0.001
R57303 S.n977 S.n974 0.001
R57304 S.n22354 S.n22351 0.001
R57305 S.n21348 S.n21345 0.001
R57306 S.n21264 S.n21261 0.001
R57307 S.n20835 S.n20827 0.001
R57308 S.n20848 S.n20845 0.001
R57309 S.n20200 S.n20192 0.001
R57310 S.n19330 S.n19322 0.001
R57311 S.n18448 S.n18440 0.001
R57312 S.n17543 S.n17535 0.001
R57313 S.n16625 S.n16617 0.001
R57314 S.n15685 S.n15677 0.001
R57315 S.n14732 S.n14724 0.001
R57316 S.n13757 S.n13749 0.001
R57317 S.n12769 S.n12761 0.001
R57318 S.n11759 S.n11751 0.001
R57319 S.n10736 S.n10728 0.001
R57320 S.n9691 S.n9683 0.001
R57321 S.n8633 S.n8625 0.001
R57322 S.n7553 S.n7545 0.001
R57323 S.n6460 S.n6452 0.001
R57324 S.n5344 S.n5336 0.001
R57325 S.n4215 S.n4207 0.001
R57326 S.n3074 S.n3066 0.001
R57327 S.n1885 S.n1882 0.001
R57328 S.n809 S.n806 0.001
R57329 S.n2597 S.n2596 0.001
R57330 S.n22371 S.n22368 0.001
R57331 S.n21654 S.n21650 0.001
R57332 S.n21659 S.n21656 0.001
R57333 S.n20510 S.n20507 0.001
R57334 S.n20864 S.n20861 0.001
R57335 S.n19899 S.n19896 0.001
R57336 S.n19045 S.n19042 0.001
R57337 S.n18179 S.n18176 0.001
R57338 S.n17290 S.n17287 0.001
R57339 S.n16388 S.n16385 0.001
R57340 S.n15464 S.n15461 0.001
R57341 S.n14527 S.n14524 0.001
R57342 S.n13568 S.n13565 0.001
R57343 S.n12596 S.n12593 0.001
R57344 S.n11602 S.n11599 0.001
R57345 S.n10595 S.n10592 0.001
R57346 S.n9566 S.n9563 0.001
R57347 S.n8524 S.n8521 0.001
R57348 S.n7460 S.n7457 0.001
R57349 S.n6383 S.n6380 0.001
R57350 S.n5283 S.n5280 0.001
R57351 S.n4170 S.n4167 0.001
R57352 S.n3044 S.n3041 0.001
R57353 S.n1899 S.n1891 0.001
R57354 S.n3728 S.n3727 0.001
R57355 S.n22672 S.n22668 0.001
R57356 S.n21685 S.n21681 0.001
R57357 S.n21690 S.n21687 0.001
R57358 S.n20525 S.n20522 0.001
R57359 S.n20880 S.n20877 0.001
R57360 S.n19914 S.n19911 0.001
R57361 S.n19060 S.n19057 0.001
R57362 S.n18194 S.n18191 0.001
R57363 S.n17305 S.n17302 0.001
R57364 S.n16403 S.n16400 0.001
R57365 S.n15479 S.n15476 0.001
R57366 S.n14542 S.n14539 0.001
R57367 S.n13583 S.n13580 0.001
R57368 S.n12611 S.n12608 0.001
R57369 S.n11617 S.n11614 0.001
R57370 S.n10610 S.n10607 0.001
R57371 S.n9581 S.n9578 0.001
R57372 S.n8539 S.n8536 0.001
R57373 S.n7475 S.n7472 0.001
R57374 S.n6398 S.n6395 0.001
R57375 S.n5298 S.n5295 0.001
R57376 S.n4185 S.n4182 0.001
R57377 S.n3060 S.n3057 0.001
R57378 S.n4841 S.n4840 0.001
R57379 S.n4201 S.n4198 0.001
R57380 S.n5314 S.n5311 0.001
R57381 S.n6414 S.n6411 0.001
R57382 S.n7491 S.n7488 0.001
R57383 S.n8555 S.n8552 0.001
R57384 S.n9232 S.n9229 0.001
R57385 S.n9597 S.n9594 0.001
R57386 S.n10626 S.n10623 0.001
R57387 S.n11633 S.n11630 0.001
R57388 S.n12627 S.n12624 0.001
R57389 S.n13599 S.n13596 0.001
R57390 S.n14558 S.n14555 0.001
R57391 S.n15495 S.n15492 0.001
R57392 S.n16419 S.n16416 0.001
R57393 S.n17321 S.n17318 0.001
R57394 S.n18210 S.n18207 0.001
R57395 S.n19076 S.n19073 0.001
R57396 S.n19930 S.n19927 0.001
R57397 S.n20895 S.n20892 0.001
R57398 S.n20541 S.n20538 0.001
R57399 S.n21705 S.n21702 0.001
R57400 S.n21364 S.n21361 0.001
R57401 S.n22387 S.n22384 0.001
R57402 S.n5947 S.n5946 0.001
R57403 S.n5330 S.n5327 0.001
R57404 S.n6430 S.n6427 0.001
R57405 S.n7507 S.n7504 0.001
R57406 S.n8571 S.n8568 0.001
R57407 S.n9613 S.n9610 0.001
R57408 S.n10642 S.n10639 0.001
R57409 S.n11649 S.n11646 0.001
R57410 S.n12643 S.n12640 0.001
R57411 S.n13615 S.n13612 0.001
R57412 S.n14574 S.n14571 0.001
R57413 S.n15511 S.n15508 0.001
R57414 S.n16435 S.n16432 0.001
R57415 S.n17337 S.n17334 0.001
R57416 S.n18226 S.n18223 0.001
R57417 S.n19092 S.n19089 0.001
R57418 S.n19946 S.n19943 0.001
R57419 S.n20910 S.n20907 0.001
R57420 S.n20557 S.n20554 0.001
R57421 S.n21720 S.n21717 0.001
R57422 S.n21380 S.n21377 0.001
R57423 S.n22403 S.n22400 0.001
R57424 S.n7025 S.n7024 0.001
R57425 S.n6446 S.n6443 0.001
R57426 S.n7523 S.n7520 0.001
R57427 S.n8587 S.n8584 0.001
R57428 S.n9629 S.n9626 0.001
R57429 S.n10658 S.n10655 0.001
R57430 S.n11665 S.n11662 0.001
R57431 S.n12659 S.n12656 0.001
R57432 S.n13631 S.n13628 0.001
R57433 S.n14590 S.n14587 0.001
R57434 S.n15527 S.n15524 0.001
R57435 S.n16451 S.n16448 0.001
R57436 S.n17353 S.n17350 0.001
R57437 S.n18242 S.n18239 0.001
R57438 S.n19108 S.n19105 0.001
R57439 S.n19962 S.n19959 0.001
R57440 S.n20925 S.n20922 0.001
R57441 S.n20573 S.n20570 0.001
R57442 S.n21735 S.n21732 0.001
R57443 S.n21396 S.n21393 0.001
R57444 S.n22419 S.n22416 0.001
R57445 S.n8094 S.n8093 0.001
R57446 S.n7539 S.n7536 0.001
R57447 S.n8603 S.n8600 0.001
R57448 S.n9645 S.n9642 0.001
R57449 S.n10674 S.n10671 0.001
R57450 S.n11681 S.n11678 0.001
R57451 S.n12675 S.n12672 0.001
R57452 S.n13647 S.n13644 0.001
R57453 S.n14606 S.n14603 0.001
R57454 S.n15543 S.n15540 0.001
R57455 S.n16467 S.n16464 0.001
R57456 S.n17369 S.n17366 0.001
R57457 S.n18258 S.n18255 0.001
R57458 S.n19124 S.n19121 0.001
R57459 S.n19978 S.n19975 0.001
R57460 S.n20940 S.n20937 0.001
R57461 S.n20589 S.n20586 0.001
R57462 S.n21750 S.n21747 0.001
R57463 S.n21412 S.n21409 0.001
R57464 S.n22435 S.n22432 0.001
R57465 S.n9137 S.n9136 0.001
R57466 S.n8619 S.n8616 0.001
R57467 S.n9661 S.n9658 0.001
R57468 S.n10690 S.n10687 0.001
R57469 S.n11697 S.n11694 0.001
R57470 S.n12691 S.n12688 0.001
R57471 S.n13663 S.n13660 0.001
R57472 S.n14622 S.n14619 0.001
R57473 S.n15559 S.n15556 0.001
R57474 S.n16483 S.n16480 0.001
R57475 S.n17385 S.n17382 0.001
R57476 S.n18274 S.n18271 0.001
R57477 S.n19140 S.n19137 0.001
R57478 S.n19994 S.n19991 0.001
R57479 S.n20955 S.n20952 0.001
R57480 S.n20605 S.n20602 0.001
R57481 S.n21765 S.n21762 0.001
R57482 S.n21428 S.n21425 0.001
R57483 S.n22451 S.n22448 0.001
R57484 S.n10171 S.n10170 0.001
R57485 S.n9677 S.n9674 0.001
R57486 S.n10706 S.n10703 0.001
R57487 S.n11713 S.n11710 0.001
R57488 S.n12707 S.n12704 0.001
R57489 S.n13679 S.n13676 0.001
R57490 S.n14638 S.n14635 0.001
R57491 S.n15575 S.n15572 0.001
R57492 S.n16499 S.n16496 0.001
R57493 S.n17401 S.n17398 0.001
R57494 S.n18290 S.n18287 0.001
R57495 S.n19156 S.n19153 0.001
R57496 S.n20010 S.n20007 0.001
R57497 S.n20970 S.n20967 0.001
R57498 S.n20621 S.n20618 0.001
R57499 S.n21780 S.n21777 0.001
R57500 S.n21444 S.n21441 0.001
R57501 S.n22467 S.n22464 0.001
R57502 S.n11179 S.n11178 0.001
R57503 S.n10722 S.n10719 0.001
R57504 S.n11729 S.n11726 0.001
R57505 S.n12723 S.n12720 0.001
R57506 S.n13695 S.n13692 0.001
R57507 S.n14654 S.n14651 0.001
R57508 S.n15591 S.n15588 0.001
R57509 S.n16515 S.n16512 0.001
R57510 S.n17417 S.n17414 0.001
R57511 S.n18306 S.n18303 0.001
R57512 S.n19172 S.n19169 0.001
R57513 S.n20026 S.n20023 0.001
R57514 S.n20985 S.n20982 0.001
R57515 S.n20637 S.n20634 0.001
R57516 S.n21795 S.n21792 0.001
R57517 S.n21460 S.n21457 0.001
R57518 S.n22483 S.n22480 0.001
R57519 S.n12178 S.n12177 0.001
R57520 S.n11745 S.n11742 0.001
R57521 S.n12739 S.n12736 0.001
R57522 S.n13711 S.n13708 0.001
R57523 S.n14670 S.n14667 0.001
R57524 S.n15607 S.n15604 0.001
R57525 S.n16531 S.n16528 0.001
R57526 S.n17433 S.n17430 0.001
R57527 S.n18322 S.n18319 0.001
R57528 S.n19188 S.n19185 0.001
R57529 S.n20042 S.n20039 0.001
R57530 S.n21000 S.n20997 0.001
R57531 S.n20653 S.n20650 0.001
R57532 S.n21810 S.n21807 0.001
R57533 S.n21476 S.n21473 0.001
R57534 S.n22499 S.n22496 0.001
R57535 S.n13151 S.n13150 0.001
R57536 S.n12755 S.n12752 0.001
R57537 S.n13727 S.n13724 0.001
R57538 S.n14686 S.n14683 0.001
R57539 S.n15623 S.n15620 0.001
R57540 S.n16547 S.n16544 0.001
R57541 S.n17449 S.n17446 0.001
R57542 S.n18338 S.n18335 0.001
R57543 S.n19204 S.n19201 0.001
R57544 S.n20058 S.n20055 0.001
R57545 S.n21015 S.n21012 0.001
R57546 S.n20669 S.n20666 0.001
R57547 S.n21825 S.n21822 0.001
R57548 S.n21492 S.n21489 0.001
R57549 S.n22515 S.n22512 0.001
R57550 S.n14115 S.n14114 0.001
R57551 S.n13743 S.n13740 0.001
R57552 S.n14702 S.n14699 0.001
R57553 S.n15639 S.n15636 0.001
R57554 S.n16563 S.n16560 0.001
R57555 S.n17465 S.n17462 0.001
R57556 S.n18354 S.n18351 0.001
R57557 S.n19220 S.n19217 0.001
R57558 S.n20074 S.n20071 0.001
R57559 S.n21030 S.n21027 0.001
R57560 S.n20685 S.n20682 0.001
R57561 S.n21840 S.n21837 0.001
R57562 S.n21508 S.n21505 0.001
R57563 S.n22531 S.n22528 0.001
R57564 S.n15053 S.n15052 0.001
R57565 S.n14718 S.n14715 0.001
R57566 S.n15655 S.n15652 0.001
R57567 S.n16579 S.n16576 0.001
R57568 S.n17481 S.n17478 0.001
R57569 S.n18370 S.n18367 0.001
R57570 S.n19236 S.n19233 0.001
R57571 S.n20090 S.n20087 0.001
R57572 S.n21045 S.n21042 0.001
R57573 S.n20701 S.n20698 0.001
R57574 S.n21855 S.n21852 0.001
R57575 S.n21524 S.n21521 0.001
R57576 S.n22547 S.n22544 0.001
R57577 S.n15982 S.n15981 0.001
R57578 S.n15671 S.n15668 0.001
R57579 S.n16595 S.n16592 0.001
R57580 S.n17497 S.n17494 0.001
R57581 S.n18386 S.n18383 0.001
R57582 S.n19252 S.n19249 0.001
R57583 S.n20106 S.n20103 0.001
R57584 S.n21060 S.n21057 0.001
R57585 S.n20717 S.n20714 0.001
R57586 S.n21870 S.n21867 0.001
R57587 S.n21540 S.n21537 0.001
R57588 S.n22563 S.n22560 0.001
R57589 S.n16885 S.n16884 0.001
R57590 S.n16611 S.n16608 0.001
R57591 S.n17513 S.n17510 0.001
R57592 S.n18402 S.n18399 0.001
R57593 S.n19268 S.n19265 0.001
R57594 S.n20122 S.n20119 0.001
R57595 S.n21075 S.n21072 0.001
R57596 S.n20733 S.n20730 0.001
R57597 S.n21885 S.n21882 0.001
R57598 S.n21556 S.n21553 0.001
R57599 S.n22579 S.n22576 0.001
R57600 S.n17779 S.n17778 0.001
R57601 S.n17529 S.n17526 0.001
R57602 S.n18418 S.n18415 0.001
R57603 S.n19284 S.n19281 0.001
R57604 S.n20138 S.n20135 0.001
R57605 S.n21090 S.n21087 0.001
R57606 S.n20749 S.n20746 0.001
R57607 S.n21900 S.n21897 0.001
R57608 S.n21572 S.n21569 0.001
R57609 S.n22595 S.n22592 0.001
R57610 S.n18647 S.n18646 0.001
R57611 S.n18434 S.n18431 0.001
R57612 S.n19300 S.n19297 0.001
R57613 S.n20154 S.n20151 0.001
R57614 S.n21105 S.n21102 0.001
R57615 S.n20765 S.n20762 0.001
R57616 S.n21915 S.n21912 0.001
R57617 S.n21588 S.n21585 0.001
R57618 S.n22611 S.n22608 0.001
R57619 S.n19504 S.n19503 0.001
R57620 S.n19316 S.n19313 0.001
R57621 S.n20170 S.n20167 0.001
R57622 S.n21120 S.n21117 0.001
R57623 S.n20781 S.n20778 0.001
R57624 S.n21930 S.n21927 0.001
R57625 S.n21604 S.n21601 0.001
R57626 S.n22627 S.n22624 0.001
R57627 S.n20344 S.n20343 0.001
R57628 S.n20186 S.n20183 0.001
R57629 S.n21136 S.n21133 0.001
R57630 S.n20797 S.n20794 0.001
R57631 S.n21945 S.n21942 0.001
R57632 S.n21620 S.n21617 0.001
R57633 S.n22643 S.n22640 0.001
R57634 S.n21172 S.n21142 0.001
R57635 S.n20821 S.n20818 0.001
R57636 S.n21965 S.n21962 0.001
R57637 S.n21641 S.n21638 0.001
R57638 S.n22659 S.n22656 0.001
R57639 S.n22979 S.n22978 0.001
R57640 S.n22978 S.n22971 0.001
R57641 S.n971 S.n970 0.001
R57642 S.n1911 S.n1910 0.001
R57643 S.n2612 S.n2611 0.001
R57644 S.n3743 S.n3742 0.001
R57645 S.n4856 S.n4855 0.001
R57646 S.n5961 S.n5960 0.001
R57647 S.n7039 S.n7038 0.001
R57648 S.n8108 S.n8107 0.001
R57649 S.n9151 S.n9150 0.001
R57650 S.n10185 S.n10184 0.001
R57651 S.n11193 S.n11192 0.001
R57652 S.n12192 S.n12191 0.001
R57653 S.n13165 S.n13164 0.001
R57654 S.n14129 S.n14128 0.001
R57655 S.n15067 S.n15066 0.001
R57656 S.n15996 S.n15995 0.001
R57657 S.n16899 S.n16898 0.001
R57658 S.n17793 S.n17792 0.001
R57659 S.n18661 S.n18660 0.001
R57660 S.n19518 S.n19517 0.001
R57661 S.n21168 S.n21167 0.001
R57662 S.n21186 S.n21185 0.001
R57663 S.n22784 S.n22783 0.001
R57664 S.n22280 S.n22279 0.001
R57665 S.n22799 S.n22798 0.001
R57666 S.n1177 S.n1176 0.001
R57667 S.n1180 S.n1179 0.001
R57668 S.n22798 S.n22797 0.001
R57669 S.n970 S.n969 0.001
R57670 S.n1910 S.n1909 0.001
R57671 S.n2611 S.n2610 0.001
R57672 S.n3742 S.n3741 0.001
R57673 S.n4855 S.n4854 0.001
R57674 S.n5960 S.n5959 0.001
R57675 S.n7038 S.n7037 0.001
R57676 S.n8107 S.n8106 0.001
R57677 S.n9150 S.n9149 0.001
R57678 S.n10184 S.n10183 0.001
R57679 S.n11192 S.n11191 0.001
R57680 S.n12191 S.n12190 0.001
R57681 S.n13164 S.n13163 0.001
R57682 S.n14128 S.n14127 0.001
R57683 S.n15066 S.n15065 0.001
R57684 S.n15995 S.n15994 0.001
R57685 S.n16898 S.n16897 0.001
R57686 S.n17792 S.n17791 0.001
R57687 S.n18660 S.n18659 0.001
R57688 S.n19517 S.n19516 0.001
R57689 S.n21167 S.n21166 0.001
R57690 S.n21185 S.n21184 0.001
R57691 S.n22789 S.n22787 0.001
R57692 S.n21187 S.n21177 0.001
R57693 S.n972 S.n962 0.001
R57694 S.n1912 S.n1903 0.001
R57695 S.n2613 S.n2603 0.001
R57696 S.n3744 S.n3734 0.001
R57697 S.n4857 S.n4847 0.001
R57698 S.n5962 S.n5952 0.001
R57699 S.n7040 S.n7030 0.001
R57700 S.n8109 S.n8099 0.001
R57701 S.n9152 S.n9142 0.001
R57702 S.n10186 S.n10176 0.001
R57703 S.n11194 S.n11184 0.001
R57704 S.n12193 S.n12183 0.001
R57705 S.n13166 S.n13156 0.001
R57706 S.n14130 S.n14120 0.001
R57707 S.n15068 S.n15058 0.001
R57708 S.n15997 S.n15987 0.001
R57709 S.n16900 S.n16890 0.001
R57710 S.n17794 S.n17784 0.001
R57711 S.n18662 S.n18652 0.001
R57712 S.n19519 S.n19509 0.001
R57713 S.n21169 S.n21159 0.001
R57714 S.n22802 S.n22801 0.001
R57715 S.n22783 S.n22782 0.001
R57716 S.n22980 S.n22979 0.001
R57717 S.n22971 S.n22970 0.001
R57718 S.n22332 S.n22328 0.001
R57719 PW PW.n0 2.027
C0 S D 8331.87fF
C1 G D 3947.35fF
C2 S G 5238.35fF
.ends

