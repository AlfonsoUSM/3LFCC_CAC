**.subckt prelayout_cap_pmos
VG VP GND PULSE(0 {VGS} 20n 0 0 100n 120n)
.save i(vg)
VSS VSS GND 0
.save i(vss)
R1 G VP 100 m=1
VG1 VP2 GND {VGS}
.save i(vg1)
XM1 VSS G VP2 VP2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4.38 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4512 m=4512
**** begin user architecture code


.param VGS = 5
.option temp=70
.lib /foss/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice tt

.control
compose voltage values (2.5) 5
foreach volt $&voltage
alterparam VGS=$volt
reset
save v(G)
tran 50f 120n
wrdata SPICE_files/PMOS/PRELAYOUT_CAP/PMOS_cap_calc_PRELAYOUT.txt v(G)
set appendwrite
end

.endc



**** end user architecture code
**.ends
.GLOBAL GND
.end
.control
quit
.endc