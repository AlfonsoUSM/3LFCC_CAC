* NGSPICE file created from nmos_24x24_flat.ext - technology: sky130A

.subckt nmos_24x24_flat
X0 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=1.53148e+15p pd=1.0396e+10u as=0p ps=0u w=4.38e+06u l=500000u
X1 S.t1141 G D S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X2 S.t1140 G D S.t168 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X3 D G S.t1139 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X4 D G S.t1138 S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X5 S.t1137 G D S.t48 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X6 S.t1136 G D S.t48 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X7 D G S.t1135 S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X8 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X9 S.t1133 G D S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X10 S.t1132 G D S.t164 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X11 D G S.t1131 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X12 S.t1130 G D S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X13 D G S.t1129 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X14 S.t1128 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X15 D G S.t1127 S.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X16 D G S.t1126 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X17 D G S.t1125 S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X18 S.t1124 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X19 D G S.t1123 S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X20 S.t1122 G D S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X21 D G S.t1121 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X22 D G S.t1120 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X23 S.t1119 G D S.t162 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X24 S.t1118 G D S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X25 D G S.t1117 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X26 S.t1116 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X27 S.t1115 G D S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X28 D G S.t1114 S.t164 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X29 D G S.t1113 S.t162 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X30 D G S.t1112 S.t140 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X31 D G S.t1111 S.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X32 S.t1110 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X33 D G S.t1109 S.t151 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X34 S.t1108 G D S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X35 S.t1107 G D S.t164 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X36 D G S.t1106 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X37 S.t1105 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X38 D G S.t1104 S.t151 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X39 S.t1103 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X40 D G S.t1102 S.t168 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X41 S.t1101 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X42 S.t1100 G D S.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X43 S.t1099 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X44 S.t1098 G D S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X45 S.t1097 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X46 D G S.t1096 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X47 D G S.t1095 S.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X48 D G S.t1094 S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X49 S.t1093 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X50 S.t1092 G D S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X51 D G S.t1091 S.t154 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X52 S.t1090 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X53 D G S.t1089 S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X54 S.t1088 G D S.t140 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X55 S.t1087 G D S.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X56 S.t1086 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X57 S.t1085 G D S.t95 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X58 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X59 D G S.t1083 S.t154 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X60 S.t1082 G D S.t135 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X61 S.t1081 G D S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X62 D G S.t1080 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X63 D G S.t1079 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X64 D G S.t1078 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X65 D G S.t1077 S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X66 S.t1076 G D S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X67 S.t1075 G D S.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X68 S.t1074 G D S.t127 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X69 S.t1073 G D S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X70 S.t1072 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X71 D G S.t1071 S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X72 D G S.t1070 S.t135 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X73 D G S.t1069 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X74 D G S.t1068 S.t162 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X75 S.t1067 G D S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X76 S.t1066 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X77 D G S.t1065 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X78 S.t1064 G D S.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X79 D G S.t1063 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X80 S.t1062 G D S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X81 S.t1061 G D S.t151 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X82 S.t1060 G D S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X83 D G S.t1059 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X84 D G S.t1058 S.t164 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X85 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X86 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X87 S.t1055 G D S.t168 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X88 S.t1054 G D S.t107 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X89 D G S.t1053 S.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X90 D G S.t1052 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X91 D G S.t1051 S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X92 S.t1050 G D S.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X93 D G S.t1049 S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X94 D G S.t1048 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X95 S.t1047 G D S.t95 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X96 D G S.t1046 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X97 S.t1045 G D S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X98 S.t1044 G D S.t154 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X99 D G S.t1043 S.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X100 D G S.t1042 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X101 D G S.t1041 S.t95 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X102 S.t1040 G D S.t154 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X103 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X104 D G S.t1038 S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X105 S.t1037 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X106 S.t1036 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X107 D G S.t1035 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X108 S.t1034 G D S.t162 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X109 S.t1033 G D S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X110 D G S.t1032 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X111 S.t1031 G D S.t95 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X112 S.t1030 G D S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X113 D G S.t1029 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X114 D G S.t1028 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X115 D G S.t1027 S.t151 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X116 S.t1026 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X117 S.t1025 G D S.t164 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X118 D G S.t1024 S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X119 D G S.t1023 S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X120 D G S.t1022 S.t168 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X121 S.t1021 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X122 S.t1020 G D S.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X123 D G S.t1019 S.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X124 D G S.t1018 S.t107 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X125 S.t1017 G D S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X126 D G S.t1016 S.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X127 S.t1015 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X128 D G S.t1014 S.t95 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X129 D G S.t1013 S.t154 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X130 D G S.t1012 S.t127 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X131 S.t1011 G D S.t95 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X132 D G S.t1010 S.t154 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X133 S.t1009 G D S.t135 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X134 D G S.t1008 S.t140 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X135 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X136 D G S.t1006 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X137 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X138 D G S.t1004 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X139 S.t1003 G D S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X140 S.t1002 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X141 D G S.t1001 S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X142 D G S.t1000 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X143 D G S.t999 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X144 S.t998 G D S.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X145 S.t997 G D S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X146 S.t996 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X147 D G S.t995 S.t107 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X148 D G S.t994 S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X149 S.t993 G D S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X150 S.t992 G D S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X151 S.t991 G D S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X152 S.t990 G D S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X153 S.t989 G D S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X154 S.t988 G D S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X155 D G S.t987 S.t162 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X156 S.t986 G D S.t107 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X157 D G S.t985 S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X158 S.t984 G D S.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X159 S.t983 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X160 D G S.t982 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X161 S.t981 G D S.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X162 S.t980 G D S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X163 S.t979 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X164 S.t978 G D S.t127 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X165 S.t977 G D S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X166 D G S.t976 S.t48 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X167 D G S.t975 S.t135 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X168 S.t974 G D S.t140 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X169 S.t973 G D S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X170 S.t972 G D S.t168 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X171 D G S.t971 S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X172 D G S.t970 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X173 D G S.t969 S.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X174 S.t968 G D S.t135 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X175 S.t967 G D S.t107 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X176 D G S.t966 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X177 D G S.t965 S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X178 D G S.t964 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X179 S.t963 G D S.t127 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X180 D G S.t962 S.t48 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X181 S.t961 G D S.t168 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X182 D G S.t960 S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X183 D G S.t959 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X184 D G S.t958 S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X185 D G S.t957 S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X186 S.t956 G D S.t164 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X187 S.t955 G D S.t162 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X188 D G S.t954 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X189 D G S.t953 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X190 D G S.t952 S.t107 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X191 S.t951 G D S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X192 S.t950 G D S.t151 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X193 D G S.t949 S.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X194 D G S.t948 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X195 D G S.t947 S.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X196 D G S.t946 S.t127 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X197 D G S.t945 S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X198 S.t944 G D S.t48 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X199 S.t943 G D S.t135 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X200 S.t942 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X201 D G S.t941 S.t140 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X202 D G S.t940 S.t140 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X203 D G S.t939 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X204 S.t938 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X205 S.t937 G D S.t151 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X206 D G S.t936 S.t135 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X207 S.t935 G D S.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X208 S.t934 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X209 S.t933 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X210 D G S.t932 S.t107 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X211 D G S.t931 S.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X212 D G S.t930 S.t127 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X213 S.t929 G D S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X214 S.t928 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X215 S.t927 G D S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X216 S.t926 G D S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X217 D G S.t925 S.t168 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X218 S.t924 G D S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X219 S.t923 G D S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X220 D G S.t922 S.t164 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X221 D G S.t921 S.t162 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X222 D G S.t920 S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X223 S.t919 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X224 S.t918 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X225 D G S.t917 S.t151 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X226 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X227 D G S.t915 S.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X228 S.t914 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X229 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X230 D G S.t912 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X231 S.t911 G D S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X232 S.t910 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X233 D G S.t909 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X234 S.t908 G D S.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X235 S.t907 G D S.t140 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X236 S.t906 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X237 D G S.t905 S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X238 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X239 D G S.t903 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X240 S.t902 G D S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X241 S.t901 G D S.t135 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X242 D G S.t900 S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X243 D G S.t899 S.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X244 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X245 S.t897 G D S.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X246 S.t896 G D S.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X247 S.t895 G D S.t127 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X248 D G S.t894 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X249 D G S.t893 S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X250 S.t892 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X251 S.t891 G D S.t168 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X252 S.t890 G D S.t164 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X253 S.t889 G D S.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X254 S.t888 G D S.t95 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X255 D G S.t887 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X256 D G S.t886 S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X257 S.t885 G D S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X258 S.t884 G D S.t95 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X259 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X260 S.t882 G D S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X261 D G S.t881 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X262 S.t880 G D S.t154 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X263 D G S.t879 S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X264 S.t878 G D S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X265 D G S.t877 S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X266 D G S.t876 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X267 S.t875 G D S.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X268 S.t874 G D S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X269 D G S.t873 S.t140 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X270 D G S.t872 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X271 D G S.t871 S.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X272 D G S.t870 S.t135 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X273 D G S.t869 S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X274 S.t868 G D S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X275 D G S.t867 S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X276 D G S.t866 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X277 S.t865 G D S.t48 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X278 D G S.t864 S.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X279 D G S.t863 S.t154 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X280 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X281 S.t861 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X282 S.t860 G D S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X283 D G S.t859 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X284 D G S.t858 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X285 S.t857 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X286 D G S.t856 S.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X287 S.t855 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X288 D G S.t854 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X289 S.t853 G D S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X290 S.t852 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X291 D G S.t851 S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X292 S.t850 G D S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X293 D G S.t849 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X294 S.t848 G D S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X295 D G S.t847 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X296 S.t846 G D S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X297 D G S.t845 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X298 S.t844 G D S.t107 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X299 D G S.t843 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X300 S.t842 G D S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X301 D G S.t841 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X302 D G S.t840 S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X303 D G S.t839 S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X304 S.t838 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X305 D G S.t837 S.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X306 S.t836 G D S.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X307 D G S.t835 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X308 S.t834 G D S.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X309 D G S.t833 S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X310 S.t832 G D S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X311 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X312 S.t830 G D S.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X313 D G S.t829 S.t48 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X314 D G S.t828 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X315 S.t827 G D S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X316 D G S.t826 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X317 S.t825 G D S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X318 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X319 S.t823 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X320 D G S.t822 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X321 D G S.t821 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X322 S.t820 G D S.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X323 D G S.t819 S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X324 D G S.t818 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X325 S.t817 G D S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X326 D G S.t816 S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X327 S.t815 G D S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X328 D G S.t814 S.t48 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X329 D G S.t813 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X330 S.t812 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X331 D G S.t811 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X332 S.t810 G D S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X333 D G S.t809 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X334 D G S.t808 S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X335 D G S.t807 S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X336 S.t806 G D S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X337 S.t805 G D S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X338 D G S.t804 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X339 D G S.t803 S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X340 S.t802 G D S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X341 D G S.t801 S.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X342 S.t800 G D S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X343 S.t799 G D S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X344 S.t798 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X345 S.t797 G D S.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X346 D G S.t796 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X347 S.t795 G D S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X348 S.t794 G D S.t48 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X349 S.t793 G D S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X350 D G S.t792 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X351 S.t791 G D S.t162 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X352 D G S.t790 S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X353 D G S.t789 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X354 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X355 D G S.t787 S.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X356 S.t786 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X357 S.t785 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X358 S.t784 G D S.t151 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X359 D G S.t783 S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X360 D G S.t782 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X361 S.t781 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X362 S.t780 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X363 D G S.t779 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X364 S.t778 G D S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X365 D G S.t777 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X366 D G S.t776 S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X367 D G S.t775 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X368 S.t774 G D S.t162 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X369 S.t773 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X370 D G S.t772 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X371 D G S.t771 S.t162 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X372 D G S.t770 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X373 D G S.t769 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X374 S.t768 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X375 S.t767 G D S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X376 D G S.t766 S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X377 S.t765 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X378 D G S.t764 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X379 S.t763 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X380 S.t762 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X381 D G S.t761 S.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X382 D G S.t760 S.t127 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X383 D G S.t759 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X384 S.t758 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X385 S.t757 G D S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X386 D G S.t756 S.t168 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X387 S.t755 G D S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X388 D G S.t754 S.t48 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X389 D G S.t753 S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X390 S.t752 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X391 S.t751 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X392 D G S.t750 S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X393 S.t749 G D S.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X394 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X395 S.t747 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X396 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X397 S.t745 G D S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X398 D G S.t744 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X399 D G S.t743 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X400 S.t742 G D S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X401 S.t741 G D S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X402 D G S.t740 S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X403 S.t739 G D S.t127 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X404 S.t738 G D S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X405 D G S.t737 S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X406 S.t736 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X407 D G S.t735 S.t162 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X408 D G S.t734 S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X409 S.t733 G D S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X410 D G S.t732 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X411 S.t731 G D S.t168 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X412 D G S.t730 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X413 D G S.t729 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X414 S.t728 G D S.t164 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X415 S.t727 G D S.t151 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X416 D G S.t726 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X417 D G S.t725 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X418 D G S.t724 S.t164 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X419 S.t723 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X420 D G S.t722 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X421 S.t721 G D S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X422 S.t720 G D S.t168 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X423 D G S.t719 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X424 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X425 D G S.t717 S.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X426 D G S.t716 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X427 S.t715 G D S.t107 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X428 D G S.t714 S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X429 S.t713 G D S.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X430 D G S.t712 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X431 S.t711 G D S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X432 D G S.t710 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X433 S.t709 G D S.t95 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X434 D G S.t708 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X435 D G S.t707 S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X436 D G S.t706 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X437 S.t705 G D S.t154 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X438 D G S.t704 S.t140 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X439 D G S.t703 S.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X440 S.t702 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X441 S.t701 G D S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X442 D G S.t700 S.t95 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X443 S.t699 G D S.t154 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X444 D G S.t698 S.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X445 S.t697 G D S.t127 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X446 D G S.t696 S.t135 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X447 S.t695 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X448 D G S.t694 S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X449 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X450 S.t692 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X451 D G S.t691 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X452 D G S.t690 S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X453 S.t689 G D S.t162 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X454 S.t688 G D S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X455 D G S.t687 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X456 D G S.t686 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X457 S.t685 G D S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X458 S.t684 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X459 D G S.t683 S.t151 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X460 D G S.t682 S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X461 S.t681 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X462 S.t680 G D S.t164 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X463 S.t679 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X464 S.t678 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X465 D G S.t677 S.t168 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X466 D G S.t676 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X467 D G S.t675 S.t107 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X468 S.t674 G D S.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X469 S.t673 G D S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X470 S.t672 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X471 S.t671 G D S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X472 D G S.t670 S.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X473 S.t669 G D S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X474 S.t668 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X475 S.t667 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X476 D G S.t666 S.t95 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X477 S.t665 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X478 D G S.t664 S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X479 D G S.t663 S.t154 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X480 S.t662 G D S.t95 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X481 S.t661 G D S.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X482 D G S.t660 S.t154 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X483 D G S.t659 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X484 D G S.t658 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X485 D G S.t657 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X486 S.t656 G D S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X487 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X488 D G S.t654 S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X489 S.t653 G D S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X490 S.t652 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X491 D G S.t651 S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X492 S.t650 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X493 D G S.t649 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X494 S.t648 G D S.t151 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X495 D G S.t647 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X496 D G S.t646 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X497 S.t645 G D S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X498 D G S.t644 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X499 D G S.t643 S.t164 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X500 S.t642 G D S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X501 S.t641 G D S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X502 S.t640 G D S.t168 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X503 D G S.t639 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X504 S.t638 G D S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X505 D G S.t637 S.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X506 S.t636 G D S.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X507 S.t635 G D S.t107 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X508 D G S.t634 S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X509 S.t633 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X510 S.t632 G D S.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X511 D G S.t631 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X512 S.t630 G D S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X513 S.t629 G D S.t95 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X514 S.t628 G D S.t127 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X515 S.t627 G D S.t154 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X516 D G S.t626 S.t48 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X517 D G S.t625 S.t135 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X518 D G S.t624 S.t95 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X519 S.t623 G D S.t154 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X520 S.t622 G D S.t140 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X521 S.t621 G D S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X522 S.t620 G D S.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X523 D G S.t619 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X524 S.t618 G D S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X525 D G S.t617 S.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X526 D G S.t616 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X527 S.t615 G D S.t107 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X528 D G S.t614 S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X529 D G S.t613 S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X530 D G S.t612 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X531 D G S.t611 S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X532 D G S.t610 S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X533 D G S.t609 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X534 S.t608 G D S.t162 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X535 D G S.t607 S.t107 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X536 S.t606 G D S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X537 D G S.t605 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X538 D G S.t604 S.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X539 D G S.t603 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X540 S.t602 G D S.t151 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X541 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X542 D G S.t600 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X543 D G S.t599 S.t127 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X544 D G S.t598 S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X545 S.t597 G D S.t135 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X546 S.t596 G D S.t48 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X547 D G S.t595 S.t140 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X548 D G S.t594 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X549 S.t593 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X550 D G S.t592 S.t140 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X551 D G S.t591 S.t135 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X552 S.t590 G D S.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X553 D G S.t589 S.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X554 S.t588 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X555 S.t587 G D S.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X556 D G S.t586 S.t107 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X557 S.t585 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X558 D G S.t584 S.t127 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X559 S.t583 G D S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X560 S.t582 G D S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X561 S.t581 G D S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X562 S.t580 G D S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X563 D G S.t579 S.t168 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X564 D G S.t578 S.t162 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X565 S.t577 G D S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X566 S.t576 G D S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X567 D G S.t575 S.t164 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X568 D G S.t574 S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X569 S.t573 G D S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X570 S.t572 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X571 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X572 D G S.t570 S.t151 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X573 S.t569 G D S.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X574 S.t568 G D S.t127 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X575 D G S.t567 S.t48 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X576 D G S.t566 S.t164 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X577 D G S.t565 S.t135 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X578 S.t564 G D S.t140 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X579 D G S.t563 S.t164 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X580 S.t562 G D S.t140 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X581 S.t561 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X582 D G S.t560 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X583 D G S.t559 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X584 D G S.t558 S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X585 S.t557 G D S.t135 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X586 D G S.t556 S.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X587 D G S.t555 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X588 S.t554 G D S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X589 S.t553 G D S.t107 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X590 D G S.t552 S.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X591 S.t551 G D S.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X592 S.t550 G D S.t127 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X593 D G S.t549 S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X594 D G S.t548 S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X595 S.t547 G D S.t168 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X596 D G S.t546 S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X597 S.t545 G D S.t164 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X598 S.t544 G D S.t162 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X599 S.t543 G D S.t151 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X600 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X601 D G S.t541 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X602 S.t540 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X603 D G S.t539 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X604 S.t538 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X605 S.t537 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X606 D G S.t536 S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X607 S.t535 G D S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X608 D G S.t534 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X609 D G S.t533 S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X610 S.t532 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X611 S.t531 G D S.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X612 D G S.t530 S.t140 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X613 D G S.t529 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X614 D G S.t528 S.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X615 S.t527 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X616 D G S.t526 S.t135 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X617 S.t525 G D S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X618 D G S.t524 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X619 D G S.t523 S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X620 D G S.t522 S.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X621 D G S.t521 S.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X622 D G S.t520 S.t127 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X623 S.t519 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X624 S.t518 G D S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X625 D G S.t517 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X626 D G S.t516 S.t168 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X627 D G S.t515 S.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X628 D G S.t514 S.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X629 D G S.t513 S.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X630 S.t512 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X631 S.t511 G D S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X632 D G S.t510 S.t95 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X633 S.t509 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X634 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X635 S.t507 G D S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X636 D G S.t506 S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X637 D G S.t505 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X638 S.t504 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X639 D G S.t503 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X640 S.t502 G D S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X641 D G S.t501 S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X642 S.t500 G D S.t140 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X643 D G S.t499 S.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X644 S.t498 G D S.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X645 S.t497 G D S.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X646 S.t496 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X647 D G S.t495 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X648 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X649 S.t493 G D S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X650 S.t492 G D S.t95 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X651 S.t491 G D S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X652 S.t490 G D S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X653 D G S.t489 S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X654 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X655 D G S.t487 S.t48 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X656 S.t486 G D S.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X657 S.t485 G D S.t154 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X658 D G S.t484 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X659 D G S.t483 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X660 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X661 S.t481 G D S.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X662 D G S.t480 S.t154 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X663 S.t479 G D S.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X664 D G S.t478 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X665 D G S.t477 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X666 S.t476 G D S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X667 S.t475 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X668 D G S.t474 S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X669 S.t473 G D S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X670 S.t472 G D S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X671 D G S.t471 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X672 D G S.t470 S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X673 S.t469 G D S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X674 D G S.t468 S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X675 S.t467 G D S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X676 S.t466 G D S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X677 D G S.t465 S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X678 S.t464 G D S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X679 D G S.t463 S.t107 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X680 S.t462 G D S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X681 D G S.t461 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X682 S.t460 G D S.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X683 S.t459 G D S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X684 D G S.t458 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X685 S.t457 G D S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X686 S.t456 G D S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X687 D G S.t455 S.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X688 D G S.t454 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X689 S.t453 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X690 S.t452 G D S.t48 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X691 S.t451 G D S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X692 S.t450 G D S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X693 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X694 D G S.t448 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X695 S.t447 G D S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X696 S.t446 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X697 D G S.t445 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X698 S.t444 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X699 D G S.t443 S.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X700 S.t442 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X701 S.t441 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X702 D G S.t440 S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X703 S.t439 G D S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X704 S.t438 G D S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X705 D G S.t437 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X706 S.t436 G D S.t48 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X707 D G S.t435 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X708 D G S.t434 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X709 S.t433 G D S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X710 D G S.t432 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X711 S.t431 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X712 S.t430 G D S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X713 D G S.t429 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X714 S.t428 G D S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X715 D G S.t427 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X716 D G S.t426 S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X717 D G S.t425 S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X718 D G S.t424 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X719 S.t423 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X720 D G S.t422 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X721 S.t421 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X722 D G S.t420 S.t48 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X723 S.t419 G D S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X724 S.t418 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X725 S.t417 G D S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X726 D G S.t416 S.t48 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X727 D G S.t415 S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X728 D G S.t414 S.t164 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X729 S.t413 G D S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X730 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X731 S.t411 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X732 D G S.t410 S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X733 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X734 D G S.t408 S.t151 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X735 S.t407 G D S.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X736 D G S.t406 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X737 S.t405 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X738 S.t404 G D S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X739 S.t403 G D S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X740 D G S.t402 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X741 S.t401 G D S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X742 D G S.t400 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X743 D G S.t399 S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X744 S.t398 G D S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X745 D G S.t397 S.t162 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X746 S.t396 G D S.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X747 S.t395 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X748 D G S.t394 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X749 D G S.t393 S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X750 S.t392 G D S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X751 D G S.t391 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X752 S.t390 G D S.t162 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X753 S.t389 G D S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X754 D G S.t388 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X755 D G S.t387 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X756 S.t386 G D S.t151 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X757 S.t385 G D S.t135 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X758 S.t384 G D S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X759 D G S.t383 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X760 S.t382 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X761 D G S.t381 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X762 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X763 D G S.t379 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X764 S.t378 G D S.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X765 D G S.t377 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X766 D G S.t376 S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X767 D G S.t375 S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X768 D G S.t374 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X769 S.t373 G D S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X770 D G S.t372 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X771 S.t371 G D S.t154 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X772 D G S.t370 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X773 S.t369 G D S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X774 D G S.t368 S.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X775 D G S.t367 S.t95 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X776 S.t366 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X777 D G S.t365 S.t135 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X778 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X779 D G S.t363 S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X780 D G S.t362 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X781 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X782 S.t360 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X783 S.t359 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X784 D G S.t358 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X785 S.t357 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X786 S.t356 G D S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X787 D G S.t355 S.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X788 D G S.t354 S.t127 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X789 D G S.t353 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X790 S.t352 G D S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X791 D G S.t351 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X792 S.t350 G D S.t162 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X793 D G S.t349 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X794 S.t348 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X795 D G S.t347 S.t168 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X796 S.t346 G D S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X797 D G S.t345 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X798 D G S.t344 S.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X799 S.t343 G D S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X800 D G S.t342 S.t151 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X801 S.t341 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X802 D G S.t340 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X803 S.t339 G D S.t164 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X804 D G S.t338 S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X805 S.t337 G D S.t140 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X806 S.t336 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X807 S.t335 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X808 D G S.t334 S.t168 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X809 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X810 S.t332 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X811 D G S.t331 S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X812 S.t330 G D S.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X813 D G S.t329 S.t107 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X814 S.t328 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X815 S.t327 G D S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X816 D G S.t326 S.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X817 S.t325 G D S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X818 S.t324 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X819 D G S.t323 S.t95 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X820 S.t322 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X821 D G S.t321 S.t162 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X822 D G S.t320 S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X823 D G S.t319 S.t154 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X824 S.t318 G D S.t140 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X825 S.t317 G D S.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X826 S.t316 G D S.t95 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X827 D G S.t315 S.t154 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X828 S.t314 G D S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X829 S.t313 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X830 D G S.t312 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X831 D G S.t311 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X832 D G S.t310 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X833 S.t309 G D S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X834 D G S.t308 S.t162 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X835 D G S.t307 S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X836 S.t306 G D S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X837 D G S.t305 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X838 D G S.t304 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X839 D G S.t303 S.t154 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X840 S.t302 G D S.t151 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X841 S.t301 G D S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X842 D G S.t300 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X843 S.t299 G D S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X844 D G S.t298 S.t164 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X845 S.t297 G D S.t168 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X846 D G S.t296 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X847 S.t295 G D S.t107 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X848 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X849 D G S.t293 S.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X850 D G S.t292 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X851 S.t291 G D S.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X852 D G S.t290 S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X853 S.t289 G D S.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X854 S.t288 G D S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X855 D G S.t287 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X856 D G S.t286 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X857 S.t285 G D S.t95 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X858 S.t284 G D S.t154 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X859 D G S.t283 S.t95 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X860 S.t282 G D S.t154 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X861 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X862 S.t280 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X863 S.t279 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X864 D G S.t278 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X865 D G S.t277 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X866 D G S.t276 S.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X867 S.t275 G D S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X868 S.t274 G D S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X869 D G S.t273 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X870 D G S.t272 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X871 D G S.t271 S.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X872 S.t270 G D S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X873 D G S.t269 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X874 S.t268 G D S.t107 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X875 D G S.t267 S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X876 S.t266 G D S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X877 D G S.t265 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X878 D G S.t264 S.t151 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X879 S.t263 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X880 D G S.t262 S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X881 S.t261 G D S.t164 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X882 D G S.t260 S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X883 D G S.t259 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X884 D G S.t258 S.t168 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X885 D G S.t257 S.t107 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X886 S.t256 G D S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X887 S.t255 G D S.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X888 S.t254 G D S.t162 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X889 D G S.t253 S.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X890 D G S.t252 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X891 D G S.t251 S.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X892 D G S.t250 S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X893 D G S.t249 S.t95 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X894 D G S.t248 S.t127 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X895 S.t247 G D S.t48 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X896 S.t246 G D S.t135 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X897 D G S.t245 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X898 D G S.t244 S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X899 D G S.t243 S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X900 D G S.t242 S.t140 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X901 S.t241 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X902 S.t240 G D S.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X903 S.t239 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X904 D G S.t238 S.t107 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X905 S.t237 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X906 S.t236 G D S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X907 S.t235 G D S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X908 D G S.t234 S.t127 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X909 S.t233 G D S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X910 S.t232 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X911 S.t231 G D S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X912 S.t230 G D S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X913 S.t229 G D S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X914 S.t228 G D S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X915 D G S.t227 S.t164 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X916 D G S.t226 S.t162 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X917 D G S.t225 S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X918 S.t224 G D S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X919 S.t223 G D S.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X920 S.t222 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X921 D G S.t221 S.t151 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X922 S.t220 G D S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X923 S.t219 G D S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X924 S.t218 G D S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X925 S.t217 G D S.t127 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X926 D G S.t216 S.t48 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X927 D G S.t215 S.t135 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X928 S.t214 G D S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X929 S.t213 G D S.t140 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X930 S.t212 G D S.t140 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X931 S.t211 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X932 D G S.t210 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X933 S.t209 G D S.t135 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X934 D G S.t208 S.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X935 D G S.t207 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X936 S.t206 G D S.t107 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X937 S.t205 G D S.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X938 S.t204 G D S.t127 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X939 S.t203 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X940 D G S.t202 S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X941 D G S.t201 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X942 D G S.t200 S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X943 D G S.t199 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X944 S.t198 G D S.t168 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X945 D G S.t197 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X946 D G S.t196 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X947 D G S.t195 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X948 S.t194 G D S.t164 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X949 S.t193 G D S.t162 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X950 S.t192 G D S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X951 D G S.t191 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X952 D G S.t190 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X953 S.t189 G D S.t151 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X954 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X955 D G S.t187 S.t127 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X956 S.t186 G D S.t48 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X957 S.t185 G D S.t168 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X958 S.t184 G D S.t135 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X959 D G S.t183 S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X960 D G S.t182 S.t140 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X961 S.t181 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X962 D G S.t180 S.t140 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X963 D G S.t179 S.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X964 D G S.t178 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X965 S.t177 G D S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X966 S.t176 G D S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X967 D G S.t175 S.t135 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X968 D G S.t174 S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X969 S.t173 G D S.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X970 D G S.t172 S.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X971 D G S.t171 S.t127 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X972 D G S.t170 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X973 D G S.t169 S.t168 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X974 S.t167 G D S.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X975 D G S.t165 S.t164 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X976 D G S.t163 S.t162 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X977 D G S.t161 S.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X978 S.t160 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X979 D G S.t159 S.t151 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X980 S.t158 G D S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X981 D G S.t157 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X982 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X983 D G S.t155 S.t154 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X984 S.t153 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X985 S.t152 G D S.t151 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X986 D G S.t150 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X987 D G S.t149 S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X988 S.t148 G D S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X989 D G S.t147 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X990 S.t146 G D S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X991 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X992 S.t144 G D S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X993 S.t143 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X994 D G S.t142 S.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X995 S.t141 G D S.t140 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X996 D G S.t139 S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X997 S.t138 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X998 S.t137 G D S.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X999 S.t136 G D S.t135 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1000 S.t134 G D S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1001 D G S.t133 S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1002 S.t132 G D S.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1003 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1004 S.t130 G D S.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1005 S.t128 G D S.t127 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1006 D G S.t126 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1007 D G S.t125 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1008 S.t124 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1009 S.t123 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1010 S.t122 G D S.t107 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1011 S.t121 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1012 D G S.t120 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1013 D G S.t119 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1014 S.t118 G D S.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1015 S.t117 G D S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1016 D G S.t116 S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1017 D G S.t115 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1018 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1019 S.t113 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1020 D G S.t112 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1021 S.t111 G D S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1022 D G S.t110 S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1023 S.t109 G D S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1024 D G S.t108 S.t107 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1025 D G S.t106 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1026 S.t105 G D S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1027 D G S.t104 S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1028 S.t103 G D S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1029 S.t102 G D S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1030 S.t101 G D S.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1031 D G S.t100 S.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1032 D G S.t98 S.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1033 S.t97 G D S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1034 D G S.t96 S.t95 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1035 D G S.t94 S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1036 S.t93 G D S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1037 D G S.t92 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1038 D G S.t91 S.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1039 S.t90 G D S.t48 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1040 D G S.t89 S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1041 S.t88 G D S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1042 S.t87 G D S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1043 D G S.t86 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1044 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1045 D G S.t84 S.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1046 D G S.t83 S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1047 D G S.t82 S.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1048 S.t81 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1049 S.t80 G D S.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1050 S.t78 G D S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1051 D G S.t77 S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1052 D G S.t76 S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1053 S.t75 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1054 D G S.t74 S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1055 S.t73 G D S.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1056 S.t71 G D S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1057 D G S.t70 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1058 D G S.t69 S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1059 S.t68 G D S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1060 S.t67 G D S.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1061 S.t65 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1062 S.t64 G D S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1063 D G S.t63 S.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1064 D G S.t61 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1065 D G S.t60 S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1066 D G S.t59 S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1067 D G S.t58 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1068 S.t57 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1069 D G S.t56 S.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1070 D G S.t54 S.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1071 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1072 S.t51 G D S.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1073 D G S.t49 S.t48 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1074 D G S.t47 S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1075 D G S.t46 S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1076 D G S.t45 S.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1077 S.t43 G D S.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1078 S.t0 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1079 D G S.t40 S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1080 S.t39 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1081 S.t38 G D S.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1082 D G S.t0 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1083 D G S.t35 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1084 S.t34 G D S.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1085 S.t32 G D S.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1086 D G S.t30 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1087 D G S.t29 S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1088 D G S.t28 S.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1089 S.t26 G D S.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1090 S.t24 G D S.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1091 S.t22 G D S.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1092 S.t20 G D S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1093 D G S.t19 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1094 D G S.t18 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1095 S.t17 G D S.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1096 S.t15 G D S.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1097 S.t13 G D S.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1098 D G S.t11 S.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1099 S.t9 G D S.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1100 S.t7 G D S.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1101 S.t5 G D S.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1102 D G S.t3 S.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
X1103 D G S.t1 S.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4.38e+06u l=500000u
R0 S.n660 S.n658 169.035
R1 S.n1219 S.n1218 169.035
R2 S.n1782 S.n1781 169.035
R3 S.n2332 S.n2331 169.035
R4 S.n2873 S.n2872 169.035
R5 S.n3388 S.n3387 169.035
R6 S.n3894 S.n3893 169.035
R7 S.n4372 S.n4371 169.035
R8 S.n660 S.n659 169.035
R9 S.n4370 S.n4369 138.167
R10 S.n3892 S.n3891 138.167
R11 S.n3386 S.n3385 138.167
R12 S.n2871 S.n2870 138.167
R13 S.n2330 S.n2329 138.167
R14 S.n1780 S.n1779 138.167
R15 S.n1217 S.n1216 138.167
R16 S.n657 S.n656 138.167
R17 S.n313 S.n312 135.791
R18 S.n975 S.n974 135.791
R19 S.n1521 S.n1520 135.791
R20 S.n2135 S.n2134 135.791
R21 S.n2678 S.n2677 135.791
R22 S.n3195 S.n3194 135.791
R23 S.n3581 S.n3580 135.791
R24 S.n5238 S.n5237 91.519
R25 S.n324 S.n323 91.519
R26 S.n3207 S.n3206 91.519
R27 S.n3592 S.n3591 91.519
R28 S.n4197 S.n4196 91.519
R29 S.n4649 S.n4648 91.519
R30 S.n5032 S.n5031 91.519
R31 S.n2147 S.n2146 91.519
R32 S.n2689 S.n2688 91.519
R33 S.n987 S.n986 91.519
R34 S.n1532 S.n1531 91.519
R35 S.n646 S.n645 91.519
R36 S.n1210 S.n1209 91.519
R37 S.n1771 S.n1770 91.519
R38 S.n2321 S.n2320 91.519
R39 S.n2862 S.n2861 91.519
R40 S.n3377 S.n3376 91.519
R41 S.n3883 S.n3882 91.519
R42 S.n4363 S.n4362 91.519
R43 S.n4812 S.n4811 91.519
R44 S.n5491 S.n5490 91.519
R45 S.n5303 S.n5302 87.091
R46 S.n142 S.n141 87.091
R47 S.n139 S.n138 87.091
R48 S.n91 S.n90 87.091
R49 S.n154 S.n153 87.091
R50 S.n106 S.n105 87.091
R51 S.n120 S.n119 87.091
R52 S.n130 S.n129 87.091
R53 S.n79 S.n78 87.091
R54 S.n150 S.n149 87.091
R55 S.n67 S.n66 87.091
R56 S.n146 S.n145 87.091
R57 S.n5267 S.n5266 87.091
R58 S.n5271 S.n5270 87.091
R59 S.n5275 S.n5274 87.091
R60 S.n5279 S.n5278 87.091
R61 S.n5283 S.n5282 87.091
R62 S.n5287 S.n5286 87.091
R63 S.n5291 S.n5290 87.091
R64 S.n5295 S.n5294 87.091
R65 S.n5299 S.n5298 87.091
R66 S.n5264 S.n5263 87.091
R67 S.n662 S.t162 73.486
R68 S.n315 S.t6 73.486
R69 S.n1221 S.t166 73.486
R70 S.n977 S.t127 73.486
R71 S.n1784 S.t16 73.486
R72 S.n1523 S.t99 73.486
R73 S.n2334 S.t135 73.486
R74 S.n2137 S.t21 73.486
R75 S.n2875 S.t107 73.486
R76 S.n2680 S.t140 73.486
R77 S.n3390 S.t33 73.486
R78 S.n3197 S.t72 73.486
R79 S.n3896 S.t10 73.486
R80 S.n3583 S.t27 73.486
R81 S.n4374 S.t37 73.486
R82 S.n4187 S.t4 73.486
R83 S.t12 S.n482 70.888
R84 S.t25 S.n940 70.888
R85 S.t151 S.n1163 70.888
R86 S.t55 S.n1477 70.888
R87 S.t42 S.n1686 70.888
R88 S.t164 S.n2021 70.888
R89 S.t8 S.n2282 70.888
R90 S.t154 S.n2542 70.888
R91 S.t168 S.n2807 70.888
R92 S.t14 S.n3051 70.888
R93 S.t95 S.n3306 70.888
R94 S.t129 S.n3537 70.888
R95 S.t53 S.n3674 70.888
R96 S.t23 S.n4011 70.888
R97 S.t66 S.n4260 70.888
R98 S.t50 S.n4455 70.888
R99 S.n5303 S.t659 3.773
R100 S.n5304 S.t138 3.773
R101 S.n5301 S.t529 3.773
R102 S.n5317 S.n5316 3.773
R103 S.n5317 S.t797 3.773
R104 S.n5328 S.t63 3.773
R105 S.n5328 S.n5327 3.773
R106 S.n5325 S.t1069 3.773
R107 S.n5325 S.n5324 3.773
R108 S.n5320 S.n5319 3.773
R109 S.n5320 S.t702 3.773
R110 S.n5058 S.n5057 3.773
R111 S.n5058 S.t203 3.773
R112 S.n5076 S.t45 3.773
R113 S.n5076 S.n5075 3.773
R114 S.n5073 S.t729 3.773
R115 S.n5073 S.n5072 3.773
R116 S.n5061 S.n5060 3.773
R117 S.n5061 S.t113 3.773
R118 S.n5238 S.t808 3.773
R119 S.n5240 S.t792 3.773
R120 S.n5242 S.t652 3.773
R121 S.n5305 S.t112 3.773
R122 S.n5306 S.t170 3.773
R123 S.n324 S.t274 3.773
R124 S.n325 S.t771 3.773
R125 S.n305 S.t630 3.773
R126 S.n625 S.n624 3.773
R127 S.n625 S.t1137 3.773
R128 S.n640 S.t420 3.773
R129 S.n640 S.n639 3.773
R130 S.n643 S.t517 3.773
R131 S.n643 S.n642 3.773
R132 S.n628 S.n627 3.773
R133 S.n628 S.t390 3.773
R134 S.n142 S.t123 3.773
R135 S.n143 S.t934 3.773
R136 S.n140 S.t150 3.773
R137 S.n139 S.t942 3.773
R138 S.n135 S.t237 3.773
R139 S.n136 S.t402 3.773
R140 S.n602 S.n601 3.773
R141 S.n602 S.t1136 3.773
R142 S.n613 S.t416 3.773
R143 S.n613 S.n612 3.773
R144 S.n610 S.t300 3.773
R145 S.n610 S.n609 3.773
R146 S.n605 S.n604 3.773
R147 S.n605 S.t1034 3.773
R148 S.n921 S.n920 3.773
R149 S.n921 S.t26 3.773
R150 S.n938 S.t437 3.773
R151 S.n938 S.n937 3.773
R152 S.n935 S.t320 3.773
R153 S.n935 S.n934 3.773
R154 S.n918 S.n917 3.773
R155 S.n918 S.t327 3.773
R156 S.n5336 S.n5335 3.773
R157 S.n5336 S.t173 3.773
R158 S.n5344 S.t552 3.773
R159 S.n5344 S.n5343 3.773
R160 S.n5347 S.t647 3.773
R161 S.n5347 S.n5346 3.773
R162 S.n5333 S.n5332 3.773
R163 S.n5333 S.t538 3.773
R164 S.n5041 S.n5040 3.773
R165 S.n5041 S.t1066 3.773
R166 S.n5052 S.t286 3.773
R167 S.n5052 S.n5051 3.773
R168 S.n5049 S.t406 3.773
R169 S.n5049 S.n5048 3.773
R170 S.n5038 S.n5037 3.773
R171 S.n5038 S.t263 3.773
R172 S.n4847 S.n4846 3.773
R173 S.n4847 S.t827 3.773
R174 S.n4862 S.t89 3.773
R175 S.n4862 S.n4861 3.773
R176 S.n4859 S.t196 3.773
R177 S.n4859 S.n4858 3.773
R178 S.n4844 S.n4843 3.773
R179 S.n4844 S.t65 3.773
R180 S.n4678 S.n4677 3.773
R181 S.n4678 S.t32 3.773
R182 S.n4689 S.t945 3.773
R183 S.n4689 S.n4688 3.773
R184 S.n4686 S.t539 3.773
R185 S.n4686 S.n4685 3.773
R186 S.n4675 S.n4674 3.773
R187 S.n4675 S.t418 3.773
R188 S.n4438 S.n4437 3.773
R189 S.n4438 S.t908 3.773
R190 S.n4453 S.t179 3.773
R191 S.n4453 S.n4452 3.773
R192 S.n4450 S.t269 3.773
R193 S.n4450 S.n4449 3.773
R194 S.n4435 S.n4434 3.773
R195 S.n4435 S.t153 3.773
R196 S.n4247 S.n4246 3.773
R197 S.n4247 S.t636 3.773
R198 S.n4258 S.t1019 3.773
R199 S.n4258 S.n4257 3.773
R200 S.n4255 S.t1135 3.773
R201 S.n4255 S.n4254 3.773
R202 S.n4244 S.n4243 3.773
R203 S.n4244 S.t996 3.773
R204 S.n3994 S.n3993 3.773
R205 S.n3994 S.t398 3.773
R206 S.n4009 S.t777 3.773
R207 S.n4009 S.n4008 3.773
R208 S.n4006 S.t879 3.773
R209 S.n4006 S.n4005 3.773
R210 S.n3991 S.n3990 3.773
R211 S.n3991 S.t755 3.773
R212 S.n3661 S.n3660 3.773
R213 S.n3661 S.t134 3.773
R214 S.n3672 S.t523 3.773
R215 S.n3672 S.n3671 3.773
R216 S.n3669 S.t612 3.773
R217 S.n3669 S.n3668 3.773
R218 S.n3658 S.n3657 3.773
R219 S.n3658 S.t507 3.773
R220 S.n3520 S.n3519 3.773
R221 S.n3520 S.t897 3.773
R222 S.n3535 S.t172 3.773
R223 S.n3535 S.n3534 3.773
R224 S.n3532 S.t262 3.773
R225 S.n3532 S.n3531 3.773
R226 S.n3517 S.n3516 3.773
R227 S.n3517 S.t235 3.773
R228 S.n3293 S.n3292 3.773
R229 S.n3293 S.t629 3.773
R230 S.n3304 S.t1014 3.773
R231 S.n3304 S.n3303 3.773
R232 S.n3301 S.t1126 3.773
R233 S.n3301 S.n3300 3.773
R234 S.n3290 S.n3289 3.773
R235 S.n3290 S.t991 3.773
R236 S.n3034 S.n3033 3.773
R237 S.n3034 S.t389 3.773
R238 S.n3049 S.t770 3.773
R239 S.n3049 S.n3048 3.773
R240 S.n3046 S.t873 3.773
R241 S.n3046 S.n3045 3.773
R242 S.n3031 S.n3030 3.773
R243 S.n3031 S.t747 3.773
R244 S.n2794 S.n2793 3.773
R245 S.n2794 S.t185 3.773
R246 S.n2805 S.t516 3.773
R247 S.n2805 S.n2804 3.773
R248 S.n2802 S.t607 3.773
R249 S.n2802 S.n2801 3.773
R250 S.n2791 S.n2790 3.773
R251 S.n2791 S.t500 3.773
R252 S.n2525 S.n2524 3.773
R253 S.n2525 S.t371 3.773
R254 S.n2540 S.t303 3.773
R255 S.n2540 S.n2539 3.773
R256 S.n2537 S.t634 3.773
R257 S.n2537 S.n2536 3.773
R258 S.n2522 S.n2521 3.773
R259 S.n2522 S.t268 3.773
R260 S.n2269 S.n2268 3.773
R261 S.n2269 S.t352 3.773
R262 S.n2280 S.t737 3.773
R263 S.n2280 S.n2279 3.773
R264 S.n2277 S.t625 3.773
R265 S.n2277 S.n2276 3.773
R266 S.n2266 S.n2265 3.773
R267 S.n2266 S.t256 3.773
R268 S.n2004 S.n2003 3.773
R269 S.n2004 S.t339 3.773
R270 S.n2019 S.t724 3.773
R271 S.n2019 S.n2018 3.773
R272 S.n2016 S.t617 3.773
R273 S.n2016 S.n2015 3.773
R274 S.n2001 S.n2000 3.773
R275 S.n2001 S.t246 3.773
R276 S.n1673 S.n1672 3.773
R277 S.n1673 S.t324 3.773
R278 S.n1684 S.t710 3.773
R279 S.n1684 S.n1683 3.773
R280 S.n1681 S.t609 3.773
R281 S.n1681 S.n1680 3.773
R282 S.n1670 S.n1669 3.773
R283 S.n1670 S.t240 3.773
R284 S.n1460 S.n1459 3.773
R285 S.n1460 S.t309 3.773
R286 S.n1475 S.t691 3.773
R287 S.n1475 S.n1474 3.773
R288 S.n1472 S.t599 3.773
R289 S.n1472 S.n1471 3.773
R290 S.n1457 S.n1456 3.773
R291 S.n1457 S.t228 3.773
R292 S.n1150 S.n1149 3.773
R293 S.n1150 S.t302 3.773
R294 S.n1161 S.t683 3.773
R295 S.n1161 S.n1160 3.773
R296 S.n1158 S.t714 3.773
R297 S.n1158 S.n1157 3.773
R298 S.n1147 S.n1146 3.773
R299 S.n1147 S.t217 3.773
R300 S.n469 S.n468 3.773
R301 S.n469 S.t13 3.773
R302 S.n480 S.t427 3.773
R303 S.n480 S.n479 3.773
R304 S.n477 S.t308 3.773
R305 S.n477 S.n476 3.773
R306 S.n472 S.n471 3.773
R307 S.n472 S.t1045 3.773
R308 S.n91 S.t279 3.773
R309 S.n84 S.t1086 3.773
R310 S.n85 S.t304 3.773
R311 S.n265 S.n264 3.773
R312 S.n265 S.t186 3.773
R313 S.n276 S.t567 3.773
R314 S.n276 S.n275 3.773
R315 S.n273 S.t657 3.773
R316 S.n273 S.n272 3.773
R317 S.n268 S.n267 3.773
R318 S.n268 S.t544 3.773
R319 S.n776 S.n775 3.773
R320 S.n776 S.t685 3.773
R321 S.n789 S.t1065 3.773
R322 S.n789 S.n788 3.773
R323 S.n786 S.t59 3.773
R324 S.n786 S.n785 3.773
R325 S.n773 S.n772 3.773
R326 S.n773 S.t927 3.773
R327 S.n3207 S.t492 3.773
R328 S.n3208 S.t964 3.773
R329 S.n3188 S.t850 3.773
R330 S.n3058 S.n3057 3.773
R331 S.n3058 S.t220 3.773
R332 S.n3072 S.t600 3.773
R333 S.n3072 S.n3071 3.773
R334 S.n3075 S.t704 3.773
R335 S.n3075 S.n3074 3.773
R336 S.n3055 S.n3054 3.773
R337 S.n3055 S.t585 3.773
R338 S.n2698 S.n2697 3.773
R339 S.n2698 S.t1140 3.773
R340 S.n2709 S.t347 3.773
R341 S.n2709 S.n2708 3.773
R342 S.n2706 S.t463 3.773
R343 S.n2706 S.n2705 3.773
R344 S.n2695 S.n2694 3.773
R345 S.n2695 S.t318 3.773
R346 S.n2378 S.n2377 3.773
R347 S.n2378 S.t880 3.773
R348 S.n2393 S.t155 3.773
R349 S.n2393 S.n2392 3.773
R350 S.n2390 S.t244 3.773
R351 S.n2390 S.n2389 3.773
R352 S.n2375 S.n2374 3.773
R353 S.n2375 S.t122 3.773
R354 S.n2176 S.n2175 3.773
R355 S.n2176 S.t103 3.773
R356 S.n2184 S.t994 3.773
R357 S.n2184 S.n2183 3.773
R358 S.n2168 S.t591 3.773
R359 S.n2168 S.n2167 3.773
R360 S.n2173 S.n2172 3.773
R361 S.n2173 S.t472 3.773
R362 S.n1857 S.n1856 3.773
R363 S.n1857 S.t956 3.773
R364 S.n1872 S.t227 3.773
R365 S.n1872 S.n1871 3.773
R366 S.n1869 S.t326 3.773
R367 S.n1869 S.n1868 3.773
R368 S.n1854 S.n1853 3.773
R369 S.n1854 S.t209 3.773
R370 S.n1577 S.n1576 3.773
R371 S.n1577 S.t692 3.773
R372 S.n1588 S.t1079 3.773
R373 S.n1588 S.n1587 3.773
R374 S.n1585 S.t74 3.773
R375 S.n1585 S.n1584 3.773
R376 S.n1574 S.n1573 3.773
R377 S.n1574 S.t1050 3.773
R378 S.n1311 S.n1310 3.773
R379 S.n1311 S.t457 3.773
R380 S.n1326 S.t835 3.773
R381 S.n1326 S.n1325 3.773
R382 S.n1323 S.t930 3.773
R383 S.n1323 S.n1322 3.773
R384 S.n1308 S.n1307 3.773
R385 S.n1308 S.t810 3.773
R386 S.n1049 S.n1048 3.773
R387 S.n1049 S.t189 3.773
R388 S.n1060 S.t570 3.773
R389 S.n1060 S.n1059 3.773
R390 S.n1057 S.t200 3.773
R391 S.n1057 S.n1056 3.773
R392 S.n1046 S.n1045 3.773
R393 S.n1046 S.t550 3.773
R394 S.n154 S.t765 3.773
R395 S.n155 S.t857 3.773
R396 S.n152 S.t119 3.773
R397 S.n288 S.n287 3.773
R398 S.n288 S.t865 3.773
R399 S.n299 S.t962 3.773
R400 S.n299 S.n298 3.773
R401 S.n296 S.t3 3.773
R402 S.n296 S.n295 3.773
R403 S.n291 S.n290 3.773
R404 S.n291 S.t774 3.773
R405 S.n3592 S.t314 3.773
R406 S.n3593 S.t811 3.773
R407 S.n3572 S.t671 3.773
R408 S.n3548 S.n3547 3.773
R409 S.n3548 S.t1075 3.773
R410 S.n3563 S.t355 3.773
R411 S.n3563 S.n3562 3.773
R412 S.n3566 S.t470 3.773
R413 S.n3566 S.n3565 3.773
R414 S.n3551 S.n3550 3.773
R415 S.n3551 S.t433 3.773
R416 S.n3214 S.n3213 3.773
R417 S.n3214 S.t884 3.773
R418 S.n3225 S.t96 3.773
R419 S.n3225 S.n3224 3.773
R420 S.n3222 S.t201 3.773
R421 S.n3222 S.n3221 3.773
R422 S.n3217 S.n3216 3.773
R423 S.n3217 S.t73 3.773
R424 S.n2911 S.n2910 3.773
R425 S.n2911 S.t618 3.773
R426 S.n2931 S.t999 3.773
R427 S.n2931 S.n2930 3.773
R428 S.n2928 S.t1112 3.773
R429 S.n2928 S.n2927 3.773
R430 S.n2914 S.n2913 3.773
R431 S.n2914 S.t979 3.773
R432 S.n2715 S.n2714 3.773
R433 S.n2715 S.t961 3.773
R434 S.n2726 S.t756 3.773
R435 S.n2726 S.n2725 3.773
R436 S.n2723 S.t329 3.773
R437 S.n2723 S.n2722 3.773
R438 S.n2718 S.n2717 3.773
R439 S.n2718 S.t212 3.773
R440 S.n2402 S.n2401 3.773
R441 S.n2402 S.t699 3.773
R442 S.n2422 S.t1083 3.773
R443 S.n2422 S.n2421 3.773
R444 S.n2419 S.t76 3.773
R445 S.n2419 S.n2418 3.773
R446 S.n2405 S.n2404 3.773
R447 S.n2405 S.t1054 3.773
R448 S.n2190 S.n2189 3.773
R449 S.n2190 S.t459 3.773
R450 S.n2201 S.t840 3.773
R451 S.n2201 S.n2200 3.773
R452 S.n2198 S.t936 3.773
R453 S.n2198 S.n2197 3.773
R454 S.n2193 S.n2192 3.773
R455 S.n2193 S.t817 3.773
R456 S.n1881 S.n1880 3.773
R457 S.n1881 S.t194 3.773
R458 S.n1901 S.t575 3.773
R459 S.n1901 S.n1900 3.773
R460 S.n1898 S.t670 3.773
R461 S.n1898 S.n1897 3.773
R462 S.n1884 S.n1883 3.773
R463 S.n1884 S.t557 3.773
R464 S.n1594 S.n1593 3.773
R465 S.n1594 S.t1037 3.773
R466 S.n1605 S.t311 3.773
R467 S.n1605 S.n1604 3.773
R468 S.n1602 S.t432 3.773
R469 S.n1602 S.n1601 3.773
R470 S.n1597 S.n1596 3.773
R471 S.n1597 S.t289 3.773
R472 S.n1335 S.n1334 3.773
R473 S.n1335 S.t795 3.773
R474 S.n1355 S.t56 3.773
R475 S.n1355 S.n1354 3.773
R476 S.n1352 S.t171 3.773
R477 S.n1352 S.n1351 3.773
R478 S.n1338 S.n1337 3.773
R479 S.n1338 S.t17 3.773
R480 S.n1066 S.n1065 3.773
R481 S.n1066 S.t543 3.773
R482 S.n1079 S.t917 3.773
R483 S.n1079 S.n1078 3.773
R484 S.n1076 S.t546 3.773
R485 S.n1076 S.n1075 3.773
R486 S.n1069 S.n1068 3.773
R487 S.n1069 S.t895 3.773
R488 S.n1087 S.n1086 3.773
R489 S.n1087 S.t937 3.773
R490 S.n1101 S.t159 3.773
R491 S.n1101 S.n1100 3.773
R492 S.n1098 S.t893 3.773
R493 S.n1098 S.n1097 3.773
R494 S.n1090 S.n1089 3.773
R495 S.n1090 S.t128 3.773
R496 S.n827 S.n826 3.773
R497 S.n827 S.t117 3.773
R498 S.n851 S.t712 3.773
R499 S.n851 S.n850 3.773
R500 S.n848 S.t410 3.773
R501 S.n848 S.n847 3.773
R502 S.n830 S.n829 3.773
R503 S.n830 S.t417 3.773
R504 S.n303 S.n302 3.773
R505 S.n303 S.t105 3.773
R506 S.n501 S.t503 3.773
R507 S.n501 S.n500 3.773
R508 S.n504 S.t397 3.773
R509 S.n504 S.n503 3.773
R510 S.n507 S.n506 3.773
R511 S.n507 S.t1130 3.773
R512 S.n515 S.n514 3.773
R513 S.n515 S.t90 3.773
R514 S.n530 S.t487 3.773
R515 S.n530 S.n529 3.773
R516 S.n527 S.t381 3.773
R517 S.n527 S.n526 3.773
R518 S.n518 S.n517 3.773
R519 S.n518 S.t1119 3.773
R520 S.n106 S.t1105 3.773
R521 S.n98 S.t78 3.773
R522 S.n99 S.t478 3.773
R523 S.n1373 S.n1372 3.773
R524 S.n1373 S.t1141 3.773
R525 S.n1388 S.t422 3.773
R526 S.n1388 S.n1387 3.773
R527 S.n1385 S.t520 3.773
R528 S.n1385 S.n1384 3.773
R529 S.n1370 S.n1369 3.773
R530 S.n1370 S.t392 3.773
R531 S.n1918 S.n1917 3.773
R532 S.n1918 S.t545 3.773
R533 S.n1933 S.t922 3.773
R534 S.n1933 S.n1932 3.773
R535 S.n1930 S.t1016 3.773
R536 S.n1930 S.n1929 3.773
R537 S.n1915 S.n1914 3.773
R538 S.n1915 S.t901 3.773
R539 S.n2439 S.n2438 3.773
R540 S.n2439 S.t1040 3.773
R541 S.n2454 S.t315 3.773
R542 S.n2454 S.n2453 3.773
R543 S.n2451 S.t440 3.773
R544 S.n2451 S.n2450 3.773
R545 S.n2436 S.n2435 3.773
R546 S.n2436 S.t295 3.773
R547 S.n2948 S.n2947 3.773
R548 S.n2948 S.t466 3.773
R549 S.n2963 S.t847 3.773
R550 S.n2963 S.n2962 3.773
R551 S.n2960 S.t940 3.773
R552 S.n2960 S.n2959 3.773
R553 S.n2945 S.n2944 3.773
R554 S.n2945 S.t823 3.773
R555 S.n3434 S.n3433 3.773
R556 S.n3434 S.t378 3.773
R557 S.n3449 S.t761 3.773
R558 S.n3449 S.n3448 3.773
R559 S.n3446 S.t867 3.773
R560 S.n3446 S.n3445 3.773
R561 S.n3431 S.n3430 3.773
R562 S.n3431 S.t832 3.773
R563 S.n4021 S.n4020 3.773
R564 S.n4021 S.t923 3.773
R565 S.n4035 S.t197 3.773
R566 S.n4035 S.n4034 3.773
R567 S.n4038 S.t290 3.773
R568 S.n4038 S.n4037 3.773
R569 S.n4018 S.n4017 3.773
R570 S.n4018 S.t177 3.773
R571 S.n4197 S.t67 3.773
R572 S.n4198 S.t558 3.773
R573 S.n4181 S.t441 3.773
R574 S.n3601 S.n3600 3.773
R575 S.n3601 S.t721 3.773
R576 S.n3612 S.t1038 3.773
R577 S.n3612 S.n3611 3.773
R578 S.n3609 S.t19 3.773
R579 S.n3609 S.n3608 3.773
R580 S.n3598 S.n3597 3.773
R581 S.n3598 S.t1017 3.773
R582 S.n3233 S.n3232 3.773
R583 S.n3233 S.t709 3.773
R584 S.n3244 S.t510 3.773
R585 S.n3244 S.n3243 3.773
R586 S.n3241 S.t83 3.773
R587 S.n3241 S.n3240 3.773
R588 S.n3230 S.n3229 3.773
R589 S.n3230 S.t1060 3.773
R590 S.n2734 S.n2733 3.773
R591 S.n2734 S.t198 3.773
R592 S.n2745 S.t579 3.773
R593 S.n2745 S.n2744 3.773
R594 S.n2742 S.t675 3.773
R595 S.n2742 S.n2741 3.773
R596 S.n2731 S.n2730 3.773
R597 S.n2731 S.t562 3.773
R598 S.n2209 S.n2208 3.773
R599 S.n2209 S.t800 3.773
R600 S.n2220 S.t60 3.773
R601 S.n2220 S.n2219 3.773
R602 S.n2217 S.t175 3.773
R603 S.n2217 S.n2216 3.773
R604 S.n2206 S.n2205 3.773
R605 S.n2206 S.t22 3.773
R606 S.n1613 S.n1612 3.773
R607 S.n1613 S.t280 3.773
R608 S.n1624 S.t658 3.773
R609 S.n1624 S.n1623 3.773
R610 S.n1621 S.t772 3.773
R611 S.n1621 S.n1620 3.773
R612 S.n1610 S.n1609 3.773
R613 S.n1610 S.t632 3.773
R614 S.n866 S.n865 3.773
R615 S.n866 S.t473 3.773
R616 S.n885 S.t854 3.773
R617 S.n885 S.n884 3.773
R618 S.n882 S.t750 3.773
R619 S.n882 S.n881 3.773
R620 S.n869 S.n868 3.773
R621 S.n869 S.t757 3.773
R622 S.n429 S.n428 3.773
R623 S.n429 S.t464 3.773
R624 S.n444 S.t841 3.773
R625 S.n444 S.n443 3.773
R626 S.n441 S.t735 3.773
R627 S.n441 S.n440 3.773
R628 S.n432 S.n431 3.773
R629 S.n432 S.t369 3.773
R630 S.n547 S.n546 3.773
R631 S.n547 S.t452 3.773
R632 S.n563 S.t829 3.773
R633 S.n563 S.n562 3.773
R634 S.n560 S.t722 3.773
R635 S.n560 S.n559 3.773
R636 S.n550 S.n549 3.773
R637 S.n550 S.t350 3.773
R638 S.n120 S.t335 3.773
R639 S.n109 S.t442 3.773
R640 S.n110 S.t818 3.773
R641 S.n4649 S.t926 3.773
R642 S.n4650 S.t296 3.773
R643 S.n4638 S.t181 3.773
R644 S.n4469 S.n4468 3.773
R645 S.n4469 S.t661 3.773
R646 S.n4477 S.t1043 3.773
R647 S.n4477 S.n4476 3.773
R648 S.n4480 S.t29 3.773
R649 S.n4480 S.n4479 3.773
R650 S.n4466 S.n4465 3.773
R651 S.n4466 S.t1021 3.773
R652 S.n4211 S.n4210 3.773
R653 S.n4211 S.t481 3.773
R654 S.n4219 S.t801 3.773
R655 S.n4219 S.n4218 3.773
R656 S.n4216 S.t905 3.773
R657 S.n4216 S.n4215 3.773
R658 S.n4208 S.n4207 3.773
R659 S.n4208 S.t780 3.773
R660 S.n3939 S.n3938 3.773
R661 S.n3939 S.t214 3.773
R662 S.n3957 S.t594 3.773
R663 S.n3957 S.n3956 3.773
R664 S.n3954 S.t690 3.773
R665 S.n3954 S.n3953 3.773
R666 S.n3936 S.n3935 3.773
R667 S.n3936 S.t573 3.773
R668 S.n3625 S.n3624 3.773
R669 S.n3625 S.t554 3.773
R670 S.n3633 S.t338 3.773
R671 S.n3633 S.n3632 3.773
R672 S.n3630 S.t1028 3.773
R673 S.n3630 S.n3629 3.773
R674 S.n3622 S.n3621 3.773
R675 S.n3622 S.t911 3.773
R676 S.n3465 S.n3464 3.773
R677 S.n3465 S.t205 3.773
R678 S.n3483 S.t589 3.773
R679 S.n3483 S.n3482 3.773
R680 S.n3480 S.t682 3.773
R681 S.n3480 S.n3479 3.773
R682 S.n3462 S.n3461 3.773
R683 S.n3462 S.t645 3.773
R684 S.n3257 S.n3256 3.773
R685 S.n3257 S.t1047 3.773
R686 S.n3265 S.t323 3.773
R687 S.n3265 S.n3264 3.773
R688 S.n3262 S.t445 3.773
R689 S.n3262 S.n3261 3.773
R690 S.n3254 S.n3253 3.773
R691 S.n3254 S.t301 3.773
R692 S.n2979 S.n2978 3.773
R693 S.n2979 S.t806 3.773
R694 S.n2997 S.t70 3.773
R695 S.n2997 S.n2996 3.773
R696 S.n2994 S.t180 3.773
R697 S.n2994 S.n2993 3.773
R698 S.n2976 S.n2975 3.773
R699 S.n2976 S.t34 3.773
R700 S.n2758 S.n2757 3.773
R701 S.n2758 S.t547 3.773
R702 S.n2766 S.t925 3.773
R703 S.n2766 S.n2765 3.773
R704 S.n2763 S.t1018 3.773
R705 S.n2763 S.n2762 3.773
R706 S.n2755 S.n2754 3.773
R707 S.n2755 S.t907 3.773
R708 S.n2470 S.n2469 3.773
R709 S.n2470 S.t282 3.773
R710 S.n2488 S.t660 3.773
R711 S.n2488 S.n2487 3.773
R712 S.n2485 S.t776 3.773
R713 S.n2485 S.n2484 3.773
R714 S.n2467 S.n2466 3.773
R715 S.n2467 S.t635 3.773
R716 S.n2233 S.n2232 3.773
R717 S.n2233 S.t9 3.773
R718 S.n2241 S.t426 3.773
R719 S.n2241 S.n2240 3.773
R720 S.n2238 S.t526 3.773
R721 S.n2238 S.n2237 3.773
R722 S.n2230 S.n2229 3.773
R723 S.n2230 S.t401 3.773
R724 S.n1949 S.n1948 3.773
R725 S.n1949 S.t890 3.773
R726 S.n1967 S.t165 3.773
R727 S.n1967 S.n1966 3.773
R728 S.n1964 S.t251 3.773
R729 S.n1964 S.n1963 3.773
R730 S.n1946 S.n1945 3.773
R731 S.n1946 S.t136 3.773
R732 S.n1637 S.n1636 3.773
R733 S.n1637 S.t678 3.773
R734 S.n1645 S.t1004 3.773
R735 S.n1645 S.n1644 3.773
R736 S.n1642 S.t1117 3.773
R737 S.n1642 S.n1641 3.773
R738 S.n1634 S.n1633 3.773
R739 S.n1634 S.t981 3.773
R740 S.n1404 S.n1403 3.773
R741 S.n1404 S.t741 3.773
R742 S.n1422 S.t821 3.773
R743 S.n1422 S.n1421 3.773
R744 S.n1419 S.t1012 3.773
R745 S.n1419 S.n1418 3.773
R746 S.n1401 S.n1400 3.773
R747 S.n1401 S.t638 3.773
R748 S.n1114 S.n1113 3.773
R749 S.n1114 S.t727 3.773
R750 S.n1122 S.t1109 3.773
R751 S.n1122 S.n1121 3.773
R752 S.n1119 S.t1138 3.773
R753 S.n1119 S.n1118 3.773
R754 S.n1111 S.n1110 3.773
R755 S.n1111 S.t628 3.773
R756 S.n894 S.n893 3.773
R757 S.n894 S.t815 3.773
R758 S.n913 S.t77 3.773
R759 S.n913 S.n912 3.773
R760 S.n910 S.t1089 3.773
R761 S.n910 S.n909 3.773
R762 S.n897 S.n896 3.773
R763 S.n897 S.t1098 3.773
R764 S.n449 S.n448 3.773
R765 S.n449 S.t802 3.773
R766 S.n463 S.t61 3.773
R767 S.n463 S.n462 3.773
R768 S.n460 S.t1068 3.773
R769 S.n460 S.n459 3.773
R770 S.n452 S.n451 3.773
R771 S.n452 S.t701 3.773
R772 S.n1133 S.n1132 3.773
R773 S.n1133 S.t1061 3.773
R774 S.n1142 S.t342 3.773
R775 S.n1142 S.n1141 3.773
R776 S.n1139 S.t376 3.773
R777 S.n1139 S.n1138 3.773
R778 S.n1130 S.n1129 3.773
R779 S.n1130 S.t978 3.773
R780 S.n1431 S.n1430 3.773
R781 S.n1431 S.t1076 3.773
R782 S.n1443 S.t358 3.773
R783 S.n1443 S.n1442 3.773
R784 S.n1440 S.t248 3.773
R785 S.n1440 S.n1439 3.773
R786 S.n1434 S.n1433 3.773
R787 S.n1434 S.t988 3.773
R788 S.n1651 S.n1650 3.773
R789 S.n1651 S.t1097 3.773
R790 S.n1665 S.t374 3.773
R791 S.n1665 S.n1664 3.773
R792 S.n1662 S.t259 3.773
R793 S.n1662 S.n1661 3.773
R794 S.n1654 S.n1653 3.773
R795 S.n1654 S.t998 3.773
R796 S.n1976 S.n1975 3.773
R797 S.n1976 S.t1107 3.773
R798 S.n1987 S.t563 3.773
R799 S.n1987 S.n1986 3.773
R800 S.n1984 S.t271 3.773
R801 S.n1984 S.n1983 3.773
R802 S.n1979 S.n1978 3.773
R803 S.n1979 S.t1009 3.773
R804 S.n2247 S.n2246 3.773
R805 S.n2247 S.t447 3.773
R806 S.n2261 S.t766 3.773
R807 S.n2261 S.n2260 3.773
R808 S.n2258 S.t870 3.773
R809 S.n2258 S.n2257 3.773
R810 S.n2250 S.n2249 3.773
R811 S.n2250 S.t742 3.773
R812 S.n2497 S.n2496 3.773
R813 S.n2497 S.t623 3.773
R814 S.n2508 S.t1010 3.773
R815 S.n2508 S.n2507 3.773
R816 S.n2505 S.t1123 3.773
R817 S.n2505 S.n2504 3.773
R818 S.n2500 S.n2499 3.773
R819 S.n2500 S.t986 3.773
R820 S.n2772 S.n2771 3.773
R821 S.n2772 S.t891 3.773
R822 S.n2786 S.t169 3.773
R823 S.n2786 S.n2785 3.773
R824 S.n2783 S.t257 3.773
R825 S.n2783 S.n2782 3.773
R826 S.n2775 S.n2774 3.773
R827 S.n2775 S.t141 3.773
R828 S.n3006 S.n3005 3.773
R829 S.n3006 S.t15 3.773
R830 S.n3017 S.t429 3.773
R831 S.n3017 S.n3016 3.773
R832 S.n3014 S.t530 3.773
R833 S.n3014 S.n3013 3.773
R834 S.n3009 S.n3008 3.773
R835 S.n3009 S.t405 3.773
R836 S.n3271 S.n3270 3.773
R837 S.n3271 S.t285 3.773
R838 S.n3285 S.t666 3.773
R839 S.n3285 S.n3284 3.773
R840 S.n3282 S.t782 3.773
R841 S.n3282 S.n3281 3.773
R842 S.n3274 S.n3273 3.773
R843 S.n3274 S.t641 3.773
R844 S.n3492 S.n3491 3.773
R845 S.n3492 S.t551 3.773
R846 S.n3503 S.t931 3.773
R847 S.n3503 S.n3502 3.773
R848 S.n3500 S.t1023 3.773
R849 S.n3500 S.n3499 3.773
R850 S.n3495 S.n3494 3.773
R851 S.n3495 S.t992 3.773
R852 S.n3639 S.n3638 3.773
R853 S.n3639 S.t902 3.773
R854 S.n3653 S.t174 3.773
R855 S.n3653 S.n3652 3.773
R856 S.n3650 S.t265 3.773
R857 S.n3650 S.n3649 3.773
R858 S.n3642 S.n3641 3.773
R859 S.n3642 S.t148 3.773
R860 S.n3966 S.n3965 3.773
R861 S.n3966 S.t24 3.773
R862 S.n3977 S.t435 3.773
R863 S.n3977 S.n3976 3.773
R864 S.n3974 S.t536 3.773
R865 S.n3974 S.n3973 3.773
R866 S.n3969 S.n3968 3.773
R867 S.n3969 S.t413 3.773
R868 S.n4225 S.n4224 3.773
R869 S.n4225 S.t291 3.773
R870 S.n4239 S.t84 3.773
R871 S.n4239 S.n4238 3.773
R872 S.n4236 S.t790 3.773
R873 S.n4236 S.n4235 3.773
R874 S.n4228 S.n4227 3.773
R875 S.n4228 S.t650 3.773
R876 S.n4410 S.n4409 3.773
R877 S.n4410 S.t1064 3.773
R878 S.n4421 S.t344 3.773
R879 S.n4421 S.n4420 3.773
R880 S.n4418 S.t458 3.773
R881 S.n4418 S.n4417 3.773
R882 S.n4413 S.n4412 3.773
R883 S.n4413 S.t313 3.773
R884 S.n4656 S.n4655 3.773
R885 S.n4656 S.t219 3.773
R886 S.n4670 S.t548 3.773
R887 S.n4670 S.n4669 3.773
R888 S.n4667 S.t639 3.773
R889 S.n4667 S.n4666 3.773
R890 S.n4659 S.n4658 3.773
R891 S.n4659 S.t532 3.773
R892 S.n4875 S.n4874 3.773
R893 S.n4875 S.t430 3.773
R894 S.n4883 S.t807 3.773
R895 S.n4883 S.n4882 3.773
R896 S.n4886 S.t909 3.773
R897 S.n4886 S.n4885 3.773
R898 S.n4878 S.n4877 3.773
R899 S.n4878 S.t785 3.773
R900 S.n5032 S.t667 3.773
R901 S.n5033 S.t35 3.773
R902 S.n5023 S.t1026 3.773
R903 S.n130 S.t681 3.773
R904 S.n125 S.t781 3.773
R905 S.n126 S.t30 3.773
R906 S.n573 S.n572 3.773
R907 S.n573 S.t794 3.773
R908 S.n592 S.t49 3.773
R909 S.n592 S.n591 3.773
R910 S.n589 S.t1059 3.773
R911 S.n589 S.n588 3.773
R912 S.n576 S.n575 3.773
R913 S.n576 S.t689 3.773
R914 S.n798 S.n797 3.773
R915 S.n798 S.t1030 3.773
R916 S.n817 S.t305 3.773
R917 S.n817 S.n816 3.773
R918 S.n814 S.t425 3.773
R919 S.n814 S.n813 3.773
R920 S.n801 S.n800 3.773
R921 S.n801 S.t167 3.773
R922 S.n413 S.n412 3.773
R923 S.n413 S.t848 3.773
R924 S.n424 S.t40 3.773
R925 S.n424 S.n423 3.773
R926 S.n421 S.t163 3.773
R927 S.n421 S.n420 3.773
R928 S.n416 S.n415 3.773
R929 S.n416 S.t7 3.773
R930 S.n396 S.n395 3.773
R931 S.n396 S.t451 3.773
R932 S.n407 S.t826 3.773
R933 S.n407 S.n406 3.773
R934 S.n404 S.t921 3.773
R935 S.n404 S.n403 3.773
R936 S.n399 S.n398 3.773
R937 S.n399 S.t799 3.773
R938 S.n79 S.t695 3.773
R939 S.n72 S.t341 3.773
R940 S.n73 S.t725 3.773
R941 S.n221 S.n220 3.773
R942 S.n221 S.t596 3.773
R943 S.n232 S.t976 3.773
R944 S.n232 S.n231 3.773
R945 S.n229 S.t1078 3.773
R946 S.n229 S.n228 3.773
R947 S.n224 S.n223 3.773
R948 S.n224 S.t955 3.773
R949 S.n717 S.n716 3.773
R950 S.n717 S.t1115 3.773
R951 S.n730 S.t391 3.773
R952 S.n730 S.n729 3.773
R953 S.n727 S.t501 3.773
R954 S.n727 S.n726 3.773
R955 S.n714 S.n713 3.773
R956 S.n714 S.t233 3.773
R957 S.n2147 S.t977 3.773
R958 S.n2148 S.t365 3.773
R959 S.n2128 S.t231 3.773
R960 S.n2028 S.n2027 3.773
R961 S.n2028 S.t728 3.773
R962 S.n2042 S.t1114 3.773
R963 S.n2042 S.n2041 3.773
R964 S.n2045 S.t100 3.773
R965 S.n2045 S.n2044 3.773
R966 S.n2025 S.n2024 3.773
R967 S.n2025 S.t1082 3.773
R968 S.n1541 S.n1540 3.773
R969 S.n1541 S.t537 3.773
R970 S.n1552 S.t859 3.773
R971 S.n1552 S.n1551 3.773
R972 S.n1549 S.t953 3.773
R973 S.n1549 S.n1548 3.773
R974 S.n1538 S.n1537 3.773
R975 S.n1538 S.t836 3.773
R976 S.n1250 S.n1249 3.773
R977 S.n1250 S.t266 3.773
R978 S.n1265 S.t646 3.773
R979 S.n1265 S.n1264 3.773
R980 S.n1262 S.t760 3.773
R981 S.n1262 S.n1261 3.773
R982 S.n1247 S.n1246 3.773
R983 S.n1247 S.t621 3.773
R984 S.n1013 S.n1012 3.773
R985 S.n1013 S.t602 3.773
R986 S.n1024 S.t408 3.773
R987 S.n1024 S.n1023 3.773
R988 S.n1021 S.t613 3.773
R989 S.n1021 S.n1020 3.773
R990 S.n1010 S.n1009 3.773
R991 S.n1010 S.t963 3.773
R992 S.n150 S.t1036 3.773
R993 S.n151 S.t684 3.773
R994 S.n148 S.t1063 3.773
R995 S.n244 S.n243 3.773
R996 S.n244 S.t944 3.773
R997 S.n255 S.t216 3.773
R998 S.n255 S.n254 3.773
R999 S.n252 S.t310 3.773
R1000 S.n252 S.n251 3.773
R1001 S.n247 S.n246 3.773
R1002 S.n247 S.t193 3.773
R1003 S.n2689 S.t731 3.773
R1004 S.n2690 S.t108 3.773
R1005 S.n2669 S.t1088 3.773
R1006 S.n2553 S.n2552 3.773
R1007 S.n2553 S.t485 3.773
R1008 S.n2568 S.t863 3.773
R1009 S.n2568 S.n2567 3.773
R1010 S.n2571 S.t958 3.773
R1011 S.n2571 S.n2570 3.773
R1012 S.n2556 S.n2555 3.773
R1013 S.n2556 S.t844 3.773
R1014 S.n2154 S.n2153 3.773
R1015 S.n2154 S.t270 3.773
R1016 S.n2165 S.t598 3.773
R1017 S.n2165 S.n2164 3.773
R1018 S.n2162 S.t696 3.773
R1019 S.n2162 S.n2161 3.773
R1020 S.n2157 S.n2156 3.773
R1021 S.n2157 S.t580 3.773
R1022 S.n1820 S.n1819 3.773
R1023 S.n1820 S.t1132 3.773
R1024 S.n1840 S.t414 3.773
R1025 S.n1840 S.n1839 3.773
R1026 S.n1837 S.t515 3.773
R1027 S.n1837 S.n1836 3.773
R1028 S.n1823 S.n1822 3.773
R1029 S.n1823 S.t385 3.773
R1030 S.n1558 S.n1557 3.773
R1031 S.n1558 S.t360 3.773
R1032 S.n1569 S.t149 3.773
R1033 S.n1569 S.n1568 3.773
R1034 S.n1566 S.t849 3.773
R1035 S.n1566 S.n1565 3.773
R1036 S.n1561 S.n1560 3.773
R1037 S.n1561 S.t713 3.773
R1038 S.n1274 S.n1273 3.773
R1039 S.n1274 S.t97 3.773
R1040 S.n1294 S.t495 3.773
R1041 S.n1294 S.n1293 3.773
R1042 S.n1291 S.t584 3.773
R1043 S.n1291 S.n1290 3.773
R1044 S.n1277 S.n1276 3.773
R1045 S.n1277 S.t469 3.773
R1046 S.n1030 S.n1029 3.773
R1047 S.n1030 S.t950 3.773
R1048 S.n1041 S.t221 3.773
R1049 S.n1041 S.n1040 3.773
R1050 S.n1038 S.t960 3.773
R1051 S.n1038 S.n1037 3.773
R1052 S.n1033 S.n1032 3.773
R1053 S.n1033 S.t204 3.773
R1054 S.n739 S.n738 3.773
R1055 S.n739 S.t346 3.773
R1056 S.n759 S.t730 3.773
R1057 S.n759 S.n758 3.773
R1058 S.n756 S.t839 3.773
R1059 S.n756 S.n755 3.773
R1060 S.n742 S.n741 3.773
R1061 S.n742 S.t582 3.773
R1062 S.n380 S.n379 3.773
R1063 S.n380 S.t87 3.773
R1064 S.n391 S.t483 3.773
R1065 S.n391 S.n390 3.773
R1066 S.n388 S.t578 3.773
R1067 S.n388 S.n387 3.773
R1068 S.n383 S.n382 3.773
R1069 S.n383 S.t462 3.773
R1070 S.n363 S.n362 3.773
R1071 S.n363 S.t860 3.773
R1072 S.n374 S.t125 3.773
R1073 S.n374 S.n373 3.773
R1074 S.n371 S.t226 3.773
R1075 S.n371 S.n370 3.773
R1076 S.n366 S.n365 3.773
R1077 S.n366 S.t102 3.773
R1078 S.n67 S.t1124 3.773
R1079 S.n59 S.t768 3.773
R1080 S.n60 S.t555 3.773
R1081 S.n177 S.n176 3.773
R1082 S.n177 S.t436 3.773
R1083 S.n180 S.t814 3.773
R1084 S.n180 S.n179 3.773
R1085 S.n188 S.t912 3.773
R1086 S.n188 S.n187 3.773
R1087 S.n183 S.n182 3.773
R1088 S.n183 S.t791 3.773
R1089 S.n947 S.n946 3.773
R1090 S.n947 S.t885 3.773
R1091 S.n959 S.t157 3.773
R1092 S.n959 S.n958 3.773
R1093 S.n962 S.t250 3.773
R1094 S.n962 S.n961 3.773
R1095 S.n944 S.n943 3.773
R1096 S.n944 S.t1118 3.773
R1097 S.n987 S.t386 3.773
R1098 S.n988 S.t393 3.773
R1099 S.n968 S.t739 3.773
R1100 S.n146 S.t359 3.773
R1101 S.n147 S.t1110 3.773
R1102 S.n144 S.t388 3.773
R1103 S.n200 S.n199 3.773
R1104 S.n200 S.t247 3.773
R1105 S.n211 S.t626 3.773
R1106 S.n211 S.n210 3.773
R1107 S.n208 S.t743 3.773
R1108 S.n208 S.n207 3.773
R1109 S.n203 S.n202 3.773
R1110 S.n203 S.t608 3.773
R1111 S.n1532 S.t124 3.773
R1112 S.n1533 S.t605 3.773
R1113 S.n1512 S.t498 3.773
R1114 S.n1488 S.n1487 3.773
R1115 S.n1488 S.t973 3.773
R1116 S.n1503 S.t245 3.773
R1117 S.n1503 S.n1502 3.773
R1118 S.n1506 S.t354 3.773
R1119 S.n1506 S.n1505 3.773
R1120 S.n1491 S.n1490 3.773
R1121 S.n1491 S.t224 3.773
R1122 S.n994 S.n993 3.773
R1123 S.n994 S.t784 3.773
R1124 S.n1005 S.t1104 3.773
R1125 S.n1005 S.n1004 3.773
R1126 S.n1002 S.t734 3.773
R1127 S.n1002 S.n1001 3.773
R1128 S.n997 S.n996 3.773
R1129 S.n997 S.t1074 3.773
R1130 S.n680 S.n679 3.773
R1131 S.n680 S.t176 3.773
R1132 S.n700 S.t560 3.773
R1133 S.n700 S.n699 3.773
R1134 S.n697 S.t651 3.773
R1135 S.n697 S.n696 3.773
R1136 S.n683 S.n682 3.773
R1137 S.n683 S.t419 3.773
R1138 S.n347 S.n346 3.773
R1139 S.n347 S.t518 3.773
R1140 S.n358 S.t292 3.773
R1141 S.n358 S.n357 3.773
R1142 S.n355 S.t987 3.773
R1143 S.n355 S.n354 3.773
R1144 S.n350 S.n349 3.773
R1145 S.n350 S.t874 3.773
R1146 S.n330 S.n329 3.773
R1147 S.n330 S.t673 3.773
R1148 S.n341 S.t1000 3.773
R1149 S.n341 S.n340 3.773
R1150 S.n338 S.t1113 3.773
R1151 S.n338 S.n337 3.773
R1152 S.n333 S.n332 3.773
R1153 S.n333 S.t980 3.773
R1154 S.n54 S.t540 3.773
R1155 S.n34 S.t892 3.773
R1156 S.n646 S.t754 3.773
R1157 S.n648 S.t400 3.773
R1158 S.n650 S.t254 3.773
R1159 S.n486 S.n485 3.773
R1160 S.n486 S.t146 3.773
R1161 S.n495 S.t769 3.773
R1162 S.n495 S.n494 3.773
R1163 S.n498 S.t321 3.773
R1164 S.n498 S.n497 3.773
R1165 S.n489 S.n488 3.773
R1166 S.n489 S.t825 3.773
R1167 S.n1195 S.n1194 3.773
R1168 S.n1195 S.t403 3.773
R1169 S.n1204 S.t779 3.773
R1170 S.n1204 S.n1203 3.773
R1171 S.n1207 S.t664 3.773
R1172 S.n1207 S.n1206 3.773
R1173 S.n1198 S.n1197 3.773
R1174 S.n1198 S.t669 3.773
R1175 S.n966 S.n965 3.773
R1176 S.n966 S.t648 3.773
R1177 S.n1181 S.t1027 3.773
R1178 S.n1181 S.n1180 3.773
R1179 S.n1184 S.t1051 3.773
R1180 S.n1184 S.n1183 3.773
R1181 S.n1187 S.n1186 3.773
R1182 S.n1187 S.t568 3.773
R1183 S.n1738 S.n1737 3.773
R1184 S.n1738 S.t656 3.773
R1185 S.n1750 S.t1035 3.773
R1186 S.n1750 S.n1749 3.773
R1187 S.n1753 S.t946 3.773
R1188 S.n1753 S.n1752 3.773
R1189 S.n1741 S.n1740 3.773
R1190 S.n1741 S.t576 3.773
R1191 S.n1510 S.n1509 3.773
R1192 S.n1510 S.t668 3.773
R1193 S.n1723 S.t1048 3.773
R1194 S.n1723 S.n1722 3.773
R1195 S.n1726 S.t954 3.773
R1196 S.n1726 S.n1725 3.773
R1197 S.n1729 S.n1728 3.773
R1198 S.n1729 S.t590 3.773
R1199 S.n2067 S.n2066 3.773
R1200 S.n2067 S.t680 3.773
R1201 S.n2079 S.t1058 3.773
R1202 S.n2079 S.n2078 3.773
R1203 S.n2082 S.t969 3.773
R1204 S.n2082 S.n2081 3.773
R1205 S.n2070 S.n2069 3.773
R1206 S.n2070 S.t597 3.773
R1207 S.n2049 S.n2048 3.773
R1208 S.n2049 S.t688 3.773
R1209 S.n2052 S.t1071 3.773
R1210 S.n2052 S.n2051 3.773
R1211 S.n2055 S.t975 3.773
R1212 S.n2055 S.n2054 3.773
R1213 S.n2058 S.n2057 3.773
R1214 S.n2058 S.t606 3.773
R1215 S.n2593 S.n2592 3.773
R1216 S.n2593 S.t705 3.773
R1217 S.n2605 S.t1091 3.773
R1218 S.n2605 S.n2604 3.773
R1219 S.n2608 S.t985 3.773
R1220 S.n2608 S.n2607 3.773
R1221 S.n2596 S.n2595 3.773
R1222 S.n2596 S.t615 3.773
R1223 S.n2575 S.n2574 3.773
R1224 S.n2575 S.t720 3.773
R1225 S.n2578 S.t1102 3.773
R1226 S.n2578 S.n2577 3.773
R1227 S.n2581 S.t995 3.773
R1228 S.n2581 S.n2580 3.773
R1229 S.n2584 S.n2583 3.773
R1230 S.n2584 S.t622 3.773
R1231 S.n3097 S.n3096 3.773
R1232 S.n3097 S.t733 3.773
R1233 S.n3109 S.t47 3.773
R1234 S.n3109 S.n3108 3.773
R1235 S.n3112 S.t1008 3.773
R1236 S.n3112 S.n3111 3.773
R1237 S.n3100 S.n3099 3.773
R1238 S.n3100 S.t633 3.773
R1239 S.n3079 S.n3078 3.773
R1240 S.n3079 S.t1031 3.773
R1241 S.n3082 S.t249 3.773
R1242 S.n3082 S.n3081 3.773
R1243 S.n3085 S.t362 3.773
R1244 S.n3085 S.n3084 3.773
R1245 S.n3088 S.n3087 3.773
R1246 S.n3088 S.t229 3.773
R1247 S.n3774 S.n3773 3.773
R1248 S.n3774 S.t130 3.773
R1249 S.n3786 S.t521 3.773
R1250 S.n3786 S.n3785 3.773
R1251 S.n3789 S.t611 3.773
R1252 S.n3789 S.n3788 3.773
R1253 S.n3777 S.n3776 3.773
R1254 S.n3777 S.t581 3.773
R1255 S.n3570 S.n3569 3.773
R1256 S.n3570 S.t491 3.773
R1257 S.n3759 S.t869 3.773
R1258 S.n3759 S.n3758 3.773
R1259 S.n3762 S.t959 3.773
R1260 S.n3762 S.n3761 3.773
R1261 S.n3765 S.n3764 3.773
R1262 S.n3765 S.t846 3.773
R1263 S.n4060 S.n4059 3.773
R1264 S.n4060 S.t738 3.773
R1265 S.n4072 S.t1121 3.773
R1266 S.n4072 S.n4071 3.773
R1267 S.n4075 S.t110 3.773
R1268 S.n4075 S.n4074 3.773
R1269 S.n4063 S.n4062 3.773
R1270 S.n4063 S.t1092 3.773
R1271 S.n4042 S.n4041 3.773
R1272 S.n4042 S.t984 3.773
R1273 S.n4045 S.t253 3.773
R1274 S.n4045 S.n4044 3.773
R1275 S.n4048 S.t375 3.773
R1276 S.n4048 S.n4047 3.773
R1277 S.n4051 S.n4050 3.773
R1278 S.n4051 S.t239 3.773
R1279 S.n4502 S.n4501 3.773
R1280 S.n4502 S.t137 3.773
R1281 S.n4514 S.t528 3.773
R1282 S.n4514 S.n4513 3.773
R1283 S.n4517 S.t616 3.773
R1284 S.n4517 S.n4516 3.773
R1285 S.n4505 S.n4504 3.773
R1286 S.n4505 S.t509 3.773
R1287 S.n4484 S.n4483 3.773
R1288 S.n4484 S.t404 3.773
R1289 S.n4487 S.t783 3.773
R1290 S.n4487 S.n4486 3.773
R1291 S.n4490 S.t881 3.773
R1292 S.n4490 S.n4489 3.773
R1293 S.n4493 S.n4492 3.773
R1294 S.n4493 S.t758 3.773
R1295 S.n4891 S.n4890 3.773
R1296 S.n4891 S.t642 3.773
R1297 S.n4903 S.t1024 3.773
R1298 S.n4903 S.n4902 3.773
R1299 S.n4906 S.t1139 3.773
R1300 S.n4906 S.n4905 3.773
R1301 S.n4894 S.n4893 3.773
R1302 S.n4894 S.t1002 3.773
R1303 S.n5080 S.n5079 3.773
R1304 S.n5080 S.t910 3.773
R1305 S.n5090 S.t686 3.773
R1306 S.n5090 S.n5089 3.773
R1307 S.n5093 S.t273 3.773
R1308 S.n5093 S.n5092 3.773
R1309 S.n5083 S.n5082 3.773
R1310 S.n5083 S.t160 3.773
R1311 S.n5351 S.n5350 3.773
R1312 S.n5351 S.t569 3.773
R1313 S.n5362 S.t947 3.773
R1314 S.n5362 S.n5361 3.773
R1315 S.n5365 S.t1042 3.773
R1316 S.n5365 S.n5364 3.773
R1317 S.n5354 S.n5353 3.773
R1318 S.n5354 S.t928 3.773
R1319 S.n5267 S.t277 3.773
R1320 S.n5268 S.t527 3.773
R1321 S.n5265 S.t903 3.773
R1322 S.n1210 S.t644 3.773
R1323 S.n1212 S.t139 3.773
R1324 S.n1214 S.t990 3.773
R1325 S.n1167 S.n1166 3.773
R1326 S.n1167 S.t152 3.773
R1327 S.n1175 S.t264 3.773
R1328 S.n1175 S.n1174 3.773
R1329 S.n1178 S.t506 3.773
R1330 S.n1178 S.n1177 3.773
R1331 S.n1170 S.n1169 3.773
R1332 S.n1170 S.t697 3.773
R1333 S.n1761 S.n1760 3.773
R1334 S.n1761 S.t1003 3.773
R1335 S.n1765 S.t278 3.773
R1336 S.n1765 S.n1764 3.773
R1337 S.n1768 S.t187 3.773
R1338 S.n1768 S.n1767 3.773
R1339 S.n1758 S.n1757 3.773
R1340 S.n1758 S.t924 3.773
R1341 S.n5271 S.t676 3.773
R1342 S.n5272 S.t918 3.773
R1343 S.n5269 S.t190 3.773
R1344 S.n5373 S.n5372 3.773
R1345 S.n5373 S.t407 3.773
R1346 S.n5377 S.t787 3.773
R1347 S.n5377 S.n5376 3.773
R1348 S.n5380 S.t887 3.773
R1349 S.n5380 S.n5379 3.773
R1350 S.n5370 S.n5369 3.773
R1351 S.n5370 S.t762 3.773
R1352 S.n5101 S.n5100 3.773
R1353 S.n5101 S.t143 3.773
R1354 S.n5105 S.t534 3.773
R1355 S.n5105 S.n5104 3.773
R1356 S.n5108 S.t619 3.773
R1357 S.n5108 S.n5107 3.773
R1358 S.n5098 S.n5097 3.773
R1359 S.n5098 S.t512 3.773
R1360 S.n4914 S.n4913 3.773
R1361 S.n4914 S.t989 3.773
R1362 S.n4919 S.t260 3.773
R1363 S.n4919 S.n4918 3.773
R1364 S.n4922 S.t377 3.773
R1365 S.n4922 S.n4921 3.773
R1366 S.n4911 S.n4910 3.773
R1367 S.n4911 S.t241 3.773
R1368 S.n4539 S.n4538 3.773
R1369 S.n4539 S.t745 3.773
R1370 S.n4536 S.t1125 3.773
R1371 S.n4536 S.n4535 3.773
R1372 S.n4533 S.t115 3.773
R1373 S.n4533 S.n4532 3.773
R1374 S.n4530 S.n4529 3.773
R1375 S.n4530 S.t1099 3.773
R1376 S.n4525 S.n4524 3.773
R1377 S.n4525 S.t497 3.773
R1378 S.n4545 S.t871 3.773
R1379 S.n4545 S.n4544 3.773
R1380 S.n4548 S.t966 3.773
R1381 S.n4548 S.n4547 3.773
R1382 S.n4522 S.n4521 3.773
R1383 S.n4522 S.t852 3.773
R1384 S.n4097 S.n4096 3.773
R1385 S.n4097 S.t223 3.773
R1386 S.n4094 S.t604 3.773
R1387 S.n4094 S.n4093 3.773
R1388 S.n4091 S.t707 3.773
R1389 S.n4091 S.n4090 3.773
R1390 S.n4088 S.n4087 3.773
R1391 S.n4088 S.t588 3.773
R1392 S.n4083 S.n4082 3.773
R1393 S.n4083 S.t1073 3.773
R1394 S.n4103 S.t353 3.773
R1395 S.n4103 S.n4102 3.773
R1396 S.n4106 S.t468 3.773
R1397 S.n4106 S.n4105 3.773
R1398 S.n4080 S.n4079 3.773
R1399 S.n4080 S.t325 3.773
R1400 S.n3811 S.n3810 3.773
R1401 S.n3811 S.t882 3.773
R1402 S.n3808 S.t94 3.773
R1403 S.n3808 S.n3807 3.773
R1404 S.n3805 S.t199 3.773
R1405 S.n3805 S.n3804 3.773
R1406 S.n3802 S.n3801 3.773
R1407 S.n3802 S.t71 3.773
R1408 S.n3797 S.n3796 3.773
R1409 S.n3797 S.t1100 3.773
R1410 S.n3817 S.t915 3.773
R1411 S.n3817 S.n3816 3.773
R1412 S.n3820 S.t267 3.773
R1413 S.n3820 S.n3819 3.773
R1414 S.n3794 S.n3793 3.773
R1415 S.n3794 S.t64 3.773
R1416 S.n3134 S.n3133 3.773
R1417 S.n3134 S.t1085 3.773
R1418 S.n3131 S.t367 3.773
R1419 S.n3131 S.n3130 3.773
R1420 S.n3128 S.t252 3.773
R1421 S.n3128 S.n3127 3.773
R1422 S.n3125 S.n3124 3.773
R1423 S.n3125 S.t993 3.773
R1424 S.n3120 S.n3119 3.773
R1425 S.n3120 S.t1067 3.773
R1426 S.n3140 S.t349 3.773
R1427 S.n3140 S.n3139 3.773
R1428 S.n3143 S.t242 3.773
R1429 S.n3143 S.n3142 3.773
R1430 S.n3117 S.n3116 3.773
R1431 S.n3117 S.t983 3.773
R1432 S.n2630 S.n2629 3.773
R1433 S.n2630 S.t1055 3.773
R1434 S.n2627 S.t334 3.773
R1435 S.n2627 S.n2626 3.773
R1436 S.n2624 S.t238 3.773
R1437 S.n2624 S.n2623 3.773
R1438 S.n2621 S.n2620 3.773
R1439 S.n2621 S.t974 3.773
R1440 S.n2616 S.n2615 3.773
R1441 S.n2616 S.t1044 3.773
R1442 S.n2636 S.t319 3.773
R1443 S.n2636 S.n2635 3.773
R1444 S.n2639 S.t225 3.773
R1445 S.n2639 S.n2638 3.773
R1446 S.n2613 S.n2612 3.773
R1447 S.n2613 S.t967 3.773
R1448 S.n2104 S.n2103 3.773
R1449 S.n2104 S.t1033 3.773
R1450 S.n2101 S.t307 3.773
R1451 S.n2101 S.n2100 3.773
R1452 S.n2098 S.t215 3.773
R1453 S.n2098 S.n2097 3.773
R1454 S.n2095 S.n2094 3.773
R1455 S.n2095 S.t951 3.773
R1456 S.n2090 S.n2089 3.773
R1457 S.n2090 S.t1025 3.773
R1458 S.n2110 S.t298 3.773
R1459 S.n2110 S.n2109 3.773
R1460 S.n2113 S.t208 3.773
R1461 S.n2113 S.n2112 3.773
R1462 S.n2087 S.n2086 3.773
R1463 S.n2087 S.t943 3.773
R1464 S.n1693 S.n1692 3.773
R1465 S.n1693 S.t1015 3.773
R1466 S.n1697 S.t287 3.773
R1467 S.n1697 S.n1696 3.773
R1468 S.n1700 S.t195 3.773
R1469 S.n1700 S.n1699 3.773
R1470 S.n1690 S.n1689 3.773
R1471 S.n1690 S.t935 3.773
R1472 S.n1771 S.t649 3.773
R1473 S.n1773 S.t234 3.773
R1474 S.n1775 S.t111 3.773
R1475 S.n1705 S.n1704 3.773
R1476 S.n1705 S.t43 3.773
R1477 S.n1717 S.t631 3.773
R1478 S.n1717 S.n1716 3.773
R1479 S.n1720 S.t86 3.773
R1480 S.n1720 S.n1719 3.773
R1481 S.n1708 S.n1707 3.773
R1482 S.n1708 S.t587 3.773
R1483 S.n2121 S.n2120 3.773
R1484 S.n2121 S.t261 3.773
R1485 S.n2315 S.t643 3.773
R1486 S.n2315 S.n2314 3.773
R1487 S.n2318 S.t556 3.773
R1488 S.n2318 S.n2317 3.773
R1489 S.n2118 S.n2117 3.773
R1490 S.n2118 S.t184 3.773
R1491 S.n5275 S.t524 3.773
R1492 S.n5276 S.t752 3.773
R1493 S.n5273 S.t1131 3.773
R1494 S.n5388 S.n5387 3.773
R1495 S.n5388 S.t749 3.773
R1496 S.n5392 S.t1127 3.773
R1497 S.n5392 S.n5391 3.773
R1498 S.n5395 S.t120 3.773
R1499 S.n5395 S.n5394 3.773
R1500 S.n5385 S.n5384 3.773
R1501 S.n5385 S.t1103 3.773
R1502 S.n5116 S.n5115 3.773
R1503 S.n5116 S.t504 3.773
R1504 S.n5121 S.t876 3.773
R1505 S.n5121 S.n5120 3.773
R1506 S.n5124 S.t970 3.773
R1507 S.n5124 S.n5123 3.773
R1508 S.n5113 S.n5112 3.773
R1509 S.n5113 S.t855 3.773
R1510 S.n4930 S.n4929 3.773
R1511 S.n4930 S.t230 3.773
R1512 S.n4934 S.t610 3.773
R1513 S.n4934 S.n4933 3.773
R1514 S.n4937 S.t716 3.773
R1515 S.n4937 S.n4936 3.773
R1516 S.n4927 S.n4926 3.773
R1517 S.n4927 S.t593 3.773
R1518 S.n4697 S.n4696 3.773
R1519 S.n4697 S.t1081 3.773
R1520 S.n4702 S.t363 3.773
R1521 S.n4702 S.n4701 3.773
R1522 S.n4705 S.t471 3.773
R1523 S.n4705 S.n4704 3.773
R1524 S.n4694 S.n4693 3.773
R1525 S.n4694 S.t328 3.773
R1526 S.n4556 S.n4555 3.773
R1527 S.n4556 S.t834 3.773
R1528 S.n4560 S.t98 3.773
R1529 S.n4560 S.n4559 3.773
R1530 S.n4563 S.t207 3.773
R1531 S.n4563 S.n4562 3.773
R1532 S.n4553 S.n4552 3.773
R1533 S.n4553 S.t75 3.773
R1534 S.n4267 S.n4266 3.773
R1535 S.n4267 S.t620 3.773
R1536 S.n4272 S.t949 3.773
R1537 S.n4272 S.n4271 3.773
R1538 S.n4275 S.t1049 3.773
R1539 S.n4275 S.n4274 3.773
R1540 S.n4264 S.n4263 3.773
R1541 S.n4264 S.t933 3.773
R1542 S.n4114 S.n4113 3.773
R1543 S.n4114 S.t535 3.773
R1544 S.n4118 S.t759 3.773
R1545 S.n4118 S.n4117 3.773
R1546 S.n4121 S.t816 3.773
R1547 S.n4121 S.n4120 3.773
R1548 S.n4111 S.n4110 3.773
R1549 S.n4111 S.t450 3.773
R1550 S.n3681 S.n3680 3.773
R1551 S.n3681 S.t525 3.773
R1552 S.n3686 S.t900 3.773
R1553 S.n3686 S.n3685 3.773
R1554 S.n3689 S.t804 3.773
R1555 S.n3689 S.n3688 3.773
R1556 S.n3678 S.n3677 3.773
R1557 S.n3678 S.t439 3.773
R1558 S.n3828 S.n3827 3.773
R1559 S.n3828 S.t330 3.773
R1560 S.n3832 S.t717 3.773
R1561 S.n3832 S.n3831 3.773
R1562 S.n3835 S.t614 3.773
R1563 S.n3835 S.n3834 3.773
R1564 S.n3825 S.n3824 3.773
R1565 S.n3825 S.t428 3.773
R1566 S.n3313 S.n3312 3.773
R1567 S.n3313 S.t316 3.773
R1568 S.n3318 S.t700 3.773
R1569 S.n3318 S.n3317 3.773
R1570 S.n3321 S.t603 3.773
R1571 S.n3321 S.n3320 3.773
R1572 S.n3310 S.n3309 3.773
R1573 S.n3310 S.t236 3.773
R1574 S.n3151 S.n3150 3.773
R1575 S.n3151 S.t306 3.773
R1576 S.n3155 S.t687 3.773
R1577 S.n3155 S.n3154 3.773
R1578 S.n3158 S.t595 3.773
R1579 S.n3158 S.n3157 3.773
R1580 S.n3148 S.n3147 3.773
R1581 S.n3148 S.t222 3.773
R1582 S.n2814 S.n2813 3.773
R1583 S.n2814 S.t297 3.773
R1584 S.n2819 S.t677 3.773
R1585 S.n2819 S.n2818 3.773
R1586 S.n2822 S.t586 3.773
R1587 S.n2822 S.n2821 3.773
R1588 S.n2811 S.n2810 3.773
R1589 S.n2811 S.t213 3.773
R1590 S.n2647 S.n2646 3.773
R1591 S.n2647 S.t284 3.773
R1592 S.n2651 S.t663 3.773
R1593 S.n2651 S.n2650 3.773
R1594 S.n2654 S.t574 3.773
R1595 S.n2654 S.n2653 3.773
R1596 S.n2644 S.n2643 3.773
R1597 S.n2644 S.t206 3.773
R1598 S.n2310 S.n2309 3.773
R1599 S.n2310 S.t275 3.773
R1600 S.n2307 S.t654 3.773
R1601 S.n2307 S.n2306 3.773
R1602 S.n2304 S.t565 3.773
R1603 S.n2304 S.n2303 3.773
R1604 S.n2126 S.n2125 3.773
R1605 S.n2126 S.t192 3.773
R1606 S.n2321 S.t566 3.773
R1607 S.n2323 S.t1095 3.773
R1608 S.n2325 S.t968 3.773
R1609 S.n2286 S.n2285 3.773
R1610 S.n2286 S.t1062 3.773
R1611 S.n2298 S.t1001 3.773
R1612 S.n2298 S.n2297 3.773
R1613 S.n2301 S.t1070 3.773
R1614 S.n2301 S.n2300 3.773
R1615 S.n2289 S.n2288 3.773
R1616 S.n2289 S.t476 3.773
R1617 S.n2662 S.n2661 3.773
R1618 S.n2662 S.t627 3.773
R1619 S.n2856 S.t1013 3.773
R1620 S.n2856 S.n2855 3.773
R1621 S.n2859 S.t920 3.773
R1622 S.n2859 S.n2858 3.773
R1623 S.n2659 S.n2658 3.773
R1624 S.n2659 S.t553 3.773
R1625 S.n5279 S.t866 3.773
R1626 S.n5280 S.t1093 3.773
R1627 S.n5277 S.t372 3.773
R1628 S.n5403 S.n5402 3.773
R1629 S.n5403 S.t1087 3.773
R1630 S.n5407 S.t368 3.773
R1631 S.n5407 S.n5406 3.773
R1632 S.n5410 S.t477 3.773
R1633 S.n5410 S.n5409 3.773
R1634 S.n5400 S.n5399 3.773
R1635 S.n5400 S.t332 3.773
R1636 S.n5132 S.n5131 3.773
R1637 S.n5132 S.t838 3.773
R1638 S.n5137 S.t106 3.773
R1639 S.n5137 S.n5136 3.773
R1640 S.n5140 S.t210 3.773
R1641 S.n5140 S.n5139 3.773
R1642 S.n5129 S.n5128 3.773
R1643 S.n5129 S.t81 3.773
R1644 S.n4945 S.n4944 3.773
R1645 S.n4945 S.t577 3.773
R1646 S.n4949 S.t957 3.773
R1647 S.n4949 S.n4948 3.773
R1648 S.n4952 S.t1052 3.773
R1649 S.n4952 S.n4951 3.773
R1650 S.n4942 S.n4941 3.773
R1651 S.n4942 S.t938 3.773
R1652 S.n4713 S.n4712 3.773
R1653 S.n4713 S.t384 3.773
R1654 S.n4718 S.t694 3.773
R1655 S.n4718 S.n4717 3.773
R1656 S.n4721 S.t813 3.773
R1657 S.n4721 S.n4720 3.773
R1658 S.n4710 S.n4709 3.773
R1659 S.n4710 S.t672 3.773
R1660 S.n4571 S.n4570 3.773
R1661 S.n4571 S.t896 3.773
R1662 S.n4575 S.t514 3.773
R1663 S.n4575 S.n4574 3.773
R1664 S.n4578 S.t58 3.773
R1665 S.n4578 S.n4577 3.773
R1666 S.n4568 S.n4567 3.773
R1667 S.n4568 S.t812 3.773
R1668 S.n4283 S.n4282 3.773
R1669 S.n4283 S.t889 3.773
R1670 S.n4288 S.t161 3.773
R1671 S.n4288 S.n4287 3.773
R1672 S.n4291 S.t46 3.773
R1673 S.n4291 S.n4290 3.773
R1674 S.n4280 S.n4279 3.773
R1675 S.n4280 S.t798 3.773
R1676 S.n4129 S.n4128 3.773
R1677 S.n4129 S.t878 3.773
R1678 S.n4133 S.t147 3.773
R1679 S.n4133 S.n4132 3.773
R1680 S.n4136 S.t28 3.773
R1681 S.n4136 S.n4135 3.773
R1682 S.n4126 S.n4125 3.773
R1683 S.n4126 S.t793 3.773
R1684 S.n3697 S.n3696 3.773
R1685 S.n3697 S.t868 3.773
R1686 S.n3702 S.t133 3.773
R1687 S.n3702 S.n3701 3.773
R1688 S.n3705 S.t11 3.773
R1689 S.n3705 S.n3704 3.773
R1690 S.n3694 S.n3693 3.773
R1691 S.n3694 S.t778 3.773
R1692 S.n3843 S.n3842 3.773
R1693 S.n3843 S.t674 3.773
R1694 S.n3847 S.t1053 3.773
R1695 S.n3847 S.n3846 3.773
R1696 S.n3850 S.t965 3.773
R1697 S.n3850 S.n3849 3.773
R1698 S.n3840 S.n3839 3.773
R1699 S.n3840 S.t767 3.773
R1700 S.n3329 S.n3328 3.773
R1701 S.n3329 S.t662 3.773
R1702 S.n3334 S.t1041 3.773
R1703 S.n3334 S.n3333 3.773
R1704 S.n3337 S.t948 3.773
R1705 S.n3337 S.n3336 3.773
R1706 S.n3326 S.n3325 3.773
R1707 S.n3326 S.t583 3.773
R1708 S.n3166 S.n3165 3.773
R1709 S.n3166 S.t653 3.773
R1710 S.n3170 S.t1032 3.773
R1711 S.n3170 S.n3169 3.773
R1712 S.n3173 S.t941 3.773
R1713 S.n3173 S.n3172 3.773
R1714 S.n3163 S.n3162 3.773
R1715 S.n3163 S.t572 3.773
R1716 S.n2851 S.n2850 3.773
R1717 S.n2851 S.t640 3.773
R1718 S.n2848 S.t1022 3.773
R1719 S.n2848 S.n2847 3.773
R1720 S.n2845 S.t932 3.773
R1721 S.n2845 S.n2844 3.773
R1722 S.n2667 S.n2666 3.773
R1723 S.n2667 S.t564 3.773
R1724 S.n2862 S.t480 3.773
R1725 S.n2864 S.t851 3.773
R1726 S.n2866 S.t715 3.773
R1727 S.n2827 S.n2826 3.773
R1728 S.n2827 S.t972 3.773
R1729 S.n2839 S.t258 3.773
R1730 S.n2839 S.n2838 3.773
R1731 S.n2842 S.t952 3.773
R1732 S.n2842 S.n2841 3.773
R1733 S.n2830 S.n2829 3.773
R1734 S.n2830 S.t337 3.773
R1735 S.n3181 S.n3180 3.773
R1736 S.n3181 S.t997 3.773
R1737 S.n3371 S.t272 3.773
R1738 S.n3371 S.n3370 3.773
R1739 S.n3374 S.t182 3.773
R1740 S.n3374 S.n3373 3.773
R1741 S.n3178 S.n3177 3.773
R1742 S.n3178 S.t919 3.773
R1743 S.n5283 S.t92 3.773
R1744 S.n5284 S.t322 3.773
R1745 S.n5281 S.t708 3.773
R1746 S.n5418 S.n5417 3.773
R1747 S.n5418 S.t317 3.773
R1748 S.n5422 S.t698 3.773
R1749 S.n5422 S.n5421 3.773
R1750 S.n5425 S.t822 3.773
R1751 S.n5425 S.n5424 3.773
R1752 S.n5415 S.n5414 3.773
R1753 S.n5415 S.t679 3.773
R1754 S.n5148 S.n5147 3.773
R1755 S.n5148 S.t121 3.773
R1756 S.n5153 S.t461 3.773
R1757 S.n5153 S.n5152 3.773
R1758 S.n5156 S.t559 3.773
R1759 S.n5156 S.n5155 3.773
R1760 S.n5145 S.n5144 3.773
R1761 S.n5145 S.t444 3.773
R1762 S.n4960 S.n4959 3.773
R1763 S.n4960 S.t158 3.773
R1764 S.n4964 S.t243 3.773
R1765 S.n4964 S.n4963 3.773
R1766 S.n4967 S.t448 3.773
R1767 S.n4967 S.n4966 3.773
R1768 S.n4957 S.n4956 3.773
R1769 S.n4957 S.t57 3.773
R1770 S.n4729 S.n4728 3.773
R1771 S.n4729 S.t144 3.773
R1772 S.n4734 S.t533 3.773
R1773 S.n4734 S.n4733 3.773
R1774 S.n4737 S.t434 3.773
R1775 S.n4737 S.n4736 3.773
R1776 S.n4726 S.n4725 3.773
R1777 S.n4726 S.t39 3.773
R1778 S.n4586 S.n4585 3.773
R1779 S.n4586 S.t132 3.773
R1780 S.n4590 S.t522 3.773
R1781 S.n4590 S.n4589 3.773
R1782 S.n4593 S.t424 3.773
R1783 S.n4593 S.n4592 3.773
R1784 S.n4583 S.n4582 3.773
R1785 S.n4583 S.t20 3.773
R1786 S.n4299 S.n4298 3.773
R1787 S.n4299 S.t118 3.773
R1788 S.n4304 S.t513 3.773
R1789 S.n4304 S.n4303 3.773
R1790 S.n4307 S.t415 3.773
R1791 S.n4307 S.n4306 3.773
R1792 S.n4296 S.n4295 3.773
R1793 S.n4296 S.t5 3.773
R1794 S.n4144 S.n4143 3.773
R1795 S.n4144 S.t109 3.773
R1796 S.n4148 S.t505 3.773
R1797 S.n4148 S.n4147 3.773
R1798 S.n4151 S.t399 3.773
R1799 S.n4151 S.n4150 3.773
R1800 S.n4141 S.n4140 3.773
R1801 S.n4141 S.t1133 3.773
R1802 S.n3713 S.n3712 3.773
R1803 S.n3713 S.t93 3.773
R1804 S.n3718 S.t489 3.773
R1805 S.n3718 S.n3717 3.773
R1806 S.n3721 S.t387 3.773
R1807 S.n3721 S.n3720 3.773
R1808 S.n3710 S.n3709 3.773
R1809 S.n3710 S.t1122 3.773
R1810 S.n3858 S.n3857 3.773
R1811 S.n3858 S.t1020 3.773
R1812 S.n3862 S.t293 3.773
R1813 S.n3862 S.n3861 3.773
R1814 S.n3865 S.t202 3.773
R1815 S.n3865 S.n3864 3.773
R1816 S.n3855 S.n3854 3.773
R1817 S.n3855 S.t1108 3.773
R1818 S.n3366 S.n3365 3.773
R1819 S.n3366 S.t1011 3.773
R1820 S.n3363 S.t283 3.773
R1821 S.n3363 S.n3362 3.773
R1822 S.n3360 S.t191 3.773
R1823 S.n3360 S.n3359 3.773
R1824 S.n3186 S.n3185 3.773
R1825 S.n3186 S.t929 3.773
R1826 S.n3377 S.t383 3.773
R1827 S.n3379 S.t592 3.773
R1828 S.n3381 S.t475 3.773
R1829 S.n3342 S.n3341 3.773
R1830 S.n3342 S.t888 3.773
R1831 S.n3357 S.t624 3.773
R1832 S.n3357 S.n3356 3.773
R1833 S.n3345 S.t843 3.773
R1834 S.n3345 S.n3344 3.773
R1835 S.n3348 S.n3347 3.773
R1836 S.n3348 S.t218 3.773
R1837 S.n3873 S.n3872 3.773
R1838 S.n3873 S.t255 3.773
R1839 S.n3877 S.t637 3.773
R1840 S.n3877 S.n3876 3.773
R1841 S.n3880 S.t549 3.773
R1842 S.n3880 S.n3879 3.773
R1843 S.n3870 S.n3869 3.773
R1844 S.n3870 S.t343 3.773
R1845 S.n5287 S.t454 3.773
R1846 S.n5288 S.t665 3.773
R1847 S.n5285 S.t1046 3.773
R1848 S.n5433 S.n5432 3.773
R1849 S.n5433 S.t531 3.773
R1850 S.n5437 S.t1111 3.773
R1851 S.n5437 S.n5436 3.773
R1852 S.n5440 S.t809 3.773
R1853 S.n5440 S.n5439 3.773
R1854 S.n5430 S.n5429 3.773
R1855 S.n5430 S.t446 3.773
R1856 S.n5164 S.n5163 3.773
R1857 S.n5164 S.t519 3.773
R1858 S.n5169 S.t894 3.773
R1859 S.n5169 S.n5168 3.773
R1860 S.n5172 S.t796 3.773
R1861 S.n5172 S.n5171 3.773
R1862 S.n5161 S.n5160 3.773
R1863 S.n5161 S.t431 3.773
R1864 S.n4975 S.n4974 3.773
R1865 S.n4975 S.t511 3.773
R1866 S.n4979 S.t886 3.773
R1867 S.n4979 S.n4978 3.773
R1868 S.n4982 S.t789 3.773
R1869 S.n4982 S.n4981 3.773
R1870 S.n4972 S.n4971 3.773
R1871 S.n4972 S.t423 3.773
R1872 S.n4745 S.n4744 3.773
R1873 S.n4745 S.t502 3.773
R1874 S.n4750 S.t877 3.773
R1875 S.n4750 S.n4749 3.773
R1876 S.n4753 S.t775 3.773
R1877 S.n4753 S.n4752 3.773
R1878 S.n4742 S.n4741 3.773
R1879 S.n4742 S.t411 3.773
R1880 S.n4601 S.n4600 3.773
R1881 S.n4601 S.t486 3.773
R1882 S.n4605 S.t864 3.773
R1883 S.n4605 S.n4604 3.773
R1884 S.n4608 S.t764 3.773
R1885 S.n4608 S.n4607 3.773
R1886 S.n4598 S.n4597 3.773
R1887 S.n4598 S.t395 3.773
R1888 S.n4315 S.n4314 3.773
R1889 S.n4315 S.t479 3.773
R1890 S.n4320 S.t856 3.773
R1891 S.n4320 S.n4319 3.773
R1892 S.n4323 S.t753 3.773
R1893 S.n4323 S.n4322 3.773
R1894 S.n4312 S.n4311 3.773
R1895 S.n4312 S.t382 3.773
R1896 S.n4159 S.n4158 3.773
R1897 S.n4159 S.t467 3.773
R1898 S.n4163 S.t845 3.773
R1899 S.n4163 S.n4162 3.773
R1900 S.n4166 S.t740 3.773
R1901 S.n4166 S.n4165 3.773
R1902 S.n4156 S.n4155 3.773
R1903 S.n4156 S.t373 3.773
R1904 S.n3729 S.n3728 3.773
R1905 S.n3729 S.t456 3.773
R1906 S.n3733 S.t833 3.773
R1907 S.n3733 S.n3732 3.773
R1908 S.n3736 S.t726 3.773
R1909 S.n3736 S.n3735 3.773
R1910 S.n3726 S.n3725 3.773
R1911 S.n3726 S.t356 3.773
R1912 S.n3883 S.t276 3.773
R1913 S.n3885 S.t331 3.773
R1914 S.n3887 S.t299 3.773
R1915 S.n3741 S.n3740 3.773
R1916 S.n3741 S.t493 3.773
R1917 S.n3753 S.t54 3.773
R1918 S.n3753 S.n3752 3.773
R1919 S.n3756 S.t1096 3.773
R1920 S.n3756 S.n3755 3.773
R1921 S.n3744 S.n3743 3.773
R1922 S.n3744 S.t490 3.773
R1923 S.n4174 S.n4173 3.773
R1924 S.n4174 S.t805 3.773
R1925 S.n4357 S.t69 3.773
R1926 S.n4357 S.n4356 3.773
R1927 S.n4360 S.t1077 3.773
R1928 S.n4360 S.n4359 3.773
R1929 S.n4171 S.n4170 3.773
R1930 S.n4171 S.t711 3.773
R1931 S.n5291 S.t744 3.773
R1932 S.n5292 S.t211 3.773
R1933 S.n5289 S.t345 3.773
R1934 S.n5448 S.n5447 3.773
R1935 S.n5448 S.t875 3.773
R1936 S.n5452 S.t142 3.773
R1937 S.n5452 S.n5451 3.773
R1938 S.n5455 S.t18 3.773
R1939 S.n5455 S.n5454 3.773
R1940 S.n5445 S.n5444 3.773
R1941 S.n5445 S.t786 3.773
R1942 S.n5180 S.n5179 3.773
R1943 S.n5180 S.t861 3.773
R1944 S.n5185 S.t126 3.773
R1945 S.n5185 S.n5184 3.773
R1946 S.n5188 S.t1 3.773
R1947 S.n5188 S.n5187 3.773
R1948 S.n5177 S.n5176 3.773
R1949 S.n5177 S.t773 3.773
R1950 S.n4990 S.n4989 3.773
R1951 S.n4990 S.t853 3.773
R1952 S.n4994 S.t116 3.773
R1953 S.n4994 S.n4993 3.773
R1954 S.n4997 S.t1129 3.773
R1955 S.n4997 S.n4996 3.773
R1956 S.n4987 S.n4986 3.773
R1957 S.n4987 S.t763 3.773
R1958 S.n4761 S.n4760 3.773
R1959 S.n4761 S.t842 3.773
R1960 S.n4766 S.t104 3.773
R1961 S.n4766 S.n4765 3.773
R1962 S.n4769 S.t1120 3.773
R1963 S.n4769 S.n4768 3.773
R1964 S.n4758 S.n4757 3.773
R1965 S.n4758 S.t751 3.773
R1966 S.n4616 S.n4615 3.773
R1967 S.n4616 S.t830 3.773
R1968 S.n4620 S.t91 3.773
R1969 S.n4620 S.n4619 3.773
R1970 S.n4623 S.t1106 3.773
R1971 S.n4623 S.n4622 3.773
R1972 S.n4613 S.n4612 3.773
R1973 S.n4613 S.t736 3.773
R1974 S.n4352 S.n4351 3.773
R1975 S.n4352 S.t820 3.773
R1976 S.n4349 S.t82 3.773
R1977 S.n4349 S.n4348 3.773
R1978 S.n4346 S.t1094 3.773
R1979 S.n4346 S.n4345 3.773
R1980 S.n4179 S.n4178 3.773
R1981 S.n4179 S.t723 3.773
R1982 S.n4363 S.t982 3.773
R1983 S.n4365 S.t183 3.773
R1984 S.n4367 S.t38 3.773
R1985 S.n4328 S.n4327 3.773
R1986 S.n4328 S.t396 3.773
R1987 S.n4340 S.t443 3.773
R1988 S.n4340 S.n4339 3.773
R1989 S.n4343 S.t971 3.773
R1990 S.n4343 S.n4342 3.773
R1991 S.n4331 S.n4330 3.773
R1992 S.n4331 S.t357 3.773
R1993 S.n4631 S.n4630 3.773
R1994 S.n4631 S.t51 3.773
R1995 S.n4806 S.t455 3.773
R1996 S.n4806 S.n4805 3.773
R1997 S.n4809 S.t340 3.773
R1998 S.n4809 S.n4808 3.773
R1999 S.n4628 S.n4627 3.773
R2000 S.n4628 S.t1072 3.773
R2001 S.n5295 S.t1080 3.773
R2002 S.n5296 S.t561 3.773
R2003 S.n5293 S.t939 3.773
R2004 S.n5463 S.n5462 3.773
R2005 S.n5463 S.t101 3.773
R2006 S.n5467 S.t499 3.773
R2007 S.n5467 S.n5466 3.773
R2008 S.n5470 S.t394 3.773
R2009 S.n5470 S.n5469 3.773
R2010 S.n5460 S.n5459 3.773
R2011 S.n5460 S.t1128 3.773
R2012 S.n5196 S.n5195 3.773
R2013 S.n5196 S.t88 3.773
R2014 S.n5201 S.t484 3.773
R2015 S.n5201 S.n5200 3.773
R2016 S.n5204 S.t379 3.773
R2017 S.n5204 S.n5203 3.773
R2018 S.n5193 S.n5192 3.773
R2019 S.n5193 S.t1116 3.773
R2020 S.n5005 S.n5004 3.773
R2021 S.n5005 S.t80 3.773
R2022 S.n5009 S.t474 3.773
R2023 S.n5009 S.n5008 3.773
R2024 S.n5012 S.t370 3.773
R2025 S.n5012 S.n5011 3.773
R2026 S.n5002 S.n5001 3.773
R2027 S.n5002 S.t1101 3.773
R2028 S.n4801 S.n4800 3.773
R2029 S.n4801 S.t68 3.773
R2030 S.n4798 S.t465 3.773
R2031 S.n4798 S.n4797 3.773
R2032 S.n4795 S.t351 3.773
R2033 S.n4795 S.n4794 3.773
R2034 S.n4636 S.n4635 3.773
R2035 S.n4636 S.t1090 3.773
R2036 S.n4812 S.t899 3.773
R2037 S.n4814 S.t1029 3.773
R2038 S.n4816 S.t914 3.773
R2039 S.n4772 S.n4771 3.773
R2040 S.n4772 S.t288 3.773
R2041 S.n4789 S.t803 3.773
R2042 S.n4789 S.n4788 3.773
R2043 S.n4792 S.t858 3.773
R2044 S.n4792 S.n4791 3.773
R2045 S.n4775 S.n4774 3.773
R2046 S.n4775 S.t232 3.773
R2047 S.n5223 S.n5222 3.773
R2048 S.n5223 S.t438 3.773
R2049 S.n5232 S.t819 3.773
R2050 S.n5232 S.n5231 3.773
R2051 S.n5235 S.t706 3.773
R2052 S.n5235 S.n5234 3.773
R2053 S.n5226 S.n5225 3.773
R2054 S.n5226 S.t336 3.773
R2055 S.n5299 S.t312 3.773
R2056 S.n5300 S.t906 3.773
R2057 S.n5297 S.t178 3.773
R2058 S.n5477 S.n5476 3.773
R2059 S.n5477 S.t460 3.773
R2060 S.n5485 S.t837 3.773
R2061 S.n5485 S.n5484 3.773
R2062 S.n5488 S.t732 3.773
R2063 S.n5488 S.n5487 3.773
R2064 S.n5480 S.n5479 3.773
R2065 S.n5480 S.t366 3.773
R2066 S.n5021 S.n5020 3.773
R2067 S.n5021 S.t453 3.773
R2068 S.n5207 S.t828 3.773
R2069 S.n5207 S.n5206 3.773
R2070 S.n5210 S.t719 3.773
R2071 S.n5210 S.n5209 3.773
R2072 S.n5213 S.n5212 3.773
R2073 S.n5213 S.t348 3.773
R2074 S.n5264 S.t1006 3.773
R2075 S.n5261 S.t496 3.773
R2076 S.n5262 S.t872 3.773
R2077 S.n5491 S.t703 3.773
R2078 S.n5493 S.t541 3.773
R2079 S.n5495 S.t421 3.773
R2080 S.n315 S.n313 2.808
R2081 S.n977 S.n975 2.808
R2082 S.n1523 S.n1521 2.808
R2083 S.n2137 S.n2135 2.808
R2084 S.n2680 S.n2678 2.808
R2085 S.n3197 S.n3195 2.808
R2086 S.n3583 S.n3581 2.808
R2087 S.n4187 S.n4185 2.808
R2088 S.n38 S.n37 2.645
R2089 S.n309 S.n308 2.645
R2090 S.n971 S.n970 2.645
R2091 S.n1517 S.n1516 2.645
R2092 S.n2131 S.n2130 2.645
R2093 S.n2674 S.n2673 2.645
R2094 S.n3191 S.n3190 2.645
R2095 S.n3577 S.n3576 2.645
R2096 S.n4829 S.n4828 0.21
R2097 S.n664 S.n663 0.172
R2098 S.n40 S.n36 0.164
R2099 S.n5499 S.n5308 0.143
R2100 S.n1437 S.n1436 0.133
R2101 S.n1201 S.n1200 0.133
R2102 S.n164 S.n156 0.123
R2103 S.n62 S.n61 0.123
R2104 S.n30 S.n29 0.12
R2105 S.n20 S.n19 0.12
R2106 S.n5508 S.n1230 0.114
R2107 S.n5509 S.n668 0.111
R2108 S.n5507 S.n1808 0.111
R2109 S.n5506 S.n2358 0.111
R2110 S.n5505 S.n2899 0.111
R2111 S.n5504 S.n3414 0.111
R2112 S.n5503 S.n3920 0.111
R2113 S.n5502 S.n4398 0.111
R2114 S.n5501 S.n4831 0.111
R2115 S.n5499 S.n5498 0.11
R2116 S.n5500 S.n5260 0.11
R2117 S.n4664 S.n4662 0.109
R2118 S.n4233 S.n4231 0.109
R2119 S.n3647 S.n3645 0.109
R2120 S.n3279 S.n3277 0.109
R2121 S.n2780 S.n2778 0.109
R2122 S.n2255 S.n2253 0.109
R2123 S.n1659 S.n1657 0.109
R2124 S.n1713 S.n1710 0.106
R2125 S.n2294 S.n2291 0.106
R2126 S.n2835 S.n2832 0.106
R2127 S.n3353 S.n3350 0.106
R2128 S.n3749 S.n3746 0.106
R2129 S.n4336 S.n4333 0.106
R2130 S.n5069 S.n5064 0.106
R2131 S.n1397 S.n1396 0.097
R2132 S.n1942 S.n1941 0.097
R2133 S.n2463 S.n2462 0.097
R2134 S.n2972 S.n2971 0.097
R2135 S.n3458 S.n3457 0.097
R2136 S.n3932 S.n3931 0.097
R2137 S.n4463 S.n4462 0.097
R2138 S.n876 S.n875 0.097
R2139 S.n904 S.n903 0.097
R2140 S.n5253 S.n5252 0.095
R2141 S.n5026 S.n5025 0.093
R2142 S.n833 S.n832 0.087
R2143 S.n665 S.n662 0.081
R2144 S.n1224 S.n1221 0.081
R2145 S.n1787 S.n1784 0.081
R2146 S.n2337 S.n2334 0.081
R2147 S.n2878 S.n2875 0.081
R2148 S.n3393 S.n3390 0.081
R2149 S.n3899 S.n3896 0.081
R2150 S.n4377 S.n4374 0.081
R2151 S.n4458 S.n4457 0.08
R2152 S.n3927 S.n3926 0.08
R2153 S.n3453 S.n3452 0.08
R2154 S.n2967 S.n2966 0.08
R2155 S.n2458 S.n2457 0.08
R2156 S.n1937 S.n1936 0.08
R2157 S.n1392 S.n1391 0.08
R2158 S.n906 S.n905 0.08
R2159 S.n878 S.n877 0.08
R2160 S.n1801 S.n1800 0.079
R2161 S.n2351 S.n2350 0.079
R2162 S.n2892 S.n2891 0.079
R2163 S.n3407 S.n3406 0.079
R2164 S.n3913 S.n3912 0.079
R2165 S.n4391 S.n4390 0.079
R2166 S.n1106 S.n1105 0.077
R2167 S.n1629 S.n1628 0.077
R2168 S.n2225 S.n2224 0.077
R2169 S.n2750 S.n2749 0.077
R2170 S.n3249 S.n3248 0.077
R2171 S.n3617 S.n3616 0.077
R2172 S.n4203 S.n4202 0.077
R2173 S.n438 S.n437 0.077
R2174 S.n457 S.n456 0.077
R2175 S.n1804 S.n1803 0.075
R2176 S.n2354 S.n2353 0.075
R2177 S.n2895 S.n2894 0.075
R2178 S.n3410 S.n3409 0.075
R2179 S.n3916 S.n3915 0.075
R2180 S.n4394 S.n4393 0.075
R2181 S.n4192 S.n4191 0.074
R2182 S.n3588 S.n3587 0.074
R2183 S.n3202 S.n3201 0.074
R2184 S.n2685 S.n2684 0.074
R2185 S.n2142 S.n2141 0.074
R2186 S.n1528 S.n1527 0.074
R2187 S.n982 S.n981 0.074
R2188 S.n320 S.n319 0.074
R2189 S.n3934 S.n3933 0.071
R2190 S.n3460 S.n3459 0.071
R2191 S.n2974 S.n2973 0.071
R2192 S.n2465 S.n2464 0.071
R2193 S.n1944 S.n1943 0.071
R2194 S.n1399 S.n1398 0.071
R2195 S.n872 S.n871 0.071
R2196 S.n900 S.n899 0.071
R2197 S.n5067 S.n5066 0.07
R2198 S.n133 S.n131 0.067
R2199 S.n133 S.n132 0.067
R2200 S.n95 S.n93 0.067
R2201 S.n95 S.n94 0.067
R2202 S.n114 S.n112 0.067
R2203 S.n114 S.n113 0.067
R2204 S.n123 S.n121 0.067
R2205 S.n123 S.n122 0.067
R2206 S.n6 S.n4 0.067
R2207 S.n6 S.n5 0.067
R2208 S.n82 S.n80 0.067
R2209 S.n82 S.n81 0.067
R2210 S.n14 S.n12 0.067
R2211 S.n14 S.n13 0.067
R2212 S.n70 S.n68 0.067
R2213 S.n70 S.n69 0.067
R2214 S.n23 S.n21 0.067
R2215 S.n23 S.n22 0.067
R2216 S.n57 S.n55 0.067
R2217 S.n57 S.n56 0.067
R2218 S.n27 S.n26 0.067
R2219 S.n27 S.n25 0.067
R2220 S.n665 S.n655 0.067
R2221 S.n665 S.n653 0.067
R2222 S.n1787 S.n1778 0.067
R2223 S.n1787 S.n1777 0.067
R2224 S.n2337 S.n2328 0.067
R2225 S.n2337 S.n2327 0.067
R2226 S.n2878 S.n2869 0.067
R2227 S.n2878 S.n2868 0.067
R2228 S.n3393 S.n3384 0.067
R2229 S.n3393 S.n3383 0.067
R2230 S.n3899 S.n3890 0.067
R2231 S.n3899 S.n3889 0.067
R2232 S.n50 S.n49 0.066
R2233 S.n558 S.n557 0.066
R2234 S.n667 S.n666 0.065
R2235 S.n933 S.n932 0.063
R2236 S.n1156 S.n1155 0.063
R2237 S.n1470 S.n1469 0.063
R2238 S.n1679 S.n1678 0.063
R2239 S.n2014 S.n2013 0.063
R2240 S.n2275 S.n2274 0.063
R2241 S.n2535 S.n2534 0.063
R2242 S.n2800 S.n2799 0.063
R2243 S.n3044 S.n3043 0.063
R2244 S.n3299 S.n3298 0.063
R2245 S.n3530 S.n3529 0.063
R2246 S.n3667 S.n3666 0.063
R2247 S.n4004 S.n4003 0.063
R2248 S.n4253 S.n4252 0.063
R2249 S.n4448 S.n4447 0.063
R2250 S.n4684 S.n4683 0.063
R2251 S.n4857 S.n4856 0.063
R2252 S.n5047 S.n5046 0.063
R2253 S.n608 S.n595 0.063
R2254 S.n846 S.n820 0.063
R2255 S.n1096 S.n1082 0.063
R2256 S.n1383 S.n1382 0.063
R2257 S.n1619 S.n1618 0.063
R2258 S.n1928 S.n1927 0.063
R2259 S.n2215 S.n2214 0.063
R2260 S.n2449 S.n2448 0.063
R2261 S.n2740 S.n2739 0.063
R2262 S.n2958 S.n2957 0.063
R2263 S.n3239 S.n3238 0.063
R2264 S.n3444 S.n3443 0.063
R2265 S.n3607 S.n3606 0.063
R2266 S.n908 S.n888 0.063
R2267 S.n1438 S.n1425 0.063
R2268 S.n1982 S.n1970 0.063
R2269 S.n2503 S.n2491 0.063
R2270 S.n3012 S.n3000 0.063
R2271 S.n3498 S.n3486 0.063
R2272 S.n3972 S.n3960 0.063
R2273 S.n4416 S.n4404 0.063
R2274 S.n587 S.n567 0.063
R2275 S.n2926 S.n2905 0.063
R2276 S.n2417 S.n2396 0.063
R2277 S.n1896 S.n1875 0.063
R2278 S.n1350 S.n1329 0.063
R2279 S.n812 S.n793 0.063
R2280 S.n294 S.n279 0.063
R2281 S.n784 S.n783 0.063
R2282 S.n1055 S.n1054 0.063
R2283 S.n1321 S.n1320 0.063
R2284 S.n1583 S.n1582 0.063
R2285 S.n1867 S.n1866 0.063
R2286 S.n2182 S.n2181 0.063
R2287 S.n2388 S.n2387 0.063
R2288 S.n2704 S.n2703 0.063
R2289 S.n1835 S.n1814 0.063
R2290 S.n1289 S.n1268 0.063
R2291 S.n754 S.n734 0.063
R2292 S.n250 S.n235 0.063
R2293 S.n725 S.n724 0.063
R2294 S.n1019 S.n1018 0.063
R2295 S.n1260 S.n1259 0.063
R2296 S.n1547 S.n1546 0.063
R2297 S.n695 S.n675 0.063
R2298 S.n206 S.n191 0.063
R2299 S.n638 S.n637 0.063
R2300 S.n134 S.n133 0.062
R2301 S.n83 S.n82 0.062
R2302 S.n71 S.n70 0.062
R2303 S.n58 S.n57 0.062
R2304 S.n124 S.n123 0.062
R2305 S.n115 S.n114 0.061
R2306 S.n7 S.n6 0.06
R2307 S.n15 S.n14 0.06
R2308 S.n24 S.n23 0.06
R2309 S.n28 S.n27 0.06
R2310 S S.n5509 0.06
R2311 S.n4865 S.n4864 0.059
R2312 S.n1368 S.n1358 0.059
R2313 S.n96 S.n95 0.059
R2314 S.n1790 S.n1789 0.058
R2315 S.n2340 S.n2339 0.058
R2316 S.n2881 S.n2880 0.058
R2317 S.n3396 S.n3395 0.058
R2318 S.n3902 S.n3901 0.058
R2319 S.n4380 S.n4379 0.058
R2320 S.n667 S.n665 0.058
R2321 S.n5307 S.n5306 0.055
R2322 S.n53 S.n34 0.055
R2323 S.n322 S.n305 0.054
R2324 S.n3205 S.n3188 0.054
R2325 S.n3590 S.n3572 0.054
R2326 S.n4195 S.n4181 0.054
R2327 S.n4647 S.n4638 0.054
R2328 S.n5030 S.n5023 0.054
R2329 S.n2145 S.n2128 0.054
R2330 S.n2687 S.n2669 0.054
R2331 S.n985 S.n968 0.054
R2332 S.n1530 S.n1512 0.054
R2333 S.n5241 S.n5240 0.054
R2334 S.n649 S.n648 0.054
R2335 S.n1213 S.n1212 0.054
R2336 S.n1774 S.n1773 0.054
R2337 S.n2324 S.n2323 0.054
R2338 S.n2865 S.n2864 0.054
R2339 S.n3380 S.n3379 0.054
R2340 S.n3886 S.n3885 0.054
R2341 S.n4366 S.n4365 0.054
R2342 S.n4815 S.n4814 0.054
R2343 S.n5494 S.n5493 0.054
R2344 S.n318 S.n317 0.053
R2345 S.n980 S.n979 0.053
R2346 S.n1526 S.n1525 0.053
R2347 S.n2140 S.n2139 0.053
R2348 S.n2683 S.n2682 0.053
R2349 S.n3200 S.n3199 0.053
R2350 S.n3586 S.n3585 0.053
R2351 S.n4190 S.n4189 0.053
R2352 S.n5326 S.n5325 0.053
R2353 S.n5074 S.n5073 0.053
R2354 S.n644 S.n643 0.053
R2355 S.n611 S.n610 0.053
R2356 S.n936 S.n935 0.053
R2357 S.n5348 S.n5347 0.053
R2358 S.n5050 S.n5049 0.053
R2359 S.n4860 S.n4859 0.053
R2360 S.n4687 S.n4686 0.053
R2361 S.n4451 S.n4450 0.053
R2362 S.n4256 S.n4255 0.053
R2363 S.n4007 S.n4006 0.053
R2364 S.n3670 S.n3669 0.053
R2365 S.n3533 S.n3532 0.053
R2366 S.n3302 S.n3301 0.053
R2367 S.n3047 S.n3046 0.053
R2368 S.n2803 S.n2802 0.053
R2369 S.n2538 S.n2537 0.053
R2370 S.n2278 S.n2277 0.053
R2371 S.n2017 S.n2016 0.053
R2372 S.n1682 S.n1681 0.053
R2373 S.n1473 S.n1472 0.053
R2374 S.n1159 S.n1158 0.053
R2375 S.n478 S.n477 0.053
R2376 S.n274 S.n273 0.053
R2377 S.n787 S.n786 0.053
R2378 S.n3076 S.n3075 0.053
R2379 S.n2707 S.n2706 0.053
R2380 S.n2391 S.n2390 0.053
R2381 S.n2169 S.n2168 0.053
R2382 S.n1870 S.n1869 0.053
R2383 S.n1586 S.n1585 0.053
R2384 S.n1324 S.n1323 0.053
R2385 S.n1058 S.n1057 0.053
R2386 S.n297 S.n296 0.053
R2387 S.n3567 S.n3566 0.053
R2388 S.n3223 S.n3222 0.053
R2389 S.n2929 S.n2928 0.053
R2390 S.n2724 S.n2723 0.053
R2391 S.n2420 S.n2419 0.053
R2392 S.n2199 S.n2198 0.053
R2393 S.n1899 S.n1898 0.053
R2394 S.n1603 S.n1602 0.053
R2395 S.n1353 S.n1352 0.053
R2396 S.n1077 S.n1076 0.053
R2397 S.n1099 S.n1098 0.053
R2398 S.n849 S.n848 0.053
R2399 S.n505 S.n504 0.053
R2400 S.n528 S.n527 0.053
R2401 S.n1386 S.n1385 0.053
R2402 S.n1931 S.n1930 0.053
R2403 S.n2452 S.n2451 0.053
R2404 S.n2961 S.n2960 0.053
R2405 S.n3447 S.n3446 0.053
R2406 S.n4039 S.n4038 0.053
R2407 S.n3610 S.n3609 0.053
R2408 S.n3242 S.n3241 0.053
R2409 S.n2743 S.n2742 0.053
R2410 S.n2218 S.n2217 0.053
R2411 S.n1622 S.n1621 0.053
R2412 S.n883 S.n882 0.053
R2413 S.n442 S.n441 0.053
R2414 S.n561 S.n560 0.053
R2415 S.n4481 S.n4480 0.053
R2416 S.n4217 S.n4216 0.053
R2417 S.n3955 S.n3954 0.053
R2418 S.n3631 S.n3630 0.053
R2419 S.n3481 S.n3480 0.053
R2420 S.n3263 S.n3262 0.053
R2421 S.n2995 S.n2994 0.053
R2422 S.n2764 S.n2763 0.053
R2423 S.n2486 S.n2485 0.053
R2424 S.n2239 S.n2238 0.053
R2425 S.n1965 S.n1964 0.053
R2426 S.n1643 S.n1642 0.053
R2427 S.n1420 S.n1419 0.053
R2428 S.n1120 S.n1119 0.053
R2429 S.n911 S.n910 0.053
R2430 S.n461 S.n460 0.053
R2431 S.n1140 S.n1139 0.053
R2432 S.n1441 S.n1440 0.053
R2433 S.n1663 S.n1662 0.053
R2434 S.n1985 S.n1984 0.053
R2435 S.n2259 S.n2258 0.053
R2436 S.n2506 S.n2505 0.053
R2437 S.n2784 S.n2783 0.053
R2438 S.n3015 S.n3014 0.053
R2439 S.n3283 S.n3282 0.053
R2440 S.n3501 S.n3500 0.053
R2441 S.n3651 S.n3650 0.053
R2442 S.n3975 S.n3974 0.053
R2443 S.n4237 S.n4236 0.053
R2444 S.n4419 S.n4418 0.053
R2445 S.n4668 S.n4667 0.053
R2446 S.n4887 S.n4886 0.053
R2447 S.n590 S.n589 0.053
R2448 S.n815 S.n814 0.053
R2449 S.n422 S.n421 0.053
R2450 S.n405 S.n404 0.053
R2451 S.n230 S.n229 0.053
R2452 S.n728 S.n727 0.053
R2453 S.n2046 S.n2045 0.053
R2454 S.n1550 S.n1549 0.053
R2455 S.n1263 S.n1262 0.053
R2456 S.n1022 S.n1021 0.053
R2457 S.n253 S.n252 0.053
R2458 S.n2572 S.n2571 0.053
R2459 S.n2163 S.n2162 0.053
R2460 S.n1838 S.n1837 0.053
R2461 S.n1567 S.n1566 0.053
R2462 S.n1292 S.n1291 0.053
R2463 S.n1039 S.n1038 0.053
R2464 S.n757 S.n756 0.053
R2465 S.n389 S.n388 0.053
R2466 S.n372 S.n371 0.053
R2467 S.n189 S.n188 0.053
R2468 S.n963 S.n962 0.053
R2469 S.n209 S.n208 0.053
R2470 S.n1507 S.n1506 0.053
R2471 S.n1003 S.n1002 0.053
R2472 S.n698 S.n697 0.053
R2473 S.n356 S.n355 0.053
R2474 S.n339 S.n338 0.053
R2475 S.n499 S.n498 0.053
R2476 S.n1208 S.n1207 0.053
R2477 S.n1185 S.n1184 0.053
R2478 S.n1754 S.n1753 0.053
R2479 S.n1727 S.n1726 0.053
R2480 S.n2083 S.n2082 0.053
R2481 S.n2056 S.n2055 0.053
R2482 S.n2609 S.n2608 0.053
R2483 S.n2582 S.n2581 0.053
R2484 S.n3113 S.n3112 0.053
R2485 S.n3086 S.n3085 0.053
R2486 S.n3790 S.n3789 0.053
R2487 S.n3763 S.n3762 0.053
R2488 S.n4076 S.n4075 0.053
R2489 S.n4049 S.n4048 0.053
R2490 S.n4518 S.n4517 0.053
R2491 S.n4491 S.n4490 0.053
R2492 S.n4907 S.n4906 0.053
R2493 S.n5094 S.n5093 0.053
R2494 S.n5366 S.n5365 0.053
R2495 S.n1179 S.n1178 0.053
R2496 S.n1769 S.n1768 0.053
R2497 S.n5381 S.n5380 0.053
R2498 S.n5109 S.n5108 0.053
R2499 S.n4923 S.n4922 0.053
R2500 S.n4534 S.n4533 0.053
R2501 S.n4549 S.n4548 0.053
R2502 S.n4092 S.n4091 0.053
R2503 S.n4107 S.n4106 0.053
R2504 S.n3806 S.n3805 0.053
R2505 S.n3821 S.n3820 0.053
R2506 S.n3129 S.n3128 0.053
R2507 S.n3144 S.n3143 0.053
R2508 S.n2625 S.n2624 0.053
R2509 S.n2640 S.n2639 0.053
R2510 S.n2099 S.n2098 0.053
R2511 S.n2114 S.n2113 0.053
R2512 S.n1701 S.n1700 0.053
R2513 S.n1721 S.n1720 0.053
R2514 S.n2319 S.n2318 0.053
R2515 S.n5396 S.n5395 0.053
R2516 S.n5125 S.n5124 0.053
R2517 S.n4938 S.n4937 0.053
R2518 S.n4706 S.n4705 0.053
R2519 S.n4564 S.n4563 0.053
R2520 S.n4276 S.n4275 0.053
R2521 S.n4122 S.n4121 0.053
R2522 S.n3690 S.n3689 0.053
R2523 S.n3836 S.n3835 0.053
R2524 S.n3322 S.n3321 0.053
R2525 S.n3159 S.n3158 0.053
R2526 S.n2823 S.n2822 0.053
R2527 S.n2655 S.n2654 0.053
R2528 S.n2305 S.n2304 0.053
R2529 S.n2302 S.n2301 0.053
R2530 S.n2860 S.n2859 0.053
R2531 S.n5411 S.n5410 0.053
R2532 S.n5141 S.n5140 0.053
R2533 S.n4953 S.n4952 0.053
R2534 S.n4722 S.n4721 0.053
R2535 S.n4579 S.n4578 0.053
R2536 S.n4292 S.n4291 0.053
R2537 S.n4137 S.n4136 0.053
R2538 S.n3706 S.n3705 0.053
R2539 S.n3851 S.n3850 0.053
R2540 S.n3338 S.n3337 0.053
R2541 S.n3174 S.n3173 0.053
R2542 S.n2846 S.n2845 0.053
R2543 S.n2843 S.n2842 0.053
R2544 S.n3375 S.n3374 0.053
R2545 S.n5426 S.n5425 0.053
R2546 S.n5157 S.n5156 0.053
R2547 S.n4968 S.n4967 0.053
R2548 S.n4738 S.n4737 0.053
R2549 S.n4594 S.n4593 0.053
R2550 S.n4308 S.n4307 0.053
R2551 S.n4152 S.n4151 0.053
R2552 S.n3722 S.n3721 0.053
R2553 S.n3866 S.n3865 0.053
R2554 S.n3361 S.n3360 0.053
R2555 S.n3346 S.n3345 0.053
R2556 S.n3881 S.n3880 0.053
R2557 S.n5441 S.n5440 0.053
R2558 S.n5173 S.n5172 0.053
R2559 S.n4983 S.n4982 0.053
R2560 S.n4754 S.n4753 0.053
R2561 S.n4609 S.n4608 0.053
R2562 S.n4324 S.n4323 0.053
R2563 S.n4167 S.n4166 0.053
R2564 S.n3737 S.n3736 0.053
R2565 S.n3757 S.n3756 0.053
R2566 S.n4361 S.n4360 0.053
R2567 S.n5456 S.n5455 0.053
R2568 S.n5189 S.n5188 0.053
R2569 S.n4998 S.n4997 0.053
R2570 S.n4770 S.n4769 0.053
R2571 S.n4624 S.n4623 0.053
R2572 S.n4347 S.n4346 0.053
R2573 S.n4344 S.n4343 0.053
R2574 S.n4810 S.n4809 0.053
R2575 S.n5471 S.n5470 0.053
R2576 S.n5205 S.n5204 0.053
R2577 S.n5013 S.n5012 0.053
R2578 S.n4796 S.n4795 0.053
R2579 S.n4793 S.n4792 0.053
R2580 S.n5236 S.n5235 0.053
R2581 S.n5489 S.n5488 0.053
R2582 S.n5211 S.n5210 0.053
R2583 S.n672 S.n671 0.052
R2584 S.n1800 S.n1799 0.052
R2585 S.n1234 S.n1233 0.052
R2586 S.n2350 S.n2349 0.052
R2587 S.n1812 S.n1811 0.052
R2588 S.n2891 S.n2890 0.052
R2589 S.n2362 S.n2361 0.052
R2590 S.n3406 S.n3405 0.052
R2591 S.n2903 S.n2902 0.052
R2592 S.n3912 S.n3911 0.052
R2593 S.n3418 S.n3417 0.052
R2594 S.n4390 S.n4389 0.052
R2595 S.n3924 S.n3923 0.052
R2596 S.n4402 S.n4401 0.052
R2597 S.n5258 S.n5257 0.052
R2598 S.n5066 S.n5065 0.052
R2599 S.n512 S.n511 0.051
R2600 S.n4031 S.n4029 0.051
R2601 S.n3540 S.n3539 0.051
R2602 S.n3068 S.n3066 0.051
R2603 S.n2545 S.n2544 0.051
R2604 S.n2038 S.n2036 0.051
R2605 S.n1480 S.n1479 0.051
R2606 S.n955 S.n953 0.051
R2607 S.n617 S.n616 0.051
R2608 S.n653 S.n652 0.051
R2609 S.n655 S.n654 0.051
R2610 S.n4033 S.n4032 0.05
R2611 S.n4881 S.n4868 0.05
R2612 S.n581 S.n578 0.05
R2613 S.n3558 S.n3555 0.05
R2614 S.n3561 S.n3542 0.05
R2615 S.n3070 S.n3069 0.05
R2616 S.n2561 S.n2560 0.05
R2617 S.n2566 S.n2547 0.05
R2618 S.n2040 S.n2039 0.05
R2619 S.n1496 S.n1495 0.05
R2620 S.n1501 S.n1482 0.05
R2621 S.n957 S.n956 0.05
R2622 S.n638 S.n619 0.05
R2623 S.n598 S.n597 0.05
R2624 S.n1109 S.n1108 0.049
R2625 S.n1632 S.n1631 0.049
R2626 S.n2228 S.n2227 0.049
R2627 S.n2753 S.n2752 0.049
R2628 S.n3252 S.n3251 0.049
R2629 S.n3620 S.n3619 0.049
R2630 S.n4206 S.n4205 0.049
R2631 S.n436 S.n435 0.049
R2632 S.n455 S.n454 0.049
R2633 S.n4829 S.n4827 0.049
R2634 S.n4786 S.n4785 0.048
R2635 S S.n164 0.048
R2636 S.n1225 S.n1224 0.048
R2637 S.n1788 S.n1787 0.048
R2638 S.n2338 S.n2337 0.048
R2639 S.n2879 S.n2878 0.048
R2640 S.n3394 S.n3393 0.048
R2641 S.n3900 S.n3899 0.048
R2642 S.n4378 S.n4377 0.048
R2643 S.n4826 S.n4825 0.048
R2644 S.n5323 S.n5321 0.047
R2645 S.n5071 S.n5062 0.047
R2646 S.n5260 S.n5243 0.047
R2647 S.n638 S.n629 0.047
R2648 S.n608 S.n606 0.047
R2649 S.n933 S.n919 0.047
R2650 S.n5342 S.n5334 0.047
R2651 S.n5047 S.n5039 0.047
R2652 S.n4857 S.n4845 0.047
R2653 S.n4684 S.n4676 0.047
R2654 S.n4448 S.n4436 0.047
R2655 S.n4253 S.n4245 0.047
R2656 S.n4004 S.n3992 0.047
R2657 S.n3667 S.n3659 0.047
R2658 S.n3530 S.n3518 0.047
R2659 S.n3299 S.n3291 0.047
R2660 S.n3044 S.n3032 0.047
R2661 S.n2800 S.n2792 0.047
R2662 S.n2535 S.n2523 0.047
R2663 S.n2275 S.n2267 0.047
R2664 S.n2014 S.n2002 0.047
R2665 S.n1679 S.n1671 0.047
R2666 S.n1470 S.n1458 0.047
R2667 S.n1156 S.n1148 0.047
R2668 S.n475 S.n473 0.047
R2669 S.n271 S.n269 0.047
R2670 S.n784 S.n774 0.047
R2671 S.n3070 S.n3056 0.047
R2672 S.n2704 S.n2696 0.047
R2673 S.n2388 S.n2376 0.047
R2674 S.n2182 S.n2174 0.047
R2675 S.n1867 S.n1855 0.047
R2676 S.n1583 S.n1575 0.047
R2677 S.n1321 S.n1309 0.047
R2678 S.n1055 S.n1047 0.047
R2679 S.n294 S.n292 0.047
R2680 S.n3561 S.n3552 0.047
R2681 S.n3220 S.n3218 0.047
R2682 S.n2926 S.n2915 0.047
R2683 S.n2721 S.n2719 0.047
R2684 S.n2417 S.n2406 0.047
R2685 S.n2196 S.n2194 0.047
R2686 S.n1896 S.n1885 0.047
R2687 S.n1600 S.n1598 0.047
R2688 S.n1350 S.n1339 0.047
R2689 S.n1074 S.n1070 0.047
R2690 S.n1096 S.n1091 0.047
R2691 S.n846 S.n831 0.047
R2692 S.n510 S.n508 0.047
R2693 S.n525 S.n519 0.047
R2694 S.n1383 S.n1371 0.047
R2695 S.n1928 S.n1916 0.047
R2696 S.n2449 S.n2437 0.047
R2697 S.n2958 S.n2946 0.047
R2698 S.n3444 S.n3432 0.047
R2699 S.n4033 S.n4019 0.047
R2700 S.n3607 S.n3599 0.047
R2701 S.n3239 S.n3231 0.047
R2702 S.n2740 S.n2732 0.047
R2703 S.n2215 S.n2207 0.047
R2704 S.n1619 S.n1611 0.047
R2705 S.n880 S.n870 0.047
R2706 S.n439 S.n433 0.047
R2707 S.n558 S.n551 0.047
R2708 S.n4475 S.n4467 0.047
R2709 S.n4214 S.n4209 0.047
R2710 S.n3952 S.n3937 0.047
R2711 S.n3628 S.n3623 0.047
R2712 S.n3478 S.n3463 0.047
R2713 S.n3260 S.n3255 0.047
R2714 S.n2992 S.n2977 0.047
R2715 S.n2761 S.n2756 0.047
R2716 S.n2483 S.n2468 0.047
R2717 S.n2236 S.n2231 0.047
R2718 S.n1962 S.n1947 0.047
R2719 S.n1640 S.n1635 0.047
R2720 S.n1417 S.n1402 0.047
R2721 S.n1117 S.n1112 0.047
R2722 S.n908 S.n898 0.047
R2723 S.n458 S.n453 0.047
R2724 S.n1137 S.n1131 0.047
R2725 S.n1438 S.n1435 0.047
R2726 S.n1660 S.n1655 0.047
R2727 S.n1982 S.n1980 0.047
R2728 S.n2256 S.n2251 0.047
R2729 S.n2503 S.n2501 0.047
R2730 S.n2781 S.n2776 0.047
R2731 S.n3012 S.n3010 0.047
R2732 S.n3280 S.n3275 0.047
R2733 S.n3498 S.n3496 0.047
R2734 S.n3648 S.n3643 0.047
R2735 S.n3972 S.n3970 0.047
R2736 S.n4234 S.n4229 0.047
R2737 S.n4416 S.n4414 0.047
R2738 S.n4665 S.n4660 0.047
R2739 S.n4881 S.n4879 0.047
R2740 S.n587 S.n577 0.047
R2741 S.n812 S.n802 0.047
R2742 S.n419 S.n417 0.047
R2743 S.n402 S.n400 0.047
R2744 S.n227 S.n225 0.047
R2745 S.n725 S.n715 0.047
R2746 S.n2040 S.n2026 0.047
R2747 S.n1547 S.n1539 0.047
R2748 S.n1260 S.n1248 0.047
R2749 S.n1019 S.n1011 0.047
R2750 S.n250 S.n248 0.047
R2751 S.n2566 S.n2557 0.047
R2752 S.n2160 S.n2158 0.047
R2753 S.n1835 S.n1824 0.047
R2754 S.n1564 S.n1562 0.047
R2755 S.n1289 S.n1278 0.047
R2756 S.n1036 S.n1034 0.047
R2757 S.n754 S.n743 0.047
R2758 S.n386 S.n384 0.047
R2759 S.n369 S.n367 0.047
R2760 S.n186 S.n184 0.047
R2761 S.n957 S.n945 0.047
R2762 S.n206 S.n204 0.047
R2763 S.n1501 S.n1492 0.047
R2764 S.n1000 S.n998 0.047
R2765 S.n695 S.n684 0.047
R2766 S.n353 S.n351 0.047
R2767 S.n336 S.n334 0.047
R2768 S.n668 S.n651 0.047
R2769 S.n493 S.n490 0.047
R2770 S.n1202 S.n1199 0.047
R2771 S.n1192 S.n1188 0.047
R2772 S.n1748 S.n1742 0.047
R2773 S.n1734 S.n1730 0.047
R2774 S.n2077 S.n2071 0.047
R2775 S.n2063 S.n2059 0.047
R2776 S.n2603 S.n2597 0.047
R2777 S.n2589 S.n2585 0.047
R2778 S.n3107 S.n3101 0.047
R2779 S.n3093 S.n3089 0.047
R2780 S.n3784 S.n3778 0.047
R2781 S.n3770 S.n3766 0.047
R2782 S.n4070 S.n4064 0.047
R2783 S.n4056 S.n4052 0.047
R2784 S.n4512 S.n4506 0.047
R2785 S.n4498 S.n4494 0.047
R2786 S.n4901 S.n4895 0.047
R2787 S.n5088 S.n5084 0.047
R2788 S.n5360 S.n5355 0.047
R2789 S.n1229 S.n1215 0.047
R2790 S.n1173 S.n1171 0.047
R2791 S.n1763 S.n1759 0.047
R2792 S.n5375 S.n5371 0.047
R2793 S.n5103 S.n5099 0.047
R2794 S.n4917 S.n4912 0.047
R2795 S.n4541 S.n4531 0.047
R2796 S.n4543 S.n4523 0.047
R2797 S.n4099 S.n4089 0.047
R2798 S.n4101 S.n4081 0.047
R2799 S.n3813 S.n3803 0.047
R2800 S.n3815 S.n3795 0.047
R2801 S.n3136 S.n3126 0.047
R2802 S.n3138 S.n3118 0.047
R2803 S.n2632 S.n2622 0.047
R2804 S.n2634 S.n2614 0.047
R2805 S.n2106 S.n2096 0.047
R2806 S.n2108 S.n2088 0.047
R2807 S.n1695 S.n1691 0.047
R2808 S.n1808 S.n1776 0.047
R2809 S.n1715 S.n1709 0.047
R2810 S.n2313 S.n2119 0.047
R2811 S.n5390 S.n5386 0.047
R2812 S.n5119 S.n5114 0.047
R2813 S.n4932 S.n4928 0.047
R2814 S.n4700 S.n4695 0.047
R2815 S.n4558 S.n4554 0.047
R2816 S.n4270 S.n4265 0.047
R2817 S.n4116 S.n4112 0.047
R2818 S.n3684 S.n3679 0.047
R2819 S.n3830 S.n3826 0.047
R2820 S.n3316 S.n3311 0.047
R2821 S.n3153 S.n3149 0.047
R2822 S.n2817 S.n2812 0.047
R2823 S.n2649 S.n2645 0.047
R2824 S.n2312 S.n2127 0.047
R2825 S.n2358 S.n2326 0.047
R2826 S.n2296 S.n2290 0.047
R2827 S.n2854 S.n2660 0.047
R2828 S.n5405 S.n5401 0.047
R2829 S.n5135 S.n5130 0.047
R2830 S.n4947 S.n4943 0.047
R2831 S.n4716 S.n4711 0.047
R2832 S.n4573 S.n4569 0.047
R2833 S.n4286 S.n4281 0.047
R2834 S.n4131 S.n4127 0.047
R2835 S.n3700 S.n3695 0.047
R2836 S.n3845 S.n3841 0.047
R2837 S.n3332 S.n3327 0.047
R2838 S.n3168 S.n3164 0.047
R2839 S.n2853 S.n2668 0.047
R2840 S.n2899 S.n2867 0.047
R2841 S.n2837 S.n2831 0.047
R2842 S.n3369 S.n3179 0.047
R2843 S.n5420 S.n5416 0.047
R2844 S.n5151 S.n5146 0.047
R2845 S.n4962 S.n4958 0.047
R2846 S.n4732 S.n4727 0.047
R2847 S.n4588 S.n4584 0.047
R2848 S.n4302 S.n4297 0.047
R2849 S.n4146 S.n4142 0.047
R2850 S.n3716 S.n3711 0.047
R2851 S.n3860 S.n3856 0.047
R2852 S.n3368 S.n3187 0.047
R2853 S.n3414 S.n3382 0.047
R2854 S.n3355 S.n3349 0.047
R2855 S.n3875 S.n3871 0.047
R2856 S.n5435 S.n5431 0.047
R2857 S.n5167 S.n5162 0.047
R2858 S.n4977 S.n4973 0.047
R2859 S.n4748 S.n4743 0.047
R2860 S.n4603 S.n4599 0.047
R2861 S.n4318 S.n4313 0.047
R2862 S.n4161 S.n4157 0.047
R2863 S.n3731 S.n3727 0.047
R2864 S.n3920 S.n3888 0.047
R2865 S.n3751 S.n3745 0.047
R2866 S.n4355 S.n4172 0.047
R2867 S.n5450 S.n5446 0.047
R2868 S.n5183 S.n5178 0.047
R2869 S.n4992 S.n4988 0.047
R2870 S.n4764 S.n4759 0.047
R2871 S.n4618 S.n4614 0.047
R2872 S.n4354 S.n4180 0.047
R2873 S.n4398 S.n4368 0.047
R2874 S.n4338 S.n4332 0.047
R2875 S.n4804 S.n4629 0.047
R2876 S.n5465 S.n5461 0.047
R2877 S.n5199 S.n5194 0.047
R2878 S.n5007 S.n5003 0.047
R2879 S.n4803 S.n4637 0.047
R2880 S.n4831 S.n4817 0.047
R2881 S.n4787 S.n4776 0.047
R2882 S.n5230 S.n5227 0.047
R2883 S.n5483 S.n5481 0.047
R2884 S.n5216 S.n5214 0.047
R2885 S.n5498 S.n5496 0.047
R2886 S.n844 S.n839 0.047
R2887 S.n3428 S.n3427 0.047
R2888 S.n2942 S.n2941 0.047
R2889 S.n2433 S.n2432 0.047
R2890 S.n1912 S.n1911 0.047
R2891 S.n1367 S.n1366 0.047
R2892 S.t2 S.n97 0.046
R2893 S.t2 S.n87 0.046
R2894 S.t2 S.n75 0.046
R2895 S.t2 S.n63 0.046
R2896 S.n1202 S.n1192 0.046
R2897 S.n2313 S.n2312 0.045
R2898 S.n2854 S.n2853 0.045
R2899 S.n3369 S.n3368 0.045
R2900 S.n4355 S.n4354 0.045
R2901 S.n4804 S.n4803 0.045
R2902 S.n104 S.n102 0.045
R2903 S.n5229 S.n5228 0.045
R2904 S.n543 S.n542 0.045
R2905 S.n861 S.n853 0.045
R2906 S.n1414 S.n1406 0.045
R2907 S.n1959 S.n1951 0.045
R2908 S.n2480 S.n2472 0.045
R2909 S.n2989 S.n2981 0.045
R2910 S.n3475 S.n3467 0.045
R2911 S.n3949 S.n3941 0.045
R2912 S.n1792 S.n1791 0.045
R2913 S.n2342 S.n2341 0.045
R2914 S.n2883 S.n2882 0.045
R2915 S.n3398 S.n3397 0.045
R2916 S.n3904 S.n3903 0.045
R2917 S.n4382 S.n4381 0.045
R2918 S.n5230 S.n5216 0.044
R2919 S.n1748 S.n1735 0.044
R2920 S.n2077 S.n2064 0.044
R2921 S.n2603 S.n2590 0.044
R2922 S.n3107 S.n3094 0.044
R2923 S.n3784 S.n3771 0.044
R2924 S.n4070 S.n4057 0.044
R2925 S.n4512 S.n4499 0.044
R2926 S.n4901 S.n4888 0.044
R2927 S.n2108 S.n2107 0.044
R2928 S.n2634 S.n2633 0.044
R2929 S.n3138 S.n3137 0.044
R2930 S.n3815 S.n3814 0.044
R2931 S.n4101 S.n4100 0.044
R2932 S.n4543 S.n4542 0.044
R2933 S.n4917 S.n4916 0.044
R2934 S.n284 S.n283 0.044
R2935 S.n240 S.n239 0.044
R2936 S.n196 S.n195 0.044
R2937 S.n522 S.n521 0.043
R2938 S.n4868 S.n4867 0.043
R2939 S.n823 S.n822 0.043
R2940 S.n795 S.n794 0.042
R2941 S.n1331 S.n1330 0.042
R2942 S.n1877 S.n1876 0.042
R2943 S.n2398 S.n2397 0.042
R2944 S.n2907 S.n2906 0.042
R2945 S.n736 S.n735 0.042
R2946 S.n1270 S.n1269 0.042
R2947 S.n1816 S.n1815 0.042
R2948 S.n677 S.n676 0.042
R2949 S.n4853 S.n4850 0.042
R2950 S.n4444 S.n4441 0.042
R2951 S.n4000 S.n3997 0.042
R2952 S.n3526 S.n3523 0.042
R2953 S.n3040 S.n3037 0.042
R2954 S.n2531 S.n2528 0.042
R2955 S.n2010 S.n2007 0.042
R2956 S.n1466 S.n1463 0.042
R2957 S.n929 S.n924 0.042
R2958 S.n2384 S.n2381 0.042
R2959 S.n1863 S.n1860 0.042
R2960 S.n1317 S.n1314 0.042
R2961 S.n3440 S.n3437 0.042
R2962 S.n2954 S.n2951 0.042
R2963 S.n2445 S.n2442 0.042
R2964 S.n1924 S.n1921 0.042
R2965 S.n1379 S.n1376 0.042
R2966 S.n1256 S.n1253 0.042
R2967 S.n4406 S.n4405 0.042
R2968 S.n3962 S.n3961 0.042
R2969 S.n3488 S.n3487 0.042
R2970 S.n3002 S.n3001 0.042
R2971 S.n2493 S.n2492 0.042
R2972 S.n1972 S.n1971 0.042
R2973 S.n1427 S.n1426 0.042
R2974 S.n890 S.n889 0.042
R2975 S.n570 S.n569 0.041
R2976 S.n4016 S.n4015 0.041
R2977 S.n168 S.n167 0.041
R2978 S.n634 S.n632 0.04
R2979 S.n318 S.n309 0.04
R2980 S.n980 S.n971 0.04
R2981 S.n1526 S.n1517 0.04
R2982 S.n2140 S.n2131 0.04
R2983 S.n2683 S.n2674 0.04
R2984 S.n3200 S.n3191 0.04
R2985 S.n3586 S.n3577 0.04
R2986 S.n51 S.n40 0.04
R2987 S.n39 S.n38 0.039
R2988 S.n5249 S.n5248 0.039
R2989 S.n1793 S.n1792 0.039
R2990 S.n1798 S.n1797 0.039
R2991 S.n2343 S.n2342 0.039
R2992 S.n2348 S.n2347 0.039
R2993 S.n2884 S.n2883 0.039
R2994 S.n2889 S.n2888 0.039
R2995 S.n3399 S.n3398 0.039
R2996 S.n3404 S.n3403 0.039
R2997 S.n3905 S.n3904 0.039
R2998 S.n3910 S.n3909 0.039
R2999 S.n4383 S.n4382 0.039
R3000 S.n4388 S.n4387 0.039
R3001 S.n317 S.n310 0.039
R3002 S.n979 S.n972 0.039
R3003 S.n1525 S.n1518 0.039
R3004 S.n2139 S.n2132 0.039
R3005 S.n2682 S.n2675 0.039
R3006 S.n3199 S.n3192 0.039
R3007 S.n3585 S.n3578 0.039
R3008 S.n4189 S.n4183 0.039
R3009 S.n5026 S.n5024 0.038
R3010 S.n4841 S.n4840 0.038
R3011 S.n4432 S.n4431 0.038
R3012 S.n3988 S.n3987 0.038
R3013 S.n3514 S.n3513 0.038
R3014 S.n3028 S.n3027 0.038
R3015 S.n2519 S.n2518 0.038
R3016 S.n1998 S.n1997 0.038
R3017 S.n1454 S.n1453 0.038
R3018 S.n2372 S.n2371 0.038
R3019 S.n1851 S.n1850 0.038
R3020 S.n1305 S.n1304 0.038
R3021 S.n770 S.n769 0.038
R3022 S.n2924 S.n2919 0.038
R3023 S.n2415 S.n2410 0.038
R3024 S.n1894 S.n1889 0.038
R3025 S.n1348 S.n1343 0.038
R3026 S.n810 S.n806 0.038
R3027 S.n1244 S.n1243 0.038
R3028 S.n711 S.n710 0.038
R3029 S.n1833 S.n1828 0.038
R3030 S.n1287 S.n1282 0.038
R3031 S.n752 S.n747 0.038
R3032 S.n693 S.n688 0.038
R3033 S.n634 S.n633 0.038
R3034 S.n4474 S.n4472 0.037
R3035 S.n5249 S.n5246 0.037
R3036 S.n5248 S.n5247 0.037
R3037 S.n1417 S.n1399 0.037
R3038 S.n1962 S.n1944 0.037
R3039 S.n2483 S.n2465 0.037
R3040 S.n2992 S.n2974 0.037
R3041 S.n3478 S.n3460 0.037
R3042 S.n3952 S.n3934 0.037
R3043 S.n4475 S.n4464 0.037
R3044 S.n908 S.n900 0.037
R3045 S.n880 S.n872 0.037
R3046 S.n1798 S.n1795 0.037
R3047 S.n1797 S.n1796 0.037
R3048 S.n2348 S.n2345 0.037
R3049 S.n2347 S.n2346 0.037
R3050 S.n2889 S.n2886 0.037
R3051 S.n2888 S.n2887 0.037
R3052 S.n3404 S.n3401 0.037
R3053 S.n3403 S.n3402 0.037
R3054 S.n3910 S.n3907 0.037
R3055 S.n3909 S.n3908 0.037
R3056 S.n4388 S.n4385 0.037
R3057 S.n4387 S.n4386 0.037
R3058 S.n5474 S.n5473 0.037
R3059 S.n5220 S.n5219 0.037
R3060 S.n668 S.n168 0.036
R3061 S.n1136 S.n1135 0.036
R3062 S.n1648 S.n1647 0.036
R3063 S.n2244 S.n2243 0.036
R3064 S.n2769 S.n2768 0.036
R3065 S.n3268 S.n3267 0.036
R3066 S.n3636 S.n3635 0.036
R3067 S.n4222 S.n4221 0.036
R3068 S.n4653 S.n4652 0.036
R3069 S.n316 S.n311 0.036
R3070 S.n978 S.n973 0.036
R3071 S.n1524 S.n1519 0.036
R3072 S.n2138 S.n2133 0.036
R3073 S.n2681 S.n2676 0.036
R3074 S.n3198 S.n3193 0.036
R3075 S.n3584 S.n3579 0.036
R3076 S.n4188 S.n4184 0.036
R3077 S.n3211 S.n3210 0.035
R3078 S.n2712 S.n2711 0.035
R3079 S.n2187 S.n2186 0.035
R3080 S.n1591 S.n1590 0.035
R3081 S.n1063 S.n1062 0.035
R3082 S.n2151 S.n2150 0.035
R3083 S.n1555 S.n1554 0.035
R3084 S.n1027 S.n1026 0.035
R3085 S.n991 S.n990 0.035
R3086 S.n5314 S.n5313 0.035
R3087 S.n5250 S.n5249 0.035
R3088 S.n4841 S.n4836 0.035
R3089 S.n4432 S.n4427 0.035
R3090 S.n3988 S.n3983 0.035
R3091 S.n3514 S.n3509 0.035
R3092 S.n3028 S.n3023 0.035
R3093 S.n2519 S.n2514 0.035
R3094 S.n1998 S.n1993 0.035
R3095 S.n1454 S.n1449 0.035
R3096 S.n2372 S.n2367 0.035
R3097 S.n1851 S.n1846 0.035
R3098 S.n1305 S.n1300 0.035
R3099 S.n770 S.n765 0.035
R3100 S.n4033 S.n4016 0.035
R3101 S.n810 S.n809 0.035
R3102 S.n1348 S.n1347 0.035
R3103 S.n1894 S.n1893 0.035
R3104 S.n2415 S.n2414 0.035
R3105 S.n2924 S.n2923 0.035
R3106 S.n1244 S.n1239 0.035
R3107 S.n711 S.n706 0.035
R3108 S.n752 S.n751 0.035
R3109 S.n1287 S.n1286 0.035
R3110 S.n1833 S.n1832 0.035
R3111 S.n693 S.n692 0.035
R3112 S.n1791 S.n1790 0.035
R3113 S.n1801 S.n1798 0.035
R3114 S.n2341 S.n2340 0.035
R3115 S.n2351 S.n2348 0.035
R3116 S.n2882 S.n2881 0.035
R3117 S.n2892 S.n2889 0.035
R3118 S.n3397 S.n3396 0.035
R3119 S.n3407 S.n3404 0.035
R3120 S.n3903 S.n3902 0.035
R3121 S.n3913 S.n3910 0.035
R3122 S.n4381 S.n4380 0.035
R3123 S.n4391 S.n4388 0.035
R3124 S.n4821 S.n4820 0.034
R3125 S.n326 S.n325 0.034
R3126 S.n3209 S.n3208 0.034
R3127 S.n3594 S.n3593 0.034
R3128 S.n4199 S.n4198 0.034
R3129 S.n4651 S.n4650 0.034
R3130 S.n5034 S.n5033 0.034
R3131 S.n2149 S.n2148 0.034
R3132 S.n2691 S.n2690 0.034
R3133 S.n989 S.n988 0.034
R3134 S.n1534 S.n1533 0.034
R3135 S.n96 S.n92 0.034
R3136 S.n89 S.n88 0.034
R3137 S.n77 S.n76 0.034
R3138 S.n65 S.n64 0.034
R3139 S.n5360 S.n5356 0.034
R3140 S.n5088 S.n5085 0.034
R3141 S.n4901 S.n4897 0.034
R3142 S.n4498 S.n4495 0.034
R3143 S.n4512 S.n4508 0.034
R3144 S.n4056 S.n4053 0.034
R3145 S.n4070 S.n4066 0.034
R3146 S.n3770 S.n3767 0.034
R3147 S.n3784 S.n3780 0.034
R3148 S.n3093 S.n3090 0.034
R3149 S.n3107 S.n3103 0.034
R3150 S.n2589 S.n2586 0.034
R3151 S.n2603 S.n2599 0.034
R3152 S.n2063 S.n2060 0.034
R3153 S.n2077 S.n2073 0.034
R3154 S.n1734 S.n1731 0.034
R3155 S.n1748 S.n1744 0.034
R3156 S.n1192 S.n1189 0.034
R3157 S.n1229 S.n669 0.034
R3158 S.n1808 S.n1231 0.034
R3159 S.n2358 S.n1809 0.034
R3160 S.n2899 S.n2359 0.034
R3161 S.n3414 S.n2900 0.034
R3162 S.n3920 S.n3415 0.034
R3163 S.n4398 S.n3921 0.034
R3164 S.n4831 S.n4399 0.034
R3165 S.n5260 S.n5259 0.034
R3166 S.n4192 S.n4182 0.034
R3167 S.n3588 S.n3575 0.034
R3168 S.n3202 S.n3189 0.034
R3169 S.n2685 S.n2672 0.034
R3170 S.n2142 S.n2129 0.034
R3171 S.n1528 S.n1515 0.034
R3172 S.n982 S.n969 0.034
R3173 S.n320 S.n307 0.034
R3174 S.t0 S.n5301 0.034
R3175 S.t0 S.n5304 0.034
R3176 S.t2 S.n140 0.034
R3177 S.t2 S.n143 0.034
R3178 S.t2 S.n136 0.034
R3179 S.t2 S.n135 0.034
R3180 S.t2 S.n85 0.034
R3181 S.t2 S.n84 0.034
R3182 S.t2 S.n152 0.034
R3183 S.t2 S.n155 0.034
R3184 S.t2 S.n99 0.034
R3185 S.t2 S.n98 0.034
R3186 S.t2 S.n110 0.034
R3187 S.t2 S.n109 0.034
R3188 S.t2 S.n126 0.034
R3189 S.t2 S.n125 0.034
R3190 S.t2 S.n73 0.034
R3191 S.t2 S.n72 0.034
R3192 S.t2 S.n148 0.034
R3193 S.t2 S.n151 0.034
R3194 S.t2 S.n60 0.034
R3195 S.t2 S.n59 0.034
R3196 S.t2 S.n144 0.034
R3197 S.t2 S.n147 0.034
R3198 S.t0 S.n5265 0.034
R3199 S.t0 S.n5268 0.034
R3200 S.t0 S.n5269 0.034
R3201 S.t0 S.n5272 0.034
R3202 S.t0 S.n5273 0.034
R3203 S.t0 S.n5276 0.034
R3204 S.t0 S.n5277 0.034
R3205 S.t0 S.n5280 0.034
R3206 S.t0 S.n5281 0.034
R3207 S.t0 S.n5284 0.034
R3208 S.t0 S.n5285 0.034
R3209 S.t0 S.n5288 0.034
R3210 S.t0 S.n5289 0.034
R3211 S.t0 S.n5292 0.034
R3212 S.t0 S.n5293 0.034
R3213 S.t0 S.n5296 0.034
R3214 S.t0 S.n5297 0.034
R3215 S.t0 S.n5300 0.034
R3216 S.t0 S.n5262 0.034
R3217 S.t0 S.n5261 0.034
R3218 S.n51 S.n50 0.033
R3219 S.n1095 S.n1094 0.033
R3220 S.n5027 S.n5026 0.032
R3221 S.n4640 S.n4639 0.032
R3222 S.n950 S.n949 0.031
R3223 S.t12 S.n326 0.031
R3224 S.t95 S.n3209 0.031
R3225 S.t53 S.n3594 0.031
R3226 S.t66 S.n4199 0.031
R3227 S.t31 S.n4651 0.031
R3228 S.t44 S.n5034 0.031
R3229 S.t8 S.n2149 0.031
R3230 S.t168 S.n2691 0.031
R3231 S.t151 S.n989 0.031
R3232 S.t42 S.n1534 0.031
R3233 S.n4836 S.n4835 0.031
R3234 S.n4427 S.n4426 0.031
R3235 S.n3983 S.n3982 0.031
R3236 S.n3509 S.n3508 0.031
R3237 S.n3023 S.n3022 0.031
R3238 S.n2514 S.n2513 0.031
R3239 S.n1993 S.n1992 0.031
R3240 S.n1449 S.n1448 0.031
R3241 S.n2367 S.n2366 0.031
R3242 S.n1846 S.n1845 0.031
R3243 S.n1300 S.n1299 0.031
R3244 S.n765 S.n764 0.031
R3245 S.n809 S.n808 0.031
R3246 S.n1347 S.n1346 0.031
R3247 S.n1893 S.n1892 0.031
R3248 S.n2414 S.n2413 0.031
R3249 S.n2923 S.n2922 0.031
R3250 S.n1239 S.n1238 0.031
R3251 S.n706 S.n705 0.031
R3252 S.n751 S.n750 0.031
R3253 S.n1286 S.n1285 0.031
R3254 S.n1832 S.n1831 0.031
R3255 S.n692 S.n691 0.031
R3256 S.n158 S.n157 0.031
R3257 S.n159 S.n158 0.031
R3258 S.n160 S.n159 0.031
R3259 S.n161 S.n160 0.031
R3260 S.n162 S.n161 0.031
R3261 S.n163 S.n162 0.031
R3262 S.n164 S.n163 0.031
R3263 S.n166 S.n165 0.031
R3264 S.n5509 S.n5508 0.031
R3265 S.n5508 S.n5507 0.031
R3266 S.n5507 S.n5506 0.031
R3267 S.n5506 S.n5505 0.031
R3268 S.n5505 S.n5504 0.031
R3269 S.n5504 S.n5503 0.031
R3270 S.n5503 S.n5502 0.031
R3271 S.n5502 S.n5501 0.031
R3272 S.n5501 S.n5500 0.031
R3273 S.n5500 S.n5499 0.031
R3274 S.n5358 S.n5357 0.031
R3275 S.n4899 S.n4898 0.031
R3276 S.n4510 S.n4509 0.031
R3277 S.n4068 S.n4067 0.031
R3278 S.n3782 S.n3781 0.031
R3279 S.n3105 S.n3104 0.031
R3280 S.n2601 S.n2600 0.031
R3281 S.n2075 S.n2074 0.031
R3282 S.n1746 S.n1745 0.031
R3283 S.n2564 S.n2563 0.031
R3284 S.n1499 S.n1498 0.031
R3285 S.n3544 S.n3543 0.03
R3286 S.n2549 S.n2548 0.03
R3287 S.n1484 S.n1483 0.03
R3288 S.n3946 S.n3945 0.03
R3289 S.n3472 S.n3471 0.03
R3290 S.n2986 S.n2985 0.03
R3291 S.n2477 S.n2476 0.03
R3292 S.n1956 S.n1955 0.03
R3293 S.n1411 S.n1410 0.03
R3294 S.n858 S.n857 0.03
R3295 S.n536 S.n535 0.03
R3296 S.n621 S.n620 0.03
R3297 S.n3063 S.n3060 0.029
R3298 S.n4026 S.n4023 0.029
R3299 S.n2033 S.n2030 0.029
R3300 S.n929 S.n928 0.029
R3301 S.n1466 S.n1465 0.029
R3302 S.n2010 S.n2009 0.029
R3303 S.n2531 S.n2530 0.029
R3304 S.n3040 S.n3039 0.029
R3305 S.n3526 S.n3525 0.029
R3306 S.n4000 S.n3999 0.029
R3307 S.n4444 S.n4443 0.029
R3308 S.n4853 S.n4852 0.029
R3309 S.n1379 S.n1378 0.029
R3310 S.n1924 S.n1923 0.029
R3311 S.n2445 S.n2444 0.029
R3312 S.n2954 S.n2953 0.029
R3313 S.n3440 S.n3439 0.029
R3314 S.n1317 S.n1316 0.029
R3315 S.n1863 S.n1862 0.029
R3316 S.n2384 S.n2383 0.029
R3317 S.n1256 S.n1255 0.029
R3318 S.n1913 S.n1912 0.029
R3319 S.n2434 S.n2433 0.029
R3320 S.n2943 S.n2942 0.029
R3321 S.n3429 S.n3428 0.029
R3322 S.n3945 S.n3944 0.029
R3323 S.n3471 S.n3470 0.029
R3324 S.n2985 S.n2984 0.029
R3325 S.n2476 S.n2475 0.029
R3326 S.n1955 S.n1954 0.029
R3327 S.n1410 S.n1409 0.029
R3328 S.n857 S.n856 0.029
R3329 S.n535 S.n534 0.029
R3330 S.n4836 S.n4833 0.028
R3331 S.n4427 S.n4424 0.028
R3332 S.n3983 S.n3980 0.028
R3333 S.n3509 S.n3506 0.028
R3334 S.n3023 S.n3020 0.028
R3335 S.n2514 S.n2511 0.028
R3336 S.n1993 S.n1990 0.028
R3337 S.n1449 S.n1446 0.028
R3338 S.n2367 S.n2364 0.028
R3339 S.n1846 S.n1843 0.028
R3340 S.n1300 S.n1297 0.028
R3341 S.n765 S.n762 0.028
R3342 S.n1347 S.n1344 0.028
R3343 S.n1893 S.n1890 0.028
R3344 S.n2414 S.n2411 0.028
R3345 S.n2923 S.n2920 0.028
R3346 S.n1239 S.n1236 0.028
R3347 S.n706 S.n703 0.028
R3348 S.n751 S.n748 0.028
R3349 S.n1286 S.n1283 0.028
R3350 S.n1832 S.n1829 0.028
R3351 S.n692 S.n689 0.028
R3352 S.n1395 S.n1394 0.028
R3353 S.n1397 S.n1395 0.028
R3354 S.n1940 S.n1939 0.028
R3355 S.n1942 S.n1940 0.028
R3356 S.n2461 S.n2460 0.028
R3357 S.n2463 S.n2461 0.028
R3358 S.n2970 S.n2969 0.028
R3359 S.n2972 S.n2970 0.028
R3360 S.n3456 S.n3455 0.028
R3361 S.n3458 S.n3456 0.028
R3362 S.n3930 S.n3929 0.028
R3363 S.n3932 S.n3930 0.028
R3364 S.n4461 S.n4460 0.028
R3365 S.n4463 S.n4461 0.028
R3366 S.n874 S.n873 0.028
R3367 S.n876 S.n874 0.028
R3368 S.n902 S.n901 0.028
R3369 S.n904 S.n902 0.028
R3370 S.n662 S.n657 0.028
R3371 S.n1221 S.n1217 0.028
R3372 S.n1784 S.n1780 0.028
R3373 S.n2334 S.n2330 0.028
R3374 S.n2875 S.n2871 0.028
R3375 S.n3390 S.n3386 0.028
R3376 S.n3896 S.n3892 0.028
R3377 S.n4374 S.n4370 0.028
R3378 S.n5340 S.n5339 0.028
R3379 S.n4026 S.n4025 0.028
R3380 S.n3063 S.n3062 0.028
R3381 S.n2033 S.n2032 0.028
R3382 S.n1368 S.n1367 0.028
R3383 S.n5474 S.n5472 0.027
R3384 S.n5220 S.n5218 0.027
R3385 S.n558 S.n553 0.027
R3386 S.n580 S.n579 0.027
R3387 S.n3557 S.n3556 0.027
R3388 S.n2563 S.n2562 0.027
R3389 S.n1498 S.n1497 0.027
R3390 S.n1229 S.n1228 0.027
R3391 S.n1744 S.n1743 0.027
R3392 S.n2073 S.n2072 0.027
R3393 S.n2599 S.n2598 0.027
R3394 S.n3103 S.n3102 0.027
R3395 S.n3780 S.n3779 0.027
R3396 S.n4066 S.n4065 0.027
R3397 S.n4508 S.n4507 0.027
R3398 S.n4897 S.n4896 0.027
R3399 S.n1072 S.n1071 0.027
R3400 S.n933 S.n930 0.026
R3401 S.n1156 S.n1153 0.026
R3402 S.n1470 S.n1467 0.026
R3403 S.n1679 S.n1676 0.026
R3404 S.n2014 S.n2011 0.026
R3405 S.n2275 S.n2272 0.026
R3406 S.n2535 S.n2532 0.026
R3407 S.n2800 S.n2797 0.026
R3408 S.n3044 S.n3041 0.026
R3409 S.n3299 S.n3296 0.026
R3410 S.n3530 S.n3527 0.026
R3411 S.n3667 S.n3664 0.026
R3412 S.n4004 S.n4001 0.026
R3413 S.n4253 S.n4250 0.026
R3414 S.n4448 S.n4445 0.026
R3415 S.n4684 S.n4681 0.026
R3416 S.n4857 S.n4854 0.026
R3417 S.n5047 S.n5044 0.026
R3418 S.n5342 S.n5341 0.026
R3419 S.n475 S.n467 0.026
R3420 S.n846 S.n824 0.026
R3421 S.n1096 S.n1084 0.026
R3422 S.n1383 S.n1380 0.026
R3423 S.n1619 S.n1616 0.026
R3424 S.n1928 S.n1925 0.026
R3425 S.n2215 S.n2212 0.026
R3426 S.n2449 S.n2446 0.026
R3427 S.n2740 S.n2737 0.026
R3428 S.n2958 S.n2955 0.026
R3429 S.n3239 S.n3236 0.026
R3430 S.n3444 S.n3441 0.026
R3431 S.n3607 S.n3604 0.026
R3432 S.n4033 S.n4027 0.026
R3433 S.n1106 S.n1104 0.026
R3434 S.n1629 S.n1627 0.026
R3435 S.n2225 S.n2223 0.026
R3436 S.n2750 S.n2748 0.026
R3437 S.n3249 S.n3247 0.026
R3438 S.n3617 S.n3615 0.026
R3439 S.n4203 S.n4201 0.026
R3440 S.n4664 S.n4663 0.026
R3441 S.n4233 S.n4232 0.026
R3442 S.n3647 S.n3646 0.026
R3443 S.n3279 S.n3278 0.026
R3444 S.n2780 S.n2779 0.026
R3445 S.n2255 S.n2254 0.026
R3446 S.n1659 S.n1658 0.026
R3447 S.n1126 S.n1125 0.026
R3448 S.n908 S.n891 0.026
R3449 S.n1438 S.n1428 0.026
R3450 S.n1982 S.n1973 0.026
R3451 S.n2503 S.n2494 0.026
R3452 S.n3012 S.n3003 0.026
R3453 S.n3498 S.n3489 0.026
R3454 S.n3972 S.n3963 0.026
R3455 S.n4416 S.n4407 0.026
R3456 S.n4881 S.n4872 0.026
R3457 S.n587 S.n571 0.026
R3458 S.n3561 S.n3545 0.026
R3459 S.n2926 S.n2908 0.026
R3460 S.n2417 S.n2399 0.026
R3461 S.n1896 S.n1878 0.026
R3462 S.n1350 S.n1332 0.026
R3463 S.n812 S.n796 0.026
R3464 S.n784 S.n779 0.026
R3465 S.n1055 S.n1052 0.026
R3466 S.n1321 S.n1318 0.026
R3467 S.n1583 S.n1580 0.026
R3468 S.n1867 S.n1864 0.026
R3469 S.n2182 S.n2179 0.026
R3470 S.n2388 S.n2385 0.026
R3471 S.n2704 S.n2701 0.026
R3472 S.n3070 S.n3064 0.026
R3473 S.n2566 S.n2550 0.026
R3474 S.n1835 S.n1817 0.026
R3475 S.n1289 S.n1271 0.026
R3476 S.n754 S.n737 0.026
R3477 S.n725 S.n720 0.026
R3478 S.n1019 S.n1016 0.026
R3479 S.n1260 S.n1257 0.026
R3480 S.n1547 S.n1544 0.026
R3481 S.n2040 S.n2034 0.026
R3482 S.n1501 S.n1485 0.026
R3483 S.n695 S.n678 0.026
R3484 S.n957 S.n951 0.026
R3485 S.n638 S.n635 0.026
R3486 S.n638 S.n622 0.026
R3487 S.n5071 S.n5055 0.026
R3488 S.n525 S.n524 0.026
R3489 S.t2 S.n32 0.025
R3490 S.t2 S.n2 0.025
R3491 S.t2 S.n10 0.025
R3492 S.t2 S.n18 0.025
R3493 S.n118 S.n117 0.024
R3494 S.n1223 S.n1222 0.024
R3495 S.n1786 S.n1785 0.024
R3496 S.n2336 S.n2335 0.024
R3497 S.n2877 S.n2876 0.024
R3498 S.n3392 S.n3391 0.024
R3499 S.n3898 S.n3897 0.024
R3500 S.n4376 S.n4375 0.024
R3501 S.n4824 S.n4823 0.024
R3502 S.n3428 S.n3423 0.024
R3503 S.n2942 S.n2937 0.024
R3504 S.n2433 S.n2428 0.024
R3505 S.n1912 S.n1907 0.024
R3506 S.n1367 S.n1362 0.024
R3507 S.n1417 S.n1393 0.024
R3508 S.n1962 S.n1938 0.024
R3509 S.n2483 S.n2459 0.024
R3510 S.n2992 S.n2968 0.024
R3511 S.n3478 S.n3454 0.024
R3512 S.n3952 S.n3928 0.024
R3513 S.n4475 S.n4459 0.024
R3514 S.n908 S.n907 0.024
R3515 S.n880 S.n879 0.024
R3516 S.n844 S.n843 0.024
R3517 S.n1228 S.n1227 0.024
R3518 S.n117 S.n116 0.024
R3519 S.n5064 S.n5063 0.023
R3520 S.n5258 S.n5245 0.023
R3521 S.n635 S.n630 0.023
R3522 S.n261 S.n260 0.023
R3523 S.n285 S.n281 0.023
R3524 S.n523 S.n520 0.023
R3525 S.n879 S.n878 0.023
R3526 S.t2 S.n118 0.023
R3527 S.n4641 S.n4640 0.023
R3528 S.n4459 S.n4458 0.023
R3529 S.n3928 S.n3927 0.023
R3530 S.n3454 S.n3453 0.023
R3531 S.n2968 S.n2967 0.023
R3532 S.n2459 S.n2458 0.023
R3533 S.n1938 S.n1937 0.023
R3534 S.n1393 S.n1392 0.023
R3535 S.n1417 S.n1397 0.023
R3536 S.n1962 S.n1942 0.023
R3537 S.n2483 S.n2463 0.023
R3538 S.n2992 S.n2972 0.023
R3539 S.n3478 S.n3458 0.023
R3540 S.n3952 S.n3932 0.023
R3541 S.n4475 S.n4463 0.023
R3542 S.n436 S.n434 0.023
R3543 S.n907 S.n906 0.023
R3544 S.n581 S.n580 0.023
R3545 S.n908 S.n904 0.023
R3546 S.n880 S.n876 0.023
R3547 S.n3558 S.n3557 0.023
R3548 S.n262 S.n258 0.023
R3549 S.n217 S.n216 0.023
R3550 S.n241 S.n237 0.023
R3551 S.n218 S.n214 0.023
R3552 S.n173 S.n172 0.023
R3553 S.n197 S.n193 0.023
R3554 S.n174 S.n170 0.023
R3555 S.n672 S.n670 0.023
R3556 S.n1226 S.n1225 0.023
R3557 S.n1234 S.n1232 0.023
R3558 S.n1795 S.n1794 0.023
R3559 S.n1812 S.n1810 0.023
R3560 S.n2345 S.n2344 0.023
R3561 S.n2362 S.n2360 0.023
R3562 S.n2886 S.n2885 0.023
R3563 S.n2903 S.n2901 0.023
R3564 S.n3401 S.n3400 0.023
R3565 S.n3418 S.n3416 0.023
R3566 S.n3907 S.n3906 0.023
R3567 S.n3924 S.n3922 0.023
R3568 S.n4385 S.n4384 0.023
R3569 S.n4402 S.n4400 0.023
R3570 S.n3423 S.n3421 0.023
R3571 S.n2937 S.n2934 0.023
R3572 S.n2428 S.n2426 0.023
R3573 S.n1907 S.n1904 0.023
R3574 S.n1362 S.n1359 0.023
R3575 S.n843 S.n840 0.023
R3576 S.n835 S.n834 0.023
R3577 S.n834 S.n833 0.022
R3578 S.n3947 S.n3943 0.022
R3579 S.n3473 S.n3469 0.022
R3580 S.n2987 S.n2983 0.022
R3581 S.n2478 S.n2474 0.022
R3582 S.n1957 S.n1953 0.022
R3583 S.n1412 S.n1408 0.022
R3584 S.n859 S.n855 0.022
R3585 S.n537 S.n533 0.022
R3586 S.n4867 S.n4866 0.022
R3587 S.n1804 S.n1802 0.022
R3588 S.n2354 S.n2352 0.022
R3589 S.n2895 S.n2893 0.022
R3590 S.n3410 S.n3408 0.022
R3591 S.n3916 S.n3914 0.022
R3592 S.n4394 S.n4392 0.022
R3593 S.n4031 S.n4030 0.022
R3594 S.n3540 S.n3538 0.022
R3595 S.n3068 S.n3067 0.022
R3596 S.n2545 S.n2543 0.022
R3597 S.n2038 S.n2037 0.022
R3598 S.n1480 S.n1478 0.022
R3599 S.n955 S.n954 0.022
R3600 S.n617 S.n615 0.022
R3601 S.n4871 S.n4870 0.022
R3602 S.n928 S.n927 0.021
R3603 S.n924 S.n923 0.021
R3604 S.n1465 S.n1464 0.021
R3605 S.n1463 S.n1462 0.021
R3606 S.n2009 S.n2008 0.021
R3607 S.n2007 S.n2006 0.021
R3608 S.n2530 S.n2529 0.021
R3609 S.n2528 S.n2527 0.021
R3610 S.n3039 S.n3038 0.021
R3611 S.n3037 S.n3036 0.021
R3612 S.n3525 S.n3524 0.021
R3613 S.n3523 S.n3522 0.021
R3614 S.n3999 S.n3998 0.021
R3615 S.n3997 S.n3996 0.021
R3616 S.n4443 S.n4442 0.021
R3617 S.n4441 S.n4440 0.021
R3618 S.n4852 S.n4851 0.021
R3619 S.n4850 S.n4849 0.021
R3620 S.n5339 S.n5338 0.021
R3621 S.n597 S.n596 0.021
R3622 S.n822 S.n821 0.021
R3623 S.n1378 S.n1377 0.021
R3624 S.n1376 S.n1375 0.021
R3625 S.n1923 S.n1922 0.021
R3626 S.n1921 S.n1920 0.021
R3627 S.n2444 S.n2443 0.021
R3628 S.n2442 S.n2441 0.021
R3629 S.n2953 S.n2952 0.021
R3630 S.n2951 S.n2950 0.021
R3631 S.n3439 S.n3438 0.021
R3632 S.n3437 S.n3436 0.021
R3633 S.n4025 S.n4024 0.021
R3634 S.n782 S.n781 0.021
R3635 S.n1316 S.n1315 0.021
R3636 S.n1314 S.n1313 0.021
R3637 S.n1862 S.n1861 0.021
R3638 S.n1860 S.n1859 0.021
R3639 S.n2383 S.n2382 0.021
R3640 S.n2381 S.n2380 0.021
R3641 S.n3062 S.n3061 0.021
R3642 S.n723 S.n722 0.021
R3643 S.n1255 S.n1254 0.021
R3644 S.n1253 S.n1252 0.021
R3645 S.n2032 S.n2031 0.021
R3646 S.n4644 S.n4643 0.021
R3647 S.n4835 S.n4834 0.021
R3648 S.n4426 S.n4425 0.021
R3649 S.n3982 S.n3981 0.021
R3650 S.n3508 S.n3507 0.021
R3651 S.n3022 S.n3021 0.021
R3652 S.n2513 S.n2512 0.021
R3653 S.n1992 S.n1991 0.021
R3654 S.n1448 S.n1447 0.021
R3655 S.n595 S.n594 0.021
R3656 S.n2366 S.n2365 0.021
R3657 S.n1845 S.n1844 0.021
R3658 S.n1299 S.n1298 0.021
R3659 S.n764 S.n763 0.021
R3660 S.n4032 S.n4031 0.021
R3661 S.n4474 S.n4473 0.021
R3662 S.n808 S.n807 0.021
R3663 S.n1346 S.n1345 0.021
R3664 S.n1892 S.n1891 0.021
R3665 S.n2413 S.n2412 0.021
R3666 S.n2922 S.n2921 0.021
R3667 S.n3542 S.n3540 0.021
R3668 S.n279 S.n278 0.021
R3669 S.n3069 S.n3068 0.021
R3670 S.n1238 S.n1237 0.021
R3671 S.n705 S.n704 0.021
R3672 S.n750 S.n749 0.021
R3673 S.n1285 S.n1284 0.021
R3674 S.n1831 S.n1830 0.021
R3675 S.n2547 S.n2545 0.021
R3676 S.n235 S.n234 0.021
R3677 S.n2039 S.n2038 0.021
R3678 S.n691 S.n690 0.021
R3679 S.n1482 S.n1480 0.021
R3680 S.n191 S.n190 0.021
R3681 S.n956 S.n955 0.021
R3682 S.n619 S.n617 0.021
R3683 S.n4830 S.n4829 0.021
R3684 S.n569 S.n568 0.02
R3685 S.n283 S.n282 0.02
R3686 S.n239 S.n238 0.02
R3687 S.n195 S.n194 0.02
R3688 S.n632 S.n631 0.02
R3689 S.n5313 S.n5312 0.02
R3690 S.n3423 S.n3422 0.02
R3691 S.n2937 S.n2936 0.02
R3692 S.n2428 S.n2427 0.02
R3693 S.n1907 S.n1906 0.02
R3694 S.n1362 S.n1361 0.02
R3695 S.n4032 S.n4028 0.02
R3696 S.n4868 S.n4865 0.02
R3697 S.n843 S.n842 0.02
R3698 S.n3542 S.n3541 0.02
R3699 S.n3069 S.n3065 0.02
R3700 S.n2547 S.n2546 0.02
R3701 S.n2039 S.n2035 0.02
R3702 S.n1482 S.n1481 0.02
R3703 S.n956 S.n952 0.02
R3704 S.n619 S.n618 0.02
R3705 S.n586 S.n585 0.02
R3706 S.t2 S.n104 0.019
R3707 S.n1109 S.n1107 0.019
R3708 S.n1632 S.n1630 0.019
R3709 S.n2228 S.n2226 0.019
R3710 S.n2753 S.n2751 0.019
R3711 S.n3252 S.n3250 0.019
R3712 S.n3620 S.n3618 0.019
R3713 S.n4206 S.n4204 0.019
R3714 S.n544 S.n543 0.019
R3715 S.n1128 S.n1127 0.019
R3716 S.n662 S.n661 0.019
R3717 S.n1221 S.n1220 0.019
R3718 S.n1784 S.n1783 0.019
R3719 S.n2334 S.n2333 0.019
R3720 S.n2875 S.n2874 0.019
R3721 S.n3390 S.n3389 0.019
R3722 S.n3896 S.n3895 0.019
R3723 S.n4374 S.n4373 0.019
R3724 S.n3951 S.n3950 0.019
R3725 S.n3477 S.n3476 0.019
R3726 S.n2991 S.n2990 0.019
R3727 S.n2482 S.n2481 0.019
R3728 S.n1961 S.n1960 0.019
R3729 S.n1416 S.n1415 0.019
R3730 S.n863 S.n862 0.019
R3731 S.n5018 S.n5017 0.019
R3732 S.n555 S.n554 0.018
R3733 S.n104 S.n103 0.018
R3734 S.n281 S.n280 0.018
R3735 S.n258 S.n257 0.018
R3736 S.n237 S.n236 0.018
R3737 S.n214 S.n213 0.018
R3738 S.n193 S.n192 0.018
R3739 S.n170 S.n169 0.018
R3740 S.n4783 S.n4782 0.018
R3741 S.n108 S.n107 0.018
R3742 S.n842 S.n841 0.018
R3743 S.n2936 S.n2935 0.018
R3744 S.n1906 S.n1905 0.018
R3745 S.n1361 S.n1360 0.018
R3746 S.n4780 S.n4779 0.017
R3747 S.n4787 S.n4784 0.017
R3748 S.n5255 S.n5254 0.017
R3749 S.n5254 S.n5253 0.017
R3750 S.n1807 S.n1806 0.017
R3751 S.n2357 S.n2356 0.017
R3752 S.n2898 S.n2897 0.017
R3753 S.n3413 S.n3412 0.017
R3754 S.n3919 S.n3918 0.017
R3755 S.n4397 S.n4396 0.017
R3756 S.n846 S.n835 0.016
R3757 S.n1096 S.n1092 0.016
R3758 S.n3561 S.n3553 0.016
R3759 S.n2566 S.n2558 0.016
R3760 S.n1501 S.n1493 0.016
R3761 S.n1805 S.n1804 0.016
R3762 S.n2355 S.n2354 0.016
R3763 S.n2896 S.n2895 0.016
R3764 S.n3411 S.n3410 0.016
R3765 S.n3917 S.n3916 0.016
R3766 S.n4395 S.n4394 0.016
R3767 S.n3421 S.n3420 0.015
R3768 S.n2426 S.n2425 0.015
R3769 S.n5218 S.n5217 0.015
R3770 S.n846 S.n845 0.015
R3771 S.n3949 S.n3948 0.015
R3772 S.n3948 S.n3947 0.015
R3773 S.n3947 S.n3946 0.015
R3774 S.n3475 S.n3474 0.015
R3775 S.n3474 S.n3473 0.015
R3776 S.n3473 S.n3472 0.015
R3777 S.n2989 S.n2988 0.015
R3778 S.n2988 S.n2987 0.015
R3779 S.n2987 S.n2986 0.015
R3780 S.n2480 S.n2479 0.015
R3781 S.n2479 S.n2478 0.015
R3782 S.n2478 S.n2477 0.015
R3783 S.n1959 S.n1958 0.015
R3784 S.n1958 S.n1957 0.015
R3785 S.n1957 S.n1956 0.015
R3786 S.n1414 S.n1413 0.015
R3787 S.n1413 S.n1412 0.015
R3788 S.n1412 S.n1411 0.015
R3789 S.n861 S.n860 0.015
R3790 S.n860 S.n859 0.015
R3791 S.n859 S.n858 0.015
R3792 S.n538 S.n537 0.015
R3793 S.n537 S.n536 0.015
R3794 S.n4870 S.n4869 0.015
R3795 S.n584 S.n583 0.015
R3796 S.n1808 S.n1788 0.015
R3797 S.n2358 S.n2338 0.015
R3798 S.n2899 S.n2879 0.015
R3799 S.n3414 S.n3394 0.015
R3800 S.n3920 S.n3900 0.015
R3801 S.n4398 S.n4378 0.015
R3802 S.n5016 S.n5015 0.015
R3803 S.n5015 S.n5014 0.015
R3804 S.n4782 S.n4781 0.015
R3805 S.n4831 S.n4826 0.015
R3806 S.n4838 S.n4837 0.015
R3807 S.n4429 S.n4428 0.015
R3808 S.n3985 S.n3984 0.015
R3809 S.n3511 S.n3510 0.015
R3810 S.n3025 S.n3024 0.015
R3811 S.n2516 S.n2515 0.015
R3812 S.n1995 S.n1994 0.015
R3813 S.n1451 S.n1450 0.015
R3814 S.n2369 S.n2368 0.015
R3815 S.n1848 S.n1847 0.015
R3816 S.n1302 S.n1301 0.015
R3817 S.n767 S.n766 0.015
R3818 S.n2917 S.n2916 0.015
R3819 S.n2408 S.n2407 0.015
R3820 S.n1887 S.n1886 0.015
R3821 S.n1341 S.n1340 0.015
R3822 S.n804 S.n803 0.015
R3823 S.n1241 S.n1240 0.015
R3824 S.n708 S.n707 0.015
R3825 S.n1826 S.n1825 0.015
R3826 S.n1280 S.n1279 0.015
R3827 S.n745 S.n744 0.015
R3828 S.n686 S.n685 0.015
R3829 S.n541 S.n540 0.014
R3830 S.n4820 S.n4818 0.014
R3831 S.n771 S.n770 0.014
R3832 S.n1349 S.n1348 0.014
R3833 S.n1895 S.n1894 0.014
R3834 S.n2416 S.n2415 0.014
R3835 S.n2925 S.n2924 0.014
R3836 S.n712 S.n711 0.014
R3837 S.n1288 S.n1287 0.014
R3838 S.n1834 S.n1833 0.014
R3839 S.n5483 S.n5474 0.014
R3840 S.n5230 S.n5220 0.014
R3841 S.n845 S.n844 0.014
R3842 S.n1073 S.n1072 0.014
R3843 S.n1714 S.n1713 0.014
R3844 S.n2295 S.n2294 0.014
R3845 S.n2836 S.n2835 0.014
R3846 S.n3354 S.n3353 0.014
R3847 S.n3750 S.n3749 0.014
R3848 S.n4337 S.n4336 0.014
R3849 S.n5070 S.n5069 0.014
R3850 S.n4842 S.n4841 0.013
R3851 S.n4433 S.n4432 0.013
R3852 S.n3989 S.n3988 0.013
R3853 S.n3515 S.n3514 0.013
R3854 S.n3029 S.n3028 0.013
R3855 S.n2520 S.n2519 0.013
R3856 S.n1999 S.n1998 0.013
R3857 S.n1455 S.n1454 0.013
R3858 S.n2373 S.n2372 0.013
R3859 S.n1852 S.n1851 0.013
R3860 S.n1306 S.n1305 0.013
R3861 S.n811 S.n810 0.013
R3862 S.n1245 S.n1244 0.013
R3863 S.n753 S.n752 0.013
R3864 S.n694 S.n693 0.013
R3865 S.n4472 S.n4471 0.013
R3866 S.n1713 S.n1712 0.013
R3867 S.n2294 S.n2293 0.013
R3868 S.n2835 S.n2834 0.013
R3869 S.n3353 S.n3352 0.013
R3870 S.n3749 S.n3748 0.013
R3871 S.n4336 S.n4335 0.013
R3872 S.n5069 S.n5068 0.013
R3873 S.t2 S.n0 0.012
R3874 S.t2 S.n8 0.012
R3875 S.t2 S.n16 0.012
R3876 S.t2 S.n33 0.012
R3877 S.n4826 S.n4822 0.012
R3878 S.n5251 S.n5250 0.012
R3879 S.n4839 S.n4838 0.012
R3880 S.n4430 S.n4429 0.012
R3881 S.n3986 S.n3985 0.012
R3882 S.n3512 S.n3511 0.012
R3883 S.n3026 S.n3025 0.012
R3884 S.n2517 S.n2516 0.012
R3885 S.n1996 S.n1995 0.012
R3886 S.n1452 S.n1451 0.012
R3887 S.n608 S.n599 0.012
R3888 S.n2370 S.n2369 0.012
R3889 S.n1849 S.n1848 0.012
R3890 S.n1303 S.n1302 0.012
R3891 S.n768 S.n767 0.012
R3892 S.n2918 S.n2917 0.012
R3893 S.n2409 S.n2408 0.012
R3894 S.n1888 S.n1887 0.012
R3895 S.n1342 S.n1341 0.012
R3896 S.n838 S.n837 0.012
R3897 S.n3426 S.n3425 0.012
R3898 S.n2940 S.n2939 0.012
R3899 S.n2431 S.n2430 0.012
R3900 S.n1910 S.n1909 0.012
R3901 S.n1365 S.n1364 0.012
R3902 S.n805 S.n804 0.012
R3903 S.n294 S.n285 0.012
R3904 S.n1242 S.n1241 0.012
R3905 S.n709 S.n708 0.012
R3906 S.n1827 S.n1826 0.012
R3907 S.n1281 S.n1280 0.012
R3908 S.n746 S.n745 0.012
R3909 S.n250 S.n241 0.012
R3910 S.n687 S.n686 0.012
R3911 S.n206 S.n197 0.012
R3912 S.n1712 S.n1711 0.012
R3913 S.n1802 S.n1801 0.012
R3914 S.n2293 S.n2292 0.012
R3915 S.n2352 S.n2351 0.012
R3916 S.n2834 S.n2833 0.012
R3917 S.n2893 S.n2892 0.012
R3918 S.n3352 S.n3351 0.012
R3919 S.n3408 S.n3407 0.012
R3920 S.n3748 S.n3747 0.012
R3921 S.n3914 S.n3913 0.012
R3922 S.n4335 S.n4334 0.012
R3923 S.n4392 S.n4391 0.012
R3924 S.n5068 S.n5067 0.012
R3925 S.n4787 S.n4780 0.01
R3926 S.n410 S.n409 0.01
R3927 S.n377 S.n376 0.01
R3928 S.n344 S.n343 0.01
R3929 S.n4014 S.n4013 0.01
R3930 S.n525 S.n523 0.01
R3931 S.n1117 S.n1109 0.01
R3932 S.n1640 S.n1632 0.01
R3933 S.n2236 S.n2228 0.01
R3934 S.n2761 S.n2753 0.01
R3935 S.n3260 S.n3252 0.01
R3936 S.n3628 S.n3620 0.01
R3937 S.n4214 S.n4206 0.01
R3938 S.n439 S.n436 0.01
R3939 S.n4665 S.n4661 0.01
R3940 S.n4234 S.n4230 0.01
R3941 S.n3648 S.n3644 0.01
R3942 S.n3280 S.n3276 0.01
R3943 S.n2781 S.n2777 0.01
R3944 S.n2256 S.n2252 0.01
R3945 S.n1660 S.n1656 0.01
R3946 S.n1137 S.n1128 0.01
R3947 S.n587 S.n586 0.01
R3948 S.n458 S.n455 0.01
R3949 S.n262 S.n261 0.01
R3950 S.n218 S.n217 0.01
R3951 S.n174 S.n173 0.01
R3952 S.n493 S.n491 0.01
R3953 S.n1229 S.n1226 0.01
R3954 S.n1229 S.n672 0.01
R3955 S.n1808 S.n1234 0.01
R3956 S.n2358 S.n1812 0.01
R3957 S.n2899 S.n2362 0.01
R3958 S.n3414 S.n2903 0.01
R3959 S.n3920 S.n3418 0.01
R3960 S.n4398 S.n3924 0.01
R3961 S.n4831 S.n4402 0.01
R3962 S.n5260 S.n5258 0.01
R3963 S.n558 S.n541 0.01
R3964 S.n285 S.n284 0.01
R3965 S.n241 S.n240 0.01
R3966 S.n197 S.n196 0.01
R3967 S.n5253 S.n5251 0.01
R3968 S.n1095 S.n1093 0.01
R3969 S.n260 S.n259 0.01
R3970 S.n216 S.n215 0.01
R3971 S.n172 S.n171 0.01
R3972 S.n4646 S.n4644 0.01
R3973 S.n3589 S.n3574 0.01
R3974 S.n2686 S.n2671 0.01
R3975 S.n1529 S.n1514 0.01
R3976 S.n5498 S.n5309 0.009
R3977 S.n5256 S.n5255 0.009
R3978 S.n4475 S.n4474 0.009
R3979 S.n5260 S.n5244 0.009
R3980 S.n4840 S.n4839 0.008
R3981 S.n4431 S.n4430 0.008
R3982 S.n3987 S.n3986 0.008
R3983 S.n3513 S.n3512 0.008
R3984 S.n3027 S.n3026 0.008
R3985 S.n2518 S.n2517 0.008
R3986 S.n1997 S.n1996 0.008
R3987 S.n1453 S.n1452 0.008
R3988 S.n2371 S.n2370 0.008
R3989 S.n1850 S.n1849 0.008
R3990 S.n1304 S.n1303 0.008
R3991 S.n769 S.n768 0.008
R3992 S.n2919 S.n2918 0.008
R3993 S.n2410 S.n2409 0.008
R3994 S.n1889 S.n1888 0.008
R3995 S.n1343 S.n1342 0.008
R3996 S.n806 S.n805 0.008
R3997 S.n1243 S.n1242 0.008
R3998 S.n710 S.n709 0.008
R3999 S.n1828 S.n1827 0.008
R4000 S.n1282 S.n1281 0.008
R4001 S.n747 S.n746 0.008
R4002 S.n688 S.n687 0.008
R4003 S.n932 S.n931 0.008
R4004 S.n1155 S.n1154 0.008
R4005 S.n1469 S.n1468 0.008
R4006 S.n1678 S.n1677 0.008
R4007 S.n2013 S.n2012 0.008
R4008 S.n2274 S.n2273 0.008
R4009 S.n2534 S.n2533 0.008
R4010 S.n2799 S.n2798 0.008
R4011 S.n3043 S.n3042 0.008
R4012 S.n3298 S.n3297 0.008
R4013 S.n3529 S.n3528 0.008
R4014 S.n3666 S.n3665 0.008
R4015 S.n4003 S.n4002 0.008
R4016 S.n4252 S.n4251 0.008
R4017 S.n4447 S.n4446 0.008
R4018 S.n4683 S.n4682 0.008
R4019 S.n4856 S.n4855 0.008
R4020 S.n5046 S.n5045 0.008
R4021 S.n926 S.n925 0.008
R4022 S.n820 S.n819 0.008
R4023 S.n1082 S.n1081 0.008
R4024 S.n1382 S.n1381 0.008
R4025 S.n1618 S.n1617 0.008
R4026 S.n1927 S.n1926 0.008
R4027 S.n2214 S.n2213 0.008
R4028 S.n2448 S.n2447 0.008
R4029 S.n2739 S.n2738 0.008
R4030 S.n2957 S.n2956 0.008
R4031 S.n3238 S.n3237 0.008
R4032 S.n3443 S.n3442 0.008
R4033 S.n3606 S.n3605 0.008
R4034 S.n1117 S.n1106 0.008
R4035 S.n1640 S.n1629 0.008
R4036 S.n2236 S.n2225 0.008
R4037 S.n2761 S.n2750 0.008
R4038 S.n3260 S.n3249 0.008
R4039 S.n3628 S.n3617 0.008
R4040 S.n4214 S.n4203 0.008
R4041 S.n439 S.n438 0.008
R4042 S.n4665 S.n4664 0.008
R4043 S.n4234 S.n4233 0.008
R4044 S.n3648 S.n3647 0.008
R4045 S.n3280 S.n3279 0.008
R4046 S.n2781 S.n2780 0.008
R4047 S.n2256 S.n2255 0.008
R4048 S.n1660 S.n1659 0.008
R4049 S.n1137 S.n1126 0.008
R4050 S.n888 S.n887 0.008
R4051 S.n1425 S.n1424 0.008
R4052 S.n1970 S.n1969 0.008
R4053 S.n2491 S.n2490 0.008
R4054 S.n3000 S.n2999 0.008
R4055 S.n3486 S.n3485 0.008
R4056 S.n3960 S.n3959 0.008
R4057 S.n4404 S.n4403 0.008
R4058 S.n567 S.n566 0.008
R4059 S.n583 S.n581 0.008
R4060 S.n583 S.n582 0.008
R4061 S.n458 S.n457 0.008
R4062 S.n3560 S.n3558 0.008
R4063 S.n2905 S.n2904 0.008
R4064 S.n2396 S.n2395 0.008
R4065 S.n1875 S.n1874 0.008
R4066 S.n1329 S.n1328 0.008
R4067 S.n793 S.n792 0.008
R4068 S.n783 S.n780 0.008
R4069 S.n1054 S.n1053 0.008
R4070 S.n1320 S.n1319 0.008
R4071 S.n1582 S.n1581 0.008
R4072 S.n1866 S.n1865 0.008
R4073 S.n2181 S.n2180 0.008
R4074 S.n2387 S.n2386 0.008
R4075 S.n2703 S.n2702 0.008
R4076 S.n2565 S.n2561 0.008
R4077 S.n1814 S.n1813 0.008
R4078 S.n1268 S.n1267 0.008
R4079 S.n734 S.n733 0.008
R4080 S.n724 S.n721 0.008
R4081 S.n1018 S.n1017 0.008
R4082 S.n1259 S.n1258 0.008
R4083 S.n1546 S.n1545 0.008
R4084 S.n1500 S.n1496 0.008
R4085 S.n675 S.n674 0.008
R4086 S.n637 S.n636 0.008
R4087 S.n493 S.n492 0.008
R4088 S.n668 S.n166 0.008
R4089 S.n4787 S.n4786 0.008
R4090 S.n5311 S.n5310 0.008
R4091 S.n557 S.n556 0.008
R4092 S.n557 S.n555 0.007
R4093 S.t2 S.n96 0.007
R4094 S.t2 S.n89 0.007
R4095 S.t2 S.n77 0.007
R4096 S.t2 S.n65 0.007
R4097 S.n540 S.n539 0.007
R4098 S.n4779 S.n4778 0.007
R4099 S.n927 S.n926 0.006
R4100 S.n783 S.n782 0.006
R4101 S.n724 S.n723 0.006
R4102 S.n5312 S.n5311 0.006
R4103 S.n271 S.n262 0.006
R4104 S.n227 S.n218 0.006
R4105 S.n186 S.n174 0.006
R4106 S.n525 S.n512 0.005
R4107 S.n839 S.n838 0.005
R4108 S.n3427 S.n3426 0.005
R4109 S.n2941 S.n2940 0.005
R4110 S.n2432 S.n2431 0.005
R4111 S.n1911 S.n1910 0.005
R4112 S.n1366 S.n1365 0.005
R4113 S.t2 S.n101 0.005
R4114 S.n3555 S.n3554 0.005
R4115 S.n2560 S.n2559 0.005
R4116 S.n1495 S.n1494 0.005
R4117 S.t2 S.n115 0.005
R4118 S.n5321 S.n5320 0.004
R4119 S.n5062 S.n5061 0.004
R4120 S.n5243 S.n5242 0.004
R4121 S.n629 S.n628 0.004
R4122 S.n606 S.n605 0.004
R4123 S.n919 S.n918 0.004
R4124 S.n5334 S.n5333 0.004
R4125 S.n5039 S.n5038 0.004
R4126 S.n4845 S.n4844 0.004
R4127 S.n4676 S.n4675 0.004
R4128 S.n4436 S.n4435 0.004
R4129 S.n4245 S.n4244 0.004
R4130 S.n3992 S.n3991 0.004
R4131 S.n3659 S.n3658 0.004
R4132 S.n3518 S.n3517 0.004
R4133 S.n3291 S.n3290 0.004
R4134 S.n3032 S.n3031 0.004
R4135 S.n2792 S.n2791 0.004
R4136 S.n2523 S.n2522 0.004
R4137 S.n2267 S.n2266 0.004
R4138 S.n2002 S.n2001 0.004
R4139 S.n1671 S.n1670 0.004
R4140 S.n1458 S.n1457 0.004
R4141 S.n1148 S.n1147 0.004
R4142 S.n473 S.n472 0.004
R4143 S.n269 S.n268 0.004
R4144 S.n774 S.n773 0.004
R4145 S.n3056 S.n3055 0.004
R4146 S.n2696 S.n2695 0.004
R4147 S.n2376 S.n2375 0.004
R4148 S.n2174 S.n2173 0.004
R4149 S.n1855 S.n1854 0.004
R4150 S.n1575 S.n1574 0.004
R4151 S.n1309 S.n1308 0.004
R4152 S.n1047 S.n1046 0.004
R4153 S.n292 S.n291 0.004
R4154 S.n3552 S.n3551 0.004
R4155 S.n3218 S.n3217 0.004
R4156 S.n2915 S.n2914 0.004
R4157 S.n2719 S.n2718 0.004
R4158 S.n2406 S.n2405 0.004
R4159 S.n2194 S.n2193 0.004
R4160 S.n1885 S.n1884 0.004
R4161 S.n1598 S.n1597 0.004
R4162 S.n1339 S.n1338 0.004
R4163 S.n1070 S.n1069 0.004
R4164 S.n1091 S.n1090 0.004
R4165 S.n831 S.n830 0.004
R4166 S.n508 S.n507 0.004
R4167 S.n519 S.n518 0.004
R4168 S.n1371 S.n1370 0.004
R4169 S.n1916 S.n1915 0.004
R4170 S.n2437 S.n2436 0.004
R4171 S.n2946 S.n2945 0.004
R4172 S.n3432 S.n3431 0.004
R4173 S.n4019 S.n4018 0.004
R4174 S.n3599 S.n3598 0.004
R4175 S.n3231 S.n3230 0.004
R4176 S.n2732 S.n2731 0.004
R4177 S.n2207 S.n2206 0.004
R4178 S.n1611 S.n1610 0.004
R4179 S.n870 S.n869 0.004
R4180 S.n433 S.n432 0.004
R4181 S.n551 S.n550 0.004
R4182 S.n4467 S.n4466 0.004
R4183 S.n4209 S.n4208 0.004
R4184 S.n3937 S.n3936 0.004
R4185 S.n3623 S.n3622 0.004
R4186 S.n3463 S.n3462 0.004
R4187 S.n3255 S.n3254 0.004
R4188 S.n2977 S.n2976 0.004
R4189 S.n2756 S.n2755 0.004
R4190 S.n2468 S.n2467 0.004
R4191 S.n2231 S.n2230 0.004
R4192 S.n1947 S.n1946 0.004
R4193 S.n1635 S.n1634 0.004
R4194 S.n1402 S.n1401 0.004
R4195 S.n1112 S.n1111 0.004
R4196 S.n898 S.n897 0.004
R4197 S.n453 S.n452 0.004
R4198 S.n1131 S.n1130 0.004
R4199 S.n1435 S.n1434 0.004
R4200 S.n1655 S.n1654 0.004
R4201 S.n1980 S.n1979 0.004
R4202 S.n2251 S.n2250 0.004
R4203 S.n2501 S.n2500 0.004
R4204 S.n2776 S.n2775 0.004
R4205 S.n3010 S.n3009 0.004
R4206 S.n3275 S.n3274 0.004
R4207 S.n3496 S.n3495 0.004
R4208 S.n3643 S.n3642 0.004
R4209 S.n3970 S.n3969 0.004
R4210 S.n4229 S.n4228 0.004
R4211 S.n4414 S.n4413 0.004
R4212 S.n4660 S.n4659 0.004
R4213 S.n4879 S.n4878 0.004
R4214 S.n577 S.n576 0.004
R4215 S.n802 S.n801 0.004
R4216 S.n417 S.n416 0.004
R4217 S.n400 S.n399 0.004
R4218 S.n225 S.n224 0.004
R4219 S.n715 S.n714 0.004
R4220 S.n2026 S.n2025 0.004
R4221 S.n1539 S.n1538 0.004
R4222 S.n1248 S.n1247 0.004
R4223 S.n1011 S.n1010 0.004
R4224 S.n248 S.n247 0.004
R4225 S.n2557 S.n2556 0.004
R4226 S.n2158 S.n2157 0.004
R4227 S.n1824 S.n1823 0.004
R4228 S.n1562 S.n1561 0.004
R4229 S.n1278 S.n1277 0.004
R4230 S.n1034 S.n1033 0.004
R4231 S.n743 S.n742 0.004
R4232 S.n384 S.n383 0.004
R4233 S.n367 S.n366 0.004
R4234 S.n184 S.n183 0.004
R4235 S.n945 S.n944 0.004
R4236 S.n204 S.n203 0.004
R4237 S.n1492 S.n1491 0.004
R4238 S.n998 S.n997 0.004
R4239 S.n684 S.n683 0.004
R4240 S.n351 S.n350 0.004
R4241 S.n334 S.n333 0.004
R4242 S.n651 S.n650 0.004
R4243 S.n490 S.n489 0.004
R4244 S.n1199 S.n1198 0.004
R4245 S.n1188 S.n1187 0.004
R4246 S.n1742 S.n1741 0.004
R4247 S.n1730 S.n1729 0.004
R4248 S.n2071 S.n2070 0.004
R4249 S.n2059 S.n2058 0.004
R4250 S.n2597 S.n2596 0.004
R4251 S.n2585 S.n2584 0.004
R4252 S.n3101 S.n3100 0.004
R4253 S.n3089 S.n3088 0.004
R4254 S.n3778 S.n3777 0.004
R4255 S.n3766 S.n3765 0.004
R4256 S.n4064 S.n4063 0.004
R4257 S.n4052 S.n4051 0.004
R4258 S.n4506 S.n4505 0.004
R4259 S.n4494 S.n4493 0.004
R4260 S.n4895 S.n4894 0.004
R4261 S.n5084 S.n5083 0.004
R4262 S.n5355 S.n5354 0.004
R4263 S.n1215 S.n1214 0.004
R4264 S.n1171 S.n1170 0.004
R4265 S.n1759 S.n1758 0.004
R4266 S.n5371 S.n5370 0.004
R4267 S.n5099 S.n5098 0.004
R4268 S.n4912 S.n4911 0.004
R4269 S.n4531 S.n4530 0.004
R4270 S.n4523 S.n4522 0.004
R4271 S.n4089 S.n4088 0.004
R4272 S.n4081 S.n4080 0.004
R4273 S.n3803 S.n3802 0.004
R4274 S.n3795 S.n3794 0.004
R4275 S.n3126 S.n3125 0.004
R4276 S.n3118 S.n3117 0.004
R4277 S.n2622 S.n2621 0.004
R4278 S.n2614 S.n2613 0.004
R4279 S.n2096 S.n2095 0.004
R4280 S.n2088 S.n2087 0.004
R4281 S.n1691 S.n1690 0.004
R4282 S.n1776 S.n1775 0.004
R4283 S.n1709 S.n1708 0.004
R4284 S.n2119 S.n2118 0.004
R4285 S.n5386 S.n5385 0.004
R4286 S.n5114 S.n5113 0.004
R4287 S.n4928 S.n4927 0.004
R4288 S.n4695 S.n4694 0.004
R4289 S.n4554 S.n4553 0.004
R4290 S.n4265 S.n4264 0.004
R4291 S.n4112 S.n4111 0.004
R4292 S.n3679 S.n3678 0.004
R4293 S.n3826 S.n3825 0.004
R4294 S.n3311 S.n3310 0.004
R4295 S.n3149 S.n3148 0.004
R4296 S.n2812 S.n2811 0.004
R4297 S.n2645 S.n2644 0.004
R4298 S.n2127 S.n2126 0.004
R4299 S.n2326 S.n2325 0.004
R4300 S.n2290 S.n2289 0.004
R4301 S.n2660 S.n2659 0.004
R4302 S.n5401 S.n5400 0.004
R4303 S.n5130 S.n5129 0.004
R4304 S.n4943 S.n4942 0.004
R4305 S.n4711 S.n4710 0.004
R4306 S.n4569 S.n4568 0.004
R4307 S.n4281 S.n4280 0.004
R4308 S.n4127 S.n4126 0.004
R4309 S.n3695 S.n3694 0.004
R4310 S.n3841 S.n3840 0.004
R4311 S.n3327 S.n3326 0.004
R4312 S.n3164 S.n3163 0.004
R4313 S.n2668 S.n2667 0.004
R4314 S.n2867 S.n2866 0.004
R4315 S.n2831 S.n2830 0.004
R4316 S.n3179 S.n3178 0.004
R4317 S.n5416 S.n5415 0.004
R4318 S.n5146 S.n5145 0.004
R4319 S.n4958 S.n4957 0.004
R4320 S.n4727 S.n4726 0.004
R4321 S.n4584 S.n4583 0.004
R4322 S.n4297 S.n4296 0.004
R4323 S.n4142 S.n4141 0.004
R4324 S.n3711 S.n3710 0.004
R4325 S.n3856 S.n3855 0.004
R4326 S.n3187 S.n3186 0.004
R4327 S.n3382 S.n3381 0.004
R4328 S.n3349 S.n3348 0.004
R4329 S.n3871 S.n3870 0.004
R4330 S.n5431 S.n5430 0.004
R4331 S.n5162 S.n5161 0.004
R4332 S.n4973 S.n4972 0.004
R4333 S.n4743 S.n4742 0.004
R4334 S.n4599 S.n4598 0.004
R4335 S.n4313 S.n4312 0.004
R4336 S.n4157 S.n4156 0.004
R4337 S.n3727 S.n3726 0.004
R4338 S.n3888 S.n3887 0.004
R4339 S.n3745 S.n3744 0.004
R4340 S.n4172 S.n4171 0.004
R4341 S.n5446 S.n5445 0.004
R4342 S.n5178 S.n5177 0.004
R4343 S.n4988 S.n4987 0.004
R4344 S.n4759 S.n4758 0.004
R4345 S.n4614 S.n4613 0.004
R4346 S.n4180 S.n4179 0.004
R4347 S.n4368 S.n4367 0.004
R4348 S.n4332 S.n4331 0.004
R4349 S.n4629 S.n4628 0.004
R4350 S.n5461 S.n5460 0.004
R4351 S.n5194 S.n5193 0.004
R4352 S.n5003 S.n5002 0.004
R4353 S.n4637 S.n4636 0.004
R4354 S.n4817 S.n4816 0.004
R4355 S.n4776 S.n4775 0.004
R4356 S.n5227 S.n5226 0.004
R4357 S.n5481 S.n5480 0.004
R4358 S.n5214 S.n5213 0.004
R4359 S.n5496 S.n5495 0.004
R4360 S.t2 S.n108 0.004
R4361 S.n608 S.n607 0.004
R4362 S.n294 S.n293 0.004
R4363 S.n271 S.n270 0.004
R4364 S.n250 S.n249 0.004
R4365 S.n227 S.n226 0.004
R4366 S.n206 S.n205 0.004
R4367 S.n186 S.n185 0.004
R4368 S.t2 S.n124 0.004
R4369 S.n321 S.n306 0.004
R4370 S.n4194 S.n4193 0.004
R4371 S.n3943 S.n3942 0.004
R4372 S.n3469 S.n3468 0.004
R4373 S.n2983 S.n2982 0.004
R4374 S.n2474 S.n2473 0.004
R4375 S.n1953 S.n1952 0.004
R4376 S.n1408 S.n1407 0.004
R4377 S.n855 S.n854 0.004
R4378 S.n533 S.n532 0.004
R4379 S.n4194 S.n4192 0.004
R4380 S.n458 S.n446 0.004
R4381 S.n1137 S.n1136 0.004
R4382 S.n1660 S.n1648 0.004
R4383 S.n2256 S.n2244 0.004
R4384 S.n2781 S.n2769 0.004
R4385 S.n3280 S.n3268 0.004
R4386 S.n3648 S.n3636 0.004
R4387 S.n4234 S.n4222 0.004
R4388 S.n4665 S.n4653 0.004
R4389 S.n5029 S.n5027 0.004
R4390 S.n3589 S.n3588 0.004
R4391 S.n419 S.n410 0.004
R4392 S.n3204 S.n3202 0.004
R4393 S.n2686 S.n2685 0.004
R4394 S.n386 S.n377 0.004
R4395 S.n2144 S.n2142 0.004
R4396 S.n1529 S.n1528 0.004
R4397 S.n353 S.n344 0.004
R4398 S.n984 S.n982 0.004
R4399 S.n321 S.n320 0.004
R4400 S.n837 S.n836 0.004
R4401 S.n3425 S.n3424 0.004
R4402 S.n2939 S.n2938 0.004
R4403 S.n2430 S.n2429 0.004
R4404 S.n1909 S.n1908 0.004
R4405 S.n1364 S.n1363 0.004
R4406 S.n4646 S.n4641 0.004
R4407 S.n3951 S.n3949 0.004
R4408 S.n3477 S.n3475 0.004
R4409 S.n2991 S.n2989 0.004
R4410 S.n2482 S.n2480 0.004
R4411 S.n1961 S.n1959 0.004
R4412 S.n1416 S.n1414 0.004
R4413 S.n863 S.n861 0.004
R4414 S.n1096 S.n1095 0.004
R4415 S.n3561 S.n3560 0.004
R4416 S.n3589 S.n3573 0.004
R4417 S.n2566 S.n2565 0.004
R4418 S.n2686 S.n2670 0.004
R4419 S.n1501 S.n1500 0.004
R4420 S.n1529 S.n1513 0.004
R4421 S.n1807 S.n1793 0.004
R4422 S.n1808 S.n1807 0.004
R4423 S.n2357 S.n2343 0.004
R4424 S.n2358 S.n2357 0.004
R4425 S.n2898 S.n2884 0.004
R4426 S.n2899 S.n2898 0.004
R4427 S.n3413 S.n3399 0.004
R4428 S.n3414 S.n3413 0.004
R4429 S.n3919 S.n3905 0.004
R4430 S.n3920 S.n3919 0.004
R4431 S.n4397 S.n4383 0.004
R4432 S.n4398 S.n4397 0.004
R4433 S.n5018 S.n5016 0.004
R4434 S.n4822 S.n4821 0.004
R4435 S.n4831 S.n4830 0.004
R4436 S.t0 S.n5303 0.004
R4437 S.t0 S.n5305 0.004
R4438 S.t12 S.n324 0.004
R4439 S.t2 S.n142 0.004
R4440 S.t2 S.n139 0.004
R4441 S.t2 S.n91 0.004
R4442 S.t95 S.n3207 0.004
R4443 S.t2 S.n154 0.004
R4444 S.t53 S.n3592 0.004
R4445 S.t2 S.n106 0.004
R4446 S.t66 S.n4197 0.004
R4447 S.t2 S.n120 0.004
R4448 S.t31 S.n4649 0.004
R4449 S.t44 S.n5032 0.004
R4450 S.t2 S.n130 0.004
R4451 S.t2 S.n79 0.004
R4452 S.t8 S.n2147 0.004
R4453 S.t2 S.n150 0.004
R4454 S.t168 S.n2689 0.004
R4455 S.t2 S.n67 0.004
R4456 S.t151 S.n987 0.004
R4457 S.t2 S.n146 0.004
R4458 S.t42 S.n1532 0.004
R4459 S.t2 S.n54 0.004
R4460 S.t0 S.n5267 0.004
R4461 S.t0 S.n5271 0.004
R4462 S.t0 S.n5275 0.004
R4463 S.t0 S.n5279 0.004
R4464 S.t0 S.n5283 0.004
R4465 S.t0 S.n5287 0.004
R4466 S.t0 S.n5291 0.004
R4467 S.t0 S.n5295 0.004
R4468 S.t0 S.n5299 0.004
R4469 S.t0 S.n5264 0.004
R4470 S.t2 S.n137 0.004
R4471 S.t2 S.n7 0.004
R4472 S.t2 S.n15 0.004
R4473 S.t2 S.n24 0.004
R4474 S.t2 S.n28 0.004
R4475 S.n510 S.n509 0.004
R4476 S.t2 S.n134 0.004
R4477 S.t2 S.n83 0.004
R4478 S.t2 S.n71 0.004
R4479 S.t2 S.n58 0.004
R4480 S.n5029 S.n5028 0.004
R4481 S.n3607 S.n3596 0.004
R4482 S.n3239 S.n3228 0.004
R4483 S.n2740 S.n2729 0.004
R4484 S.n2215 S.n2204 0.004
R4485 S.n1619 S.n1608 0.004
R4486 S.n5329 S.n5328 0.003
R4487 S.n5077 S.n5076 0.003
R4488 S.n5239 S.n5238 0.003
R4489 S.n641 S.n640 0.003
R4490 S.n614 S.n613 0.003
R4491 S.n939 S.n938 0.003
R4492 S.n5345 S.n5344 0.003
R4493 S.n5053 S.n5052 0.003
R4494 S.n4863 S.n4862 0.003
R4495 S.n4690 S.n4689 0.003
R4496 S.n4454 S.n4453 0.003
R4497 S.n4259 S.n4258 0.003
R4498 S.n4010 S.n4009 0.003
R4499 S.n3673 S.n3672 0.003
R4500 S.n3536 S.n3535 0.003
R4501 S.n3305 S.n3304 0.003
R4502 S.n3050 S.n3049 0.003
R4503 S.n2806 S.n2805 0.003
R4504 S.n2541 S.n2540 0.003
R4505 S.n2281 S.n2280 0.003
R4506 S.n2020 S.n2019 0.003
R4507 S.n1685 S.n1684 0.003
R4508 S.n1476 S.n1475 0.003
R4509 S.n1162 S.n1161 0.003
R4510 S.n481 S.n480 0.003
R4511 S.n277 S.n276 0.003
R4512 S.n790 S.n789 0.003
R4513 S.n3073 S.n3072 0.003
R4514 S.n2710 S.n2709 0.003
R4515 S.n2394 S.n2393 0.003
R4516 S.n2185 S.n2184 0.003
R4517 S.n1873 S.n1872 0.003
R4518 S.n1589 S.n1588 0.003
R4519 S.n1327 S.n1326 0.003
R4520 S.n1061 S.n1060 0.003
R4521 S.n300 S.n299 0.003
R4522 S.n3564 S.n3563 0.003
R4523 S.n3226 S.n3225 0.003
R4524 S.n2932 S.n2931 0.003
R4525 S.n2727 S.n2726 0.003
R4526 S.n2423 S.n2422 0.003
R4527 S.n2202 S.n2201 0.003
R4528 S.n1902 S.n1901 0.003
R4529 S.n1606 S.n1605 0.003
R4530 S.n1356 S.n1355 0.003
R4531 S.n1080 S.n1079 0.003
R4532 S.n1102 S.n1101 0.003
R4533 S.n852 S.n851 0.003
R4534 S.n502 S.n501 0.003
R4535 S.n531 S.n530 0.003
R4536 S.n1389 S.n1388 0.003
R4537 S.n1934 S.n1933 0.003
R4538 S.n2455 S.n2454 0.003
R4539 S.n2964 S.n2963 0.003
R4540 S.n3450 S.n3449 0.003
R4541 S.n4036 S.n4035 0.003
R4542 S.n3613 S.n3612 0.003
R4543 S.n3245 S.n3244 0.003
R4544 S.n2746 S.n2745 0.003
R4545 S.n2221 S.n2220 0.003
R4546 S.n1625 S.n1624 0.003
R4547 S.n886 S.n885 0.003
R4548 S.n445 S.n444 0.003
R4549 S.n564 S.n563 0.003
R4550 S.n4478 S.n4477 0.003
R4551 S.n4220 S.n4219 0.003
R4552 S.n3958 S.n3957 0.003
R4553 S.n3634 S.n3633 0.003
R4554 S.n3484 S.n3483 0.003
R4555 S.n3266 S.n3265 0.003
R4556 S.n2998 S.n2997 0.003
R4557 S.n2767 S.n2766 0.003
R4558 S.n2489 S.n2488 0.003
R4559 S.n2242 S.n2241 0.003
R4560 S.n1968 S.n1967 0.003
R4561 S.n1646 S.n1645 0.003
R4562 S.n1423 S.n1422 0.003
R4563 S.n1123 S.n1122 0.003
R4564 S.n914 S.n913 0.003
R4565 S.n464 S.n463 0.003
R4566 S.n1143 S.n1142 0.003
R4567 S.n1444 S.n1443 0.003
R4568 S.n1666 S.n1665 0.003
R4569 S.n1988 S.n1987 0.003
R4570 S.n2262 S.n2261 0.003
R4571 S.n2509 S.n2508 0.003
R4572 S.n2787 S.n2786 0.003
R4573 S.n3018 S.n3017 0.003
R4574 S.n3286 S.n3285 0.003
R4575 S.n3504 S.n3503 0.003
R4576 S.n3654 S.n3653 0.003
R4577 S.n3978 S.n3977 0.003
R4578 S.n4240 S.n4239 0.003
R4579 S.n4422 S.n4421 0.003
R4580 S.n4671 S.n4670 0.003
R4581 S.n4884 S.n4883 0.003
R4582 S.n593 S.n592 0.003
R4583 S.n818 S.n817 0.003
R4584 S.n425 S.n424 0.003
R4585 S.n408 S.n407 0.003
R4586 S.n233 S.n232 0.003
R4587 S.n731 S.n730 0.003
R4588 S.n2043 S.n2042 0.003
R4589 S.n1553 S.n1552 0.003
R4590 S.n1266 S.n1265 0.003
R4591 S.n1025 S.n1024 0.003
R4592 S.n256 S.n255 0.003
R4593 S.n2569 S.n2568 0.003
R4594 S.n2166 S.n2165 0.003
R4595 S.n1841 S.n1840 0.003
R4596 S.n1570 S.n1569 0.003
R4597 S.n1295 S.n1294 0.003
R4598 S.n1042 S.n1041 0.003
R4599 S.n760 S.n759 0.003
R4600 S.n392 S.n391 0.003
R4601 S.n375 S.n374 0.003
R4602 S.n181 S.n180 0.003
R4603 S.n960 S.n959 0.003
R4604 S.n212 S.n211 0.003
R4605 S.n1504 S.n1503 0.003
R4606 S.n1006 S.n1005 0.003
R4607 S.n701 S.n700 0.003
R4608 S.n359 S.n358 0.003
R4609 S.n342 S.n341 0.003
R4610 S.n647 S.n646 0.003
R4611 S.n496 S.n495 0.003
R4612 S.n1205 S.n1204 0.003
R4613 S.n1182 S.n1181 0.003
R4614 S.n1751 S.n1750 0.003
R4615 S.n1724 S.n1723 0.003
R4616 S.n2080 S.n2079 0.003
R4617 S.n2053 S.n2052 0.003
R4618 S.n2606 S.n2605 0.003
R4619 S.n2579 S.n2578 0.003
R4620 S.n3110 S.n3109 0.003
R4621 S.n3083 S.n3082 0.003
R4622 S.n3787 S.n3786 0.003
R4623 S.n3760 S.n3759 0.003
R4624 S.n4073 S.n4072 0.003
R4625 S.n4046 S.n4045 0.003
R4626 S.n4515 S.n4514 0.003
R4627 S.n4488 S.n4487 0.003
R4628 S.n4904 S.n4903 0.003
R4629 S.n5091 S.n5090 0.003
R4630 S.n5363 S.n5362 0.003
R4631 S.n1211 S.n1210 0.003
R4632 S.n1176 S.n1175 0.003
R4633 S.n1766 S.n1765 0.003
R4634 S.n5378 S.n5377 0.003
R4635 S.n5106 S.n5105 0.003
R4636 S.n4920 S.n4919 0.003
R4637 S.n4537 S.n4536 0.003
R4638 S.n4546 S.n4545 0.003
R4639 S.n4095 S.n4094 0.003
R4640 S.n4104 S.n4103 0.003
R4641 S.n3809 S.n3808 0.003
R4642 S.n3818 S.n3817 0.003
R4643 S.n3132 S.n3131 0.003
R4644 S.n3141 S.n3140 0.003
R4645 S.n2628 S.n2627 0.003
R4646 S.n2637 S.n2636 0.003
R4647 S.n2102 S.n2101 0.003
R4648 S.n2111 S.n2110 0.003
R4649 S.n1698 S.n1697 0.003
R4650 S.n1772 S.n1771 0.003
R4651 S.n1718 S.n1717 0.003
R4652 S.n2316 S.n2315 0.003
R4653 S.n5393 S.n5392 0.003
R4654 S.n5122 S.n5121 0.003
R4655 S.n4935 S.n4934 0.003
R4656 S.n4703 S.n4702 0.003
R4657 S.n4561 S.n4560 0.003
R4658 S.n4273 S.n4272 0.003
R4659 S.n4119 S.n4118 0.003
R4660 S.n3687 S.n3686 0.003
R4661 S.n3833 S.n3832 0.003
R4662 S.n3319 S.n3318 0.003
R4663 S.n3156 S.n3155 0.003
R4664 S.n2820 S.n2819 0.003
R4665 S.n2652 S.n2651 0.003
R4666 S.n2308 S.n2307 0.003
R4667 S.n2322 S.n2321 0.003
R4668 S.n2299 S.n2298 0.003
R4669 S.n2857 S.n2856 0.003
R4670 S.n5408 S.n5407 0.003
R4671 S.n5138 S.n5137 0.003
R4672 S.n4950 S.n4949 0.003
R4673 S.n4719 S.n4718 0.003
R4674 S.n4576 S.n4575 0.003
R4675 S.n4289 S.n4288 0.003
R4676 S.n4134 S.n4133 0.003
R4677 S.n3703 S.n3702 0.003
R4678 S.n3848 S.n3847 0.003
R4679 S.n3335 S.n3334 0.003
R4680 S.n3171 S.n3170 0.003
R4681 S.n2849 S.n2848 0.003
R4682 S.n2863 S.n2862 0.003
R4683 S.n2840 S.n2839 0.003
R4684 S.n3372 S.n3371 0.003
R4685 S.n5423 S.n5422 0.003
R4686 S.n5154 S.n5153 0.003
R4687 S.n4965 S.n4964 0.003
R4688 S.n4735 S.n4734 0.003
R4689 S.n4591 S.n4590 0.003
R4690 S.n4305 S.n4304 0.003
R4691 S.n4149 S.n4148 0.003
R4692 S.n3719 S.n3718 0.003
R4693 S.n3863 S.n3862 0.003
R4694 S.n3364 S.n3363 0.003
R4695 S.n3378 S.n3377 0.003
R4696 S.n3358 S.n3357 0.003
R4697 S.n3878 S.n3877 0.003
R4698 S.n5438 S.n5437 0.003
R4699 S.n5170 S.n5169 0.003
R4700 S.n4980 S.n4979 0.003
R4701 S.n4751 S.n4750 0.003
R4702 S.n4606 S.n4605 0.003
R4703 S.n4321 S.n4320 0.003
R4704 S.n4164 S.n4163 0.003
R4705 S.n3734 S.n3733 0.003
R4706 S.n3884 S.n3883 0.003
R4707 S.n3754 S.n3753 0.003
R4708 S.n4358 S.n4357 0.003
R4709 S.n5453 S.n5452 0.003
R4710 S.n5186 S.n5185 0.003
R4711 S.n4995 S.n4994 0.003
R4712 S.n4767 S.n4766 0.003
R4713 S.n4621 S.n4620 0.003
R4714 S.n4350 S.n4349 0.003
R4715 S.n4364 S.n4363 0.003
R4716 S.n4341 S.n4340 0.003
R4717 S.n4807 S.n4806 0.003
R4718 S.n5468 S.n5467 0.003
R4719 S.n5202 S.n5201 0.003
R4720 S.n5010 S.n5009 0.003
R4721 S.n4799 S.n4798 0.003
R4722 S.n4813 S.n4812 0.003
R4723 S.n4790 S.n4789 0.003
R4724 S.n5233 S.n5232 0.003
R4725 S.n5486 S.n5485 0.003
R4726 S.n5208 S.n5207 0.003
R4727 S.n5492 S.n5491 0.003
R4728 S.n1074 S.n1073 0.003
R4729 S.n5323 S.n5318 0.003
R4730 S.n5071 S.n5059 0.003
R4731 S.n638 S.n626 0.003
R4732 S.n608 S.n603 0.003
R4733 S.n933 S.n922 0.003
R4734 S.n5342 S.n5337 0.003
R4735 S.n5047 S.n5042 0.003
R4736 S.n4857 S.n4848 0.003
R4737 S.n4684 S.n4679 0.003
R4738 S.n4448 S.n4439 0.003
R4739 S.n4253 S.n4248 0.003
R4740 S.n4004 S.n3995 0.003
R4741 S.n3667 S.n3662 0.003
R4742 S.n3530 S.n3521 0.003
R4743 S.n3299 S.n3294 0.003
R4744 S.n3044 S.n3035 0.003
R4745 S.n2800 S.n2795 0.003
R4746 S.n2535 S.n2526 0.003
R4747 S.n2275 S.n2270 0.003
R4748 S.n2014 S.n2005 0.003
R4749 S.n1679 S.n1674 0.003
R4750 S.n1470 S.n1461 0.003
R4751 S.n1156 S.n1151 0.003
R4752 S.n475 S.n470 0.003
R4753 S.n271 S.n266 0.003
R4754 S.n784 S.n777 0.003
R4755 S.n3070 S.n3059 0.003
R4756 S.n2704 S.n2699 0.003
R4757 S.n2388 S.n2379 0.003
R4758 S.n2182 S.n2177 0.003
R4759 S.n1867 S.n1858 0.003
R4760 S.n1583 S.n1578 0.003
R4761 S.n1321 S.n1312 0.003
R4762 S.n1055 S.n1050 0.003
R4763 S.n294 S.n289 0.003
R4764 S.n3561 S.n3549 0.003
R4765 S.n3220 S.n3215 0.003
R4766 S.n2926 S.n2912 0.003
R4767 S.n2721 S.n2716 0.003
R4768 S.n2417 S.n2403 0.003
R4769 S.n2196 S.n2191 0.003
R4770 S.n1896 S.n1882 0.003
R4771 S.n1600 S.n1595 0.003
R4772 S.n1350 S.n1336 0.003
R4773 S.n1074 S.n1067 0.003
R4774 S.n1096 S.n1088 0.003
R4775 S.n846 S.n828 0.003
R4776 S.n510 S.n304 0.003
R4777 S.n525 S.n516 0.003
R4778 S.n1383 S.n1374 0.003
R4779 S.n1928 S.n1919 0.003
R4780 S.n2449 S.n2440 0.003
R4781 S.n2958 S.n2949 0.003
R4782 S.n3444 S.n3435 0.003
R4783 S.n4033 S.n4022 0.003
R4784 S.n3607 S.n3602 0.003
R4785 S.n3239 S.n3234 0.003
R4786 S.n2740 S.n2735 0.003
R4787 S.n2215 S.n2210 0.003
R4788 S.n1619 S.n1614 0.003
R4789 S.n880 S.n867 0.003
R4790 S.n439 S.n430 0.003
R4791 S.n558 S.n548 0.003
R4792 S.n4475 S.n4470 0.003
R4793 S.n4214 S.n4212 0.003
R4794 S.n3952 S.n3940 0.003
R4795 S.n3628 S.n3626 0.003
R4796 S.n3478 S.n3466 0.003
R4797 S.n3260 S.n3258 0.003
R4798 S.n2992 S.n2980 0.003
R4799 S.n2761 S.n2759 0.003
R4800 S.n2483 S.n2471 0.003
R4801 S.n2236 S.n2234 0.003
R4802 S.n1962 S.n1950 0.003
R4803 S.n1640 S.n1638 0.003
R4804 S.n1417 S.n1405 0.003
R4805 S.n1117 S.n1115 0.003
R4806 S.n908 S.n895 0.003
R4807 S.n458 S.n450 0.003
R4808 S.n1137 S.n1134 0.003
R4809 S.n1438 S.n1432 0.003
R4810 S.n1660 S.n1652 0.003
R4811 S.n1982 S.n1977 0.003
R4812 S.n2256 S.n2248 0.003
R4813 S.n2503 S.n2498 0.003
R4814 S.n2781 S.n2773 0.003
R4815 S.n3012 S.n3007 0.003
R4816 S.n3280 S.n3272 0.003
R4817 S.n3498 S.n3493 0.003
R4818 S.n3648 S.n3640 0.003
R4819 S.n3972 S.n3967 0.003
R4820 S.n4234 S.n4226 0.003
R4821 S.n4416 S.n4411 0.003
R4822 S.n4665 S.n4657 0.003
R4823 S.n4881 S.n4876 0.003
R4824 S.n587 S.n574 0.003
R4825 S.n812 S.n799 0.003
R4826 S.n419 S.n414 0.003
R4827 S.n402 S.n397 0.003
R4828 S.n227 S.n222 0.003
R4829 S.n725 S.n718 0.003
R4830 S.n2040 S.n2029 0.003
R4831 S.n1547 S.n1542 0.003
R4832 S.n1260 S.n1251 0.003
R4833 S.n1019 S.n1014 0.003
R4834 S.n250 S.n245 0.003
R4835 S.n2566 S.n2554 0.003
R4836 S.n2160 S.n2155 0.003
R4837 S.n1835 S.n1821 0.003
R4838 S.n1564 S.n1559 0.003
R4839 S.n1289 S.n1275 0.003
R4840 S.n1036 S.n1031 0.003
R4841 S.n754 S.n740 0.003
R4842 S.n386 S.n381 0.003
R4843 S.n369 S.n364 0.003
R4844 S.n186 S.n178 0.003
R4845 S.n957 S.n948 0.003
R4846 S.n206 S.n201 0.003
R4847 S.n1501 S.n1489 0.003
R4848 S.n1000 S.n995 0.003
R4849 S.n695 S.n681 0.003
R4850 S.n353 S.n348 0.003
R4851 S.n336 S.n331 0.003
R4852 S.n493 S.n487 0.003
R4853 S.n1202 S.n1196 0.003
R4854 S.n1192 S.n967 0.003
R4855 S.n1748 S.n1739 0.003
R4856 S.n1734 S.n1511 0.003
R4857 S.n2077 S.n2068 0.003
R4858 S.n2063 S.n2050 0.003
R4859 S.n2603 S.n2594 0.003
R4860 S.n2589 S.n2576 0.003
R4861 S.n3107 S.n3098 0.003
R4862 S.n3093 S.n3080 0.003
R4863 S.n3784 S.n3775 0.003
R4864 S.n3770 S.n3571 0.003
R4865 S.n4070 S.n4061 0.003
R4866 S.n4056 S.n4043 0.003
R4867 S.n4512 S.n4503 0.003
R4868 S.n4498 S.n4485 0.003
R4869 S.n4901 S.n4892 0.003
R4870 S.n5088 S.n5081 0.003
R4871 S.n5360 S.n5352 0.003
R4872 S.n1173 S.n1168 0.003
R4873 S.n1763 S.n1762 0.003
R4874 S.n5375 S.n5374 0.003
R4875 S.n5103 S.n5102 0.003
R4876 S.n4917 S.n4915 0.003
R4877 S.n4541 S.n4540 0.003
R4878 S.n4543 S.n4526 0.003
R4879 S.n4099 S.n4098 0.003
R4880 S.n4101 S.n4084 0.003
R4881 S.n3813 S.n3812 0.003
R4882 S.n3815 S.n3798 0.003
R4883 S.n3136 S.n3135 0.003
R4884 S.n3138 S.n3121 0.003
R4885 S.n2632 S.n2631 0.003
R4886 S.n2634 S.n2617 0.003
R4887 S.n2106 S.n2105 0.003
R4888 S.n2108 S.n2091 0.003
R4889 S.n1695 S.n1694 0.003
R4890 S.n1715 S.n1706 0.003
R4891 S.n2313 S.n2122 0.003
R4892 S.n5390 S.n5389 0.003
R4893 S.n5119 S.n5117 0.003
R4894 S.n4932 S.n4931 0.003
R4895 S.n4700 S.n4698 0.003
R4896 S.n4558 S.n4557 0.003
R4897 S.n4270 S.n4268 0.003
R4898 S.n4116 S.n4115 0.003
R4899 S.n3684 S.n3682 0.003
R4900 S.n3830 S.n3829 0.003
R4901 S.n3316 S.n3314 0.003
R4902 S.n3153 S.n3152 0.003
R4903 S.n2817 S.n2815 0.003
R4904 S.n2649 S.n2648 0.003
R4905 S.n2312 S.n2311 0.003
R4906 S.n2296 S.n2287 0.003
R4907 S.n2854 S.n2663 0.003
R4908 S.n5405 S.n5404 0.003
R4909 S.n5135 S.n5133 0.003
R4910 S.n4947 S.n4946 0.003
R4911 S.n4716 S.n4714 0.003
R4912 S.n4573 S.n4572 0.003
R4913 S.n4286 S.n4284 0.003
R4914 S.n4131 S.n4130 0.003
R4915 S.n3700 S.n3698 0.003
R4916 S.n3845 S.n3844 0.003
R4917 S.n3332 S.n3330 0.003
R4918 S.n3168 S.n3167 0.003
R4919 S.n2853 S.n2852 0.003
R4920 S.n2837 S.n2828 0.003
R4921 S.n3369 S.n3182 0.003
R4922 S.n5420 S.n5419 0.003
R4923 S.n5151 S.n5149 0.003
R4924 S.n4962 S.n4961 0.003
R4925 S.n4732 S.n4730 0.003
R4926 S.n4588 S.n4587 0.003
R4927 S.n4302 S.n4300 0.003
R4928 S.n4146 S.n4145 0.003
R4929 S.n3716 S.n3714 0.003
R4930 S.n3860 S.n3859 0.003
R4931 S.n3368 S.n3367 0.003
R4932 S.n3355 S.n3343 0.003
R4933 S.n3875 S.n3874 0.003
R4934 S.n5435 S.n5434 0.003
R4935 S.n5167 S.n5165 0.003
R4936 S.n4977 S.n4976 0.003
R4937 S.n4748 S.n4746 0.003
R4938 S.n4603 S.n4602 0.003
R4939 S.n4318 S.n4316 0.003
R4940 S.n4161 S.n4160 0.003
R4941 S.n3731 S.n3730 0.003
R4942 S.n3751 S.n3742 0.003
R4943 S.n4355 S.n4175 0.003
R4944 S.n5450 S.n5449 0.003
R4945 S.n5183 S.n5181 0.003
R4946 S.n4992 S.n4991 0.003
R4947 S.n4764 S.n4762 0.003
R4948 S.n4618 S.n4617 0.003
R4949 S.n4354 S.n4353 0.003
R4950 S.n4338 S.n4329 0.003
R4951 S.n4804 S.n4632 0.003
R4952 S.n5465 S.n5464 0.003
R4953 S.n5199 S.n5197 0.003
R4954 S.n5007 S.n5006 0.003
R4955 S.n4803 S.n4802 0.003
R4956 S.n4787 S.n4773 0.003
R4957 S.n5230 S.n5224 0.003
R4958 S.n5483 S.n5478 0.003
R4959 S.n5216 S.n5022 0.003
R4960 S.n668 S.n667 0.003
R4961 S.n2 S.n1 0.003
R4962 S.n10 S.n9 0.003
R4963 S.n18 S.n17 0.003
R4964 S.n32 S.n31 0.003
R4965 S.n4646 S.n4645 0.003
R4966 S.n635 S.n634 0.003
R4967 S.n523 S.n522 0.003
R4968 S.n4643 S.n4642 0.003
R4969 S.n3952 S.n3951 0.003
R4970 S.n3478 S.n3477 0.003
R4971 S.n2992 S.n2991 0.003
R4972 S.n2483 S.n2482 0.003
R4973 S.n1962 S.n1961 0.003
R4974 S.n1417 S.n1416 0.003
R4975 S.n880 S.n863 0.003
R4976 S.n5216 S.n5018 0.003
R4977 S.n3204 S.n3203 0.003
R4978 S.n2144 S.n2143 0.003
R4979 S.n984 S.n983 0.003
R4980 S.n4872 S.n4871 0.003
R4981 S.n3220 S.n3211 0.003
R4982 S.n2721 S.n2712 0.003
R4983 S.n2196 S.n2187 0.003
R4984 S.n1600 S.n1591 0.003
R4985 S.n1074 S.n1063 0.003
R4986 S.n2160 S.n2151 0.003
R4987 S.n1564 S.n1555 0.003
R4988 S.n1036 S.n1027 0.003
R4989 S.n1000 S.n991 0.003
R4990 S.n5323 S.n5314 0.003
R4991 S.n5498 S.n5497 0.003
R4992 S.n951 S.n950 0.003
R4993 S.n599 S.n598 0.003
R4994 S.n539 S.n538 0.003
R4995 S.n294 S.n286 0.002
R4996 S.n419 S.n411 0.002
R4997 S.n812 S.n791 0.002
R4998 S.n1074 S.n1064 0.002
R4999 S.n1350 S.n1333 0.002
R5000 S.n1600 S.n1592 0.002
R5001 S.n1896 S.n1879 0.002
R5002 S.n2196 S.n2188 0.002
R5003 S.n2417 S.n2400 0.002
R5004 S.n2721 S.n2713 0.002
R5005 S.n2926 S.n2909 0.002
R5006 S.n3220 S.n3212 0.002
R5007 S.n558 S.n545 0.002
R5008 S.n439 S.n427 0.002
R5009 S.n880 S.n864 0.002
R5010 S.n1117 S.n1103 0.002
R5011 S.n1417 S.n1390 0.002
R5012 S.n1640 S.n1626 0.002
R5013 S.n1962 S.n1935 0.002
R5014 S.n2236 S.n2222 0.002
R5015 S.n2483 S.n2456 0.002
R5016 S.n2761 S.n2747 0.002
R5017 S.n2992 S.n2965 0.002
R5018 S.n3260 S.n3246 0.002
R5019 S.n3478 S.n3451 0.002
R5020 S.n3628 S.n3614 0.002
R5021 S.n3952 S.n3925 0.002
R5022 S.n4214 S.n4200 0.002
R5023 S.n4665 S.n4654 0.002
R5024 S.n4416 S.n4408 0.002
R5025 S.n4234 S.n4223 0.002
R5026 S.n3972 S.n3964 0.002
R5027 S.n3648 S.n3637 0.002
R5028 S.n3498 S.n3490 0.002
R5029 S.n3280 S.n3269 0.002
R5030 S.n3012 S.n3004 0.002
R5031 S.n2781 S.n2770 0.002
R5032 S.n2503 S.n2495 0.002
R5033 S.n2256 S.n2245 0.002
R5034 S.n1982 S.n1974 0.002
R5035 S.n1660 S.n1649 0.002
R5036 S.n1438 S.n1429 0.002
R5037 S.n1137 S.n1124 0.002
R5038 S.n908 S.n892 0.002
R5039 S.n458 S.n447 0.002
R5040 S.n587 S.n565 0.002
R5041 S.n250 S.n242 0.002
R5042 S.n386 S.n378 0.002
R5043 S.n754 S.n732 0.002
R5044 S.n1036 S.n1028 0.002
R5045 S.n1289 S.n1272 0.002
R5046 S.n1564 S.n1556 0.002
R5047 S.n1835 S.n1818 0.002
R5048 S.n2160 S.n2152 0.002
R5049 S.n206 S.n198 0.002
R5050 S.n353 S.n345 0.002
R5051 S.n695 S.n673 0.002
R5052 S.n1000 S.n992 0.002
R5053 S.n5360 S.n5349 0.002
R5054 S.n5088 S.n5078 0.002
R5055 S.n4901 S.n4889 0.002
R5056 S.n4498 S.n4482 0.002
R5057 S.n4512 S.n4500 0.002
R5058 S.n4056 S.n4040 0.002
R5059 S.n4070 S.n4058 0.002
R5060 S.n3770 S.n3568 0.002
R5061 S.n3784 S.n3772 0.002
R5062 S.n3093 S.n3077 0.002
R5063 S.n3107 S.n3095 0.002
R5064 S.n2589 S.n2573 0.002
R5065 S.n2603 S.n2591 0.002
R5066 S.n2063 S.n2047 0.002
R5067 S.n2077 S.n2065 0.002
R5068 S.n1734 S.n1508 0.002
R5069 S.n1748 S.n1736 0.002
R5070 S.n1192 S.n964 0.002
R5071 S.n1202 S.n1193 0.002
R5072 S.n5375 S.n5367 0.002
R5073 S.n5103 S.n5095 0.002
R5074 S.n4917 S.n4908 0.002
R5075 S.n4541 S.n4527 0.002
R5076 S.n4543 S.n4519 0.002
R5077 S.n4099 S.n4085 0.002
R5078 S.n4101 S.n4077 0.002
R5079 S.n3813 S.n3799 0.002
R5080 S.n3815 S.n3791 0.002
R5081 S.n3136 S.n3122 0.002
R5082 S.n3138 S.n3114 0.002
R5083 S.n2632 S.n2618 0.002
R5084 S.n2634 S.n2610 0.002
R5085 S.n2106 S.n2092 0.002
R5086 S.n2108 S.n2084 0.002
R5087 S.n1695 S.n1687 0.002
R5088 S.n1763 S.n1755 0.002
R5089 S.n1173 S.n1165 0.002
R5090 S.n5390 S.n5382 0.002
R5091 S.n5119 S.n5110 0.002
R5092 S.n4932 S.n4924 0.002
R5093 S.n4700 S.n4691 0.002
R5094 S.n4558 S.n4550 0.002
R5095 S.n4270 S.n4261 0.002
R5096 S.n4116 S.n4108 0.002
R5097 S.n3684 S.n3675 0.002
R5098 S.n3830 S.n3822 0.002
R5099 S.n3316 S.n3307 0.002
R5100 S.n3153 S.n3145 0.002
R5101 S.n2817 S.n2808 0.002
R5102 S.n2649 S.n2641 0.002
R5103 S.n2312 S.n2123 0.002
R5104 S.n2313 S.n2115 0.002
R5105 S.n1715 S.n1703 0.002
R5106 S.n5405 S.n5397 0.002
R5107 S.n5135 S.n5126 0.002
R5108 S.n4947 S.n4939 0.002
R5109 S.n4716 S.n4707 0.002
R5110 S.n4573 S.n4565 0.002
R5111 S.n4286 S.n4277 0.002
R5112 S.n4131 S.n4123 0.002
R5113 S.n3700 S.n3691 0.002
R5114 S.n3845 S.n3837 0.002
R5115 S.n3332 S.n3323 0.002
R5116 S.n3168 S.n3160 0.002
R5117 S.n2853 S.n2664 0.002
R5118 S.n2854 S.n2656 0.002
R5119 S.n2296 S.n2284 0.002
R5120 S.n5420 S.n5412 0.002
R5121 S.n5151 S.n5142 0.002
R5122 S.n4962 S.n4954 0.002
R5123 S.n4732 S.n4723 0.002
R5124 S.n4588 S.n4580 0.002
R5125 S.n4302 S.n4293 0.002
R5126 S.n4146 S.n4138 0.002
R5127 S.n3716 S.n3707 0.002
R5128 S.n3860 S.n3852 0.002
R5129 S.n3368 S.n3183 0.002
R5130 S.n3369 S.n3175 0.002
R5131 S.n2837 S.n2825 0.002
R5132 S.n5435 S.n5427 0.002
R5133 S.n5167 S.n5158 0.002
R5134 S.n4977 S.n4969 0.002
R5135 S.n4748 S.n4739 0.002
R5136 S.n4603 S.n4595 0.002
R5137 S.n4318 S.n4309 0.002
R5138 S.n4161 S.n4153 0.002
R5139 S.n3731 S.n3723 0.002
R5140 S.n3875 S.n3867 0.002
R5141 S.n3355 S.n3340 0.002
R5142 S.n5450 S.n5442 0.002
R5143 S.n5183 S.n5174 0.002
R5144 S.n4992 S.n4984 0.002
R5145 S.n4764 S.n4755 0.002
R5146 S.n4618 S.n4610 0.002
R5147 S.n4354 S.n4176 0.002
R5148 S.n4355 S.n4168 0.002
R5149 S.n3751 S.n3739 0.002
R5150 S.n5465 S.n5457 0.002
R5151 S.n5199 S.n5190 0.002
R5152 S.n5007 S.n4999 0.002
R5153 S.n4803 S.n4633 0.002
R5154 S.n4804 S.n4625 0.002
R5155 S.n4338 S.n4326 0.002
R5156 S.n5216 S.n5019 0.002
R5157 S.n5483 S.n5475 0.002
R5158 S.n4787 S.n4777 0.002
R5159 S.n5230 S.n5221 0.002
R5160 S.n5071 S.n5056 0.002
R5161 S.n5323 S.n5315 0.002
R5162 S.n638 S.n623 0.002
R5163 S.n3561 S.n3546 0.002
R5164 S.n4475 S.n4456 0.002
R5165 S.n2566 S.n2551 0.002
R5166 S.n1501 S.n1486 0.002
R5167 S.n4881 S.n4873 0.002
R5168 S.n1806 S.n1805 0.002
R5169 S.n2356 S.n2355 0.002
R5170 S.n2897 S.n2896 0.002
R5171 S.n3412 S.n3411 0.002
R5172 S.n3918 S.n3917 0.002
R5173 S.n4396 S.n4395 0.002
R5174 S.t2 S.n128 0.002
R5175 S.n1202 S.n1201 0.002
R5176 S.n622 S.n621 0.002
R5177 S.n5341 S.n5340 0.002
R5178 S.n4027 S.n4026 0.002
R5179 S.n3064 S.n3063 0.002
R5180 S.n2034 S.n2033 0.002
R5181 S.n933 S.n916 0.002
R5182 S.n784 S.n771 0.002
R5183 S.n1350 S.n1349 0.002
R5184 S.n1600 S.n1599 0.002
R5185 S.n1896 S.n1895 0.002
R5186 S.n2196 S.n2195 0.002
R5187 S.n2417 S.n2416 0.002
R5188 S.n2721 S.n2720 0.002
R5189 S.n2926 S.n2925 0.002
R5190 S.n3220 S.n3219 0.002
R5191 S.n725 S.n712 0.002
R5192 S.n1036 S.n1035 0.002
R5193 S.n1289 S.n1288 0.002
R5194 S.n1564 S.n1563 0.002
R5195 S.n1835 S.n1834 0.002
R5196 S.n2160 S.n2159 0.002
R5197 S.n1000 S.n999 0.002
R5198 S.n1763 S.n1756 0.002
R5199 S.n2313 S.n2116 0.002
R5200 S.n2854 S.n2657 0.002
R5201 S.n3369 S.n3176 0.002
R5202 S.n3875 S.n3868 0.002
R5203 S.n4355 S.n4169 0.002
R5204 S.n4804 S.n4626 0.002
R5205 S.n5216 S.n5215 0.002
R5206 S.n5483 S.n5482 0.002
R5207 S.n5071 S.n5070 0.002
R5208 S.n5323 S.n5322 0.002
R5209 S.n3545 S.n3544 0.002
R5210 S.n2550 S.n2549 0.002
R5211 S.n1485 S.n1484 0.002
R5212 S.n48 S.n45 0.002
R5213 S.n5047 S.n5036 0.002
R5214 S.n4857 S.n4842 0.002
R5215 S.n4684 S.n4673 0.002
R5216 S.n4448 S.n4433 0.002
R5217 S.n4253 S.n4242 0.002
R5218 S.n4004 S.n3989 0.002
R5219 S.n3667 S.n3656 0.002
R5220 S.n3530 S.n3515 0.002
R5221 S.n3299 S.n3288 0.002
R5222 S.n3044 S.n3029 0.002
R5223 S.n2800 S.n2789 0.002
R5224 S.n2535 S.n2520 0.002
R5225 S.n2275 S.n2264 0.002
R5226 S.n2014 S.n1999 0.002
R5227 S.n1679 S.n1668 0.002
R5228 S.n1470 S.n1455 0.002
R5229 S.n1156 S.n1145 0.002
R5230 S.n475 S.n474 0.002
R5231 S.n2704 S.n2693 0.002
R5232 S.n2388 S.n2373 0.002
R5233 S.n2182 S.n2171 0.002
R5234 S.n1867 S.n1852 0.002
R5235 S.n1583 S.n1572 0.002
R5236 S.n1321 S.n1306 0.002
R5237 S.n1055 S.n1044 0.002
R5238 S.n812 S.n811 0.002
R5239 S.n419 S.n418 0.002
R5240 S.n402 S.n401 0.002
R5241 S.n1547 S.n1536 0.002
R5242 S.n1260 S.n1245 0.002
R5243 S.n1019 S.n1008 0.002
R5244 S.n754 S.n753 0.002
R5245 S.n386 S.n385 0.002
R5246 S.n369 S.n368 0.002
R5247 S.n695 S.n694 0.002
R5248 S.n353 S.n352 0.002
R5249 S.n336 S.n335 0.002
R5250 S.n5375 S.n5368 0.002
R5251 S.n5103 S.n5096 0.002
R5252 S.n4917 S.n4909 0.002
R5253 S.n4541 S.n4528 0.002
R5254 S.n4543 S.n4520 0.002
R5255 S.n4099 S.n4086 0.002
R5256 S.n4101 S.n4078 0.002
R5257 S.n3813 S.n3800 0.002
R5258 S.n3815 S.n3792 0.002
R5259 S.n3136 S.n3123 0.002
R5260 S.n3138 S.n3115 0.002
R5261 S.n2632 S.n2619 0.002
R5262 S.n2634 S.n2611 0.002
R5263 S.n2106 S.n2093 0.002
R5264 S.n2108 S.n2085 0.002
R5265 S.n1695 S.n1688 0.002
R5266 S.n1173 S.n1172 0.002
R5267 S.n5390 S.n5383 0.002
R5268 S.n5119 S.n5111 0.002
R5269 S.n4932 S.n4925 0.002
R5270 S.n4700 S.n4692 0.002
R5271 S.n4558 S.n4551 0.002
R5272 S.n4270 S.n4262 0.002
R5273 S.n4116 S.n4109 0.002
R5274 S.n3684 S.n3676 0.002
R5275 S.n3830 S.n3823 0.002
R5276 S.n3316 S.n3308 0.002
R5277 S.n3153 S.n3146 0.002
R5278 S.n2817 S.n2809 0.002
R5279 S.n2649 S.n2642 0.002
R5280 S.n2312 S.n2124 0.002
R5281 S.n1715 S.n1714 0.002
R5282 S.n5405 S.n5398 0.002
R5283 S.n5135 S.n5127 0.002
R5284 S.n4947 S.n4940 0.002
R5285 S.n4716 S.n4708 0.002
R5286 S.n4573 S.n4566 0.002
R5287 S.n4286 S.n4278 0.002
R5288 S.n4131 S.n4124 0.002
R5289 S.n3700 S.n3692 0.002
R5290 S.n3845 S.n3838 0.002
R5291 S.n3332 S.n3324 0.002
R5292 S.n3168 S.n3161 0.002
R5293 S.n2853 S.n2665 0.002
R5294 S.n2296 S.n2295 0.002
R5295 S.n5420 S.n5413 0.002
R5296 S.n5151 S.n5143 0.002
R5297 S.n4962 S.n4955 0.002
R5298 S.n4732 S.n4724 0.002
R5299 S.n4588 S.n4581 0.002
R5300 S.n4302 S.n4294 0.002
R5301 S.n4146 S.n4139 0.002
R5302 S.n3716 S.n3708 0.002
R5303 S.n3860 S.n3853 0.002
R5304 S.n3368 S.n3184 0.002
R5305 S.n2837 S.n2836 0.002
R5306 S.n5435 S.n5428 0.002
R5307 S.n5167 S.n5159 0.002
R5308 S.n4977 S.n4970 0.002
R5309 S.n4748 S.n4740 0.002
R5310 S.n4603 S.n4596 0.002
R5311 S.n4318 S.n4310 0.002
R5312 S.n4161 S.n4154 0.002
R5313 S.n3731 S.n3724 0.002
R5314 S.n3355 S.n3354 0.002
R5315 S.n5450 S.n5443 0.002
R5316 S.n5183 S.n5175 0.002
R5317 S.n4992 S.n4985 0.002
R5318 S.n4764 S.n4756 0.002
R5319 S.n4618 S.n4611 0.002
R5320 S.n4354 S.n4177 0.002
R5321 S.n3751 S.n3750 0.002
R5322 S.n5465 S.n5458 0.002
R5323 S.n5199 S.n5191 0.002
R5324 S.n5007 S.n5000 0.002
R5325 S.n4803 S.n4634 0.002
R5326 S.n4338 S.n4337 0.002
R5327 S.n5230 S.n5229 0.002
R5328 S.n558 S.n544 0.002
R5329 S.n587 S.n584 0.002
R5330 S.n4787 S.n4783 0.002
R5331 S.n5342 S.n5331 0.002
R5332 S.n3070 S.n3053 0.002
R5333 S.n2040 S.n2023 0.002
R5334 S.n957 S.n942 0.002
R5335 S.n52 S.n51 0.002
R5336 S.n4881 S.n4880 0.002
R5337 S.n4416 S.n4415 0.002
R5338 S.n3972 S.n3971 0.002
R5339 S.n3498 S.n3497 0.002
R5340 S.n3012 S.n3011 0.002
R5341 S.n2503 S.n2502 0.002
R5342 S.n1982 S.n1981 0.002
R5343 S.n1438 S.n1437 0.002
R5344 S.n1715 S.n1702 0.002
R5345 S.n2817 S.n2816 0.002
R5346 S.n3316 S.n3315 0.002
R5347 S.n3684 S.n3683 0.002
R5348 S.n4270 S.n4269 0.002
R5349 S.n4700 S.n4699 0.002
R5350 S.n5119 S.n5118 0.002
R5351 S.n2296 S.n2283 0.002
R5352 S.n3332 S.n3331 0.002
R5353 S.n3700 S.n3699 0.002
R5354 S.n4286 S.n4285 0.002
R5355 S.n4716 S.n4715 0.002
R5356 S.n5135 S.n5134 0.002
R5357 S.n2837 S.n2824 0.002
R5358 S.n3716 S.n3715 0.002
R5359 S.n4302 S.n4301 0.002
R5360 S.n4732 S.n4731 0.002
R5361 S.n5151 S.n5150 0.002
R5362 S.n3355 S.n3339 0.002
R5363 S.n4318 S.n4317 0.002
R5364 S.n4748 S.n4747 0.002
R5365 S.n5167 S.n5166 0.002
R5366 S.n3751 S.n3738 0.002
R5367 S.n4764 S.n4763 0.002
R5368 S.n5183 S.n5182 0.002
R5369 S.n4338 S.n4325 0.002
R5370 S.n5199 S.n5198 0.002
R5371 S.n4214 S.n4213 0.002
R5372 S.n3628 S.n3627 0.002
R5373 S.n3260 S.n3259 0.002
R5374 S.n2761 S.n2760 0.002
R5375 S.n2236 S.n2235 0.002
R5376 S.n1640 S.n1639 0.002
R5377 S.n1117 S.n1116 0.002
R5378 S.n439 S.n426 0.002
R5379 S.n493 S.n483 0.002
R5380 S.n1735 S.n1734 0.002
R5381 S.n2064 S.n2063 0.002
R5382 S.n2590 S.n2589 0.002
R5383 S.n3094 S.n3093 0.002
R5384 S.n3771 S.n3770 0.002
R5385 S.n4057 S.n4056 0.002
R5386 S.n4499 S.n4498 0.002
R5387 S.n1173 S.n1164 0.002
R5388 S.n2107 S.n2106 0.002
R5389 S.n2633 S.n2632 0.002
R5390 S.n3137 S.n3136 0.002
R5391 S.n3814 S.n3813 0.002
R5392 S.n4100 S.n4099 0.002
R5393 S.n4542 S.n4541 0.002
R5394 S.n5342 S.n5330 0.002
R5395 S.n5047 S.n5035 0.002
R5396 S.n4857 S.n4832 0.002
R5397 S.n4684 S.n4672 0.002
R5398 S.n4448 S.n4423 0.002
R5399 S.n4253 S.n4241 0.002
R5400 S.n4004 S.n3979 0.002
R5401 S.n3667 S.n3655 0.002
R5402 S.n3530 S.n3505 0.002
R5403 S.n3299 S.n3287 0.002
R5404 S.n3044 S.n3019 0.002
R5405 S.n2800 S.n2788 0.002
R5406 S.n2535 S.n2510 0.002
R5407 S.n2275 S.n2263 0.002
R5408 S.n2014 S.n1989 0.002
R5409 S.n1679 S.n1667 0.002
R5410 S.n1470 S.n1445 0.002
R5411 S.n1156 S.n1144 0.002
R5412 S.n933 S.n915 0.002
R5413 S.n475 S.n465 0.002
R5414 S.n608 S.n600 0.002
R5415 S.n4033 S.n4012 0.002
R5416 S.n3607 S.n3595 0.002
R5417 S.n3444 S.n3419 0.002
R5418 S.n3239 S.n3227 0.002
R5419 S.n2958 S.n2933 0.002
R5420 S.n2740 S.n2728 0.002
R5421 S.n2449 S.n2424 0.002
R5422 S.n2215 S.n2203 0.002
R5423 S.n1928 S.n1903 0.002
R5424 S.n1619 S.n1607 0.002
R5425 S.n1383 S.n1357 0.002
R5426 S.n1096 S.n1085 0.002
R5427 S.n846 S.n825 0.002
R5428 S.n525 S.n513 0.002
R5429 S.n510 S.n301 0.002
R5430 S.n3070 S.n3052 0.002
R5431 S.n2704 S.n2692 0.002
R5432 S.n2388 S.n2363 0.002
R5433 S.n2182 S.n2170 0.002
R5434 S.n1867 S.n1842 0.002
R5435 S.n1583 S.n1571 0.002
R5436 S.n1321 S.n1296 0.002
R5437 S.n1055 S.n1043 0.002
R5438 S.n784 S.n761 0.002
R5439 S.n402 S.n393 0.002
R5440 S.n271 S.n263 0.002
R5441 S.n2040 S.n2022 0.002
R5442 S.n1547 S.n1535 0.002
R5443 S.n1260 S.n1235 0.002
R5444 S.n1019 S.n1007 0.002
R5445 S.n725 S.n702 0.002
R5446 S.n369 S.n360 0.002
R5447 S.n227 S.n219 0.002
R5448 S.n957 S.n941 0.002
R5449 S.n336 S.n327 0.002
R5450 S.n186 S.n175 0.002
R5451 S.n571 S.n570 0.002
R5452 S.n824 S.n823 0.001
R5453 S.n779 S.n778 0.001
R5454 S.n720 S.n719 0.001
R5455 S.n53 S.n52 0.001
R5456 S.t2 S.n53 0.001
R5457 S.n4407 S.n4406 0.001
R5458 S.n3963 S.n3962 0.001
R5459 S.n3489 S.n3488 0.001
R5460 S.n3003 S.n3002 0.001
R5461 S.n2494 S.n2493 0.001
R5462 S.n1973 S.n1972 0.001
R5463 S.n1428 S.n1427 0.001
R5464 S.n891 S.n890 0.001
R5465 S.t2 S.n30 0.001
R5466 S.t2 S.n3 0.001
R5467 S.t2 S.n100 0.001
R5468 S.t2 S.n111 0.001
R5469 S.t2 S.n11 0.001
R5470 S.t2 S.n20 0.001
R5471 S.n4820 S.n4819 0.001
R5472 S.n1383 S.n1368 0.001
R5473 S.n3560 S.n3559 0.001
R5474 S.n2565 S.n2564 0.001
R5475 S.n1500 S.n1499 0.001
R5476 S.n5257 S.n5256 0.001
R5477 S.n930 S.n929 0.001
R5478 S.n1153 S.n1152 0.001
R5479 S.n1467 S.n1466 0.001
R5480 S.n1676 S.n1675 0.001
R5481 S.n2011 S.n2010 0.001
R5482 S.n2272 S.n2271 0.001
R5483 S.n2532 S.n2531 0.001
R5484 S.n2797 S.n2796 0.001
R5485 S.n3041 S.n3040 0.001
R5486 S.n3296 S.n3295 0.001
R5487 S.n3527 S.n3526 0.001
R5488 S.n3664 S.n3663 0.001
R5489 S.n4001 S.n4000 0.001
R5490 S.n4250 S.n4249 0.001
R5491 S.n4445 S.n4444 0.001
R5492 S.n4681 S.n4680 0.001
R5493 S.n4854 S.n4853 0.001
R5494 S.n5044 S.n5043 0.001
R5495 S.n467 S.n466 0.001
R5496 S.n1084 S.n1083 0.001
R5497 S.n1380 S.n1379 0.001
R5498 S.n1616 S.n1615 0.001
R5499 S.n1925 S.n1924 0.001
R5500 S.n2212 S.n2211 0.001
R5501 S.n2446 S.n2445 0.001
R5502 S.n2737 S.n2736 0.001
R5503 S.n2955 S.n2954 0.001
R5504 S.n3236 S.n3235 0.001
R5505 S.n3441 S.n3440 0.001
R5506 S.n3604 S.n3603 0.001
R5507 S.n1052 S.n1051 0.001
R5508 S.n1318 S.n1317 0.001
R5509 S.n1580 S.n1579 0.001
R5510 S.n1864 S.n1863 0.001
R5511 S.n2179 S.n2178 0.001
R5512 S.n2385 S.n2384 0.001
R5513 S.n2701 S.n2700 0.001
R5514 S.n1016 S.n1015 0.001
R5515 S.n1257 S.n1256 0.001
R5516 S.n1544 S.n1543 0.001
R5517 S.n2908 S.n2907 0.001
R5518 S.n2399 S.n2398 0.001
R5519 S.n1878 S.n1877 0.001
R5520 S.n1332 S.n1331 0.001
R5521 S.n796 S.n795 0.001
R5522 S.n1817 S.n1816 0.001
R5523 S.n1271 S.n1270 0.001
R5524 S.n737 S.n736 0.001
R5525 S.n678 S.n677 0.001
R5526 S.n493 S.n484 0.001
R5527 S.n317 S.n316 0.001
R5528 S.n979 S.n978 0.001
R5529 S.n1525 S.n1524 0.001
R5530 S.n2139 S.n2138 0.001
R5531 S.n2682 S.n2681 0.001
R5532 S.n3199 S.n3198 0.001
R5533 S.n3585 S.n3584 0.001
R5534 S.n4189 S.n4188 0.001
R5535 S.n49 S.n48 0.001
R5536 S.n3444 S.n3429 0.001
R5537 S.n2958 S.n2943 0.001
R5538 S.n2449 S.n2434 0.001
R5539 S.n1928 S.n1913 0.001
R5540 S.n156 S.t2 0.001
R5541 S.t2 S.n127 0.001
R5542 S.t2 S.n86 0.001
R5543 S.t2 S.n74 0.001
R5544 S.t2 S.n62 0.001
R5545 S.n5308 S.n5307 0.001
R5546 S.n3205 S.n3204 0.001
R5547 S.n4195 S.n4194 0.001
R5548 S.n4647 S.n4646 0.001
R5549 S.n5030 S.n5029 0.001
R5550 S.n3590 S.n3589 0.001
R5551 S.n2145 S.n2144 0.001
R5552 S.n2687 S.n2686 0.001
R5553 S.n985 S.n984 0.001
R5554 S.n1530 S.n1529 0.001
R5555 S.n322 S.n321 0.001
R5556 S.n48 S.n47 0.001
R5557 S.n4033 S.n4014 0.001
R5558 S.n5360 S.n5359 0.001
R5559 S.n5088 S.n5087 0.001
R5560 S.n4901 S.n4900 0.001
R5561 S.n4498 S.n4497 0.001
R5562 S.n4512 S.n4511 0.001
R5563 S.n4056 S.n4055 0.001
R5564 S.n4070 S.n4069 0.001
R5565 S.n3770 S.n3769 0.001
R5566 S.n3784 S.n3783 0.001
R5567 S.n3093 S.n3092 0.001
R5568 S.n3107 S.n3106 0.001
R5569 S.n2589 S.n2588 0.001
R5570 S.n2603 S.n2602 0.001
R5571 S.n2063 S.n2062 0.001
R5572 S.n2077 S.n2076 0.001
R5573 S.n1734 S.n1733 0.001
R5574 S.n1748 S.n1747 0.001
R5575 S.n1192 S.n1191 0.001
R5576 S.n315 S.n314 0.001
R5577 S.n977 S.n976 0.001
R5578 S.n1523 S.n1522 0.001
R5579 S.n2137 S.n2136 0.001
R5580 S.n2680 S.n2679 0.001
R5581 S.n3197 S.n3196 0.001
R5582 S.n3583 S.n3582 0.001
R5583 S.n4187 S.n4186 0.001
R5584 S.t12 S.n322 0.001
R5585 S.t95 S.n3205 0.001
R5586 S.t53 S.n3590 0.001
R5587 S.t66 S.n4195 0.001
R5588 S.t31 S.n4647 0.001
R5589 S.t44 S.n5030 0.001
R5590 S.t8 S.n2145 0.001
R5591 S.t168 S.n2687 0.001
R5592 S.t151 S.n985 0.001
R5593 S.t42 S.n1530 0.001
R5594 S.n5307 S.t0 0.001
R5595 S.n1230 S.n1229 0.001
R5596 S.n316 S.n315 0.001
R5597 S.n978 S.n977 0.001
R5598 S.n1524 S.n1523 0.001
R5599 S.n2138 S.n2137 0.001
R5600 S.n2681 S.n2680 0.001
R5601 S.n3198 S.n3197 0.001
R5602 S.n3584 S.n3583 0.001
R5603 S.n4188 S.n4187 0.001
R5604 S.n5055 S.n5054 0.001
R5605 S.n511 S.n510 0.001
R5606 S.n402 S.n394 0.001
R5607 S.n369 S.n361 0.001
R5608 S.n336 S.n328 0.001
R5609 S.n661 S.n660 0.001
R5610 S.n1220 S.n1219 0.001
R5611 S.n1783 S.n1782 0.001
R5612 S.n2333 S.n2332 0.001
R5613 S.n2874 S.n2873 0.001
R5614 S.n3389 S.n3388 0.001
R5615 S.n3895 S.n3894 0.001
R5616 S.n4373 S.n4372 0.001
R5617 S.n553 S.n552 0.001
R5618 S.n48 S.n41 0.001
R5619 S.n48 S.n44 0.001
R5620 S.n48 S.n43 0.001
R5621 S.n48 S.n42 0.001
R5622 S.n5318 S.n5317 0.001
R5623 S.n5059 S.n5058 0.001
R5624 S.n626 S.n625 0.001
R5625 S.n603 S.n602 0.001
R5626 S.n922 S.n921 0.001
R5627 S.n5337 S.n5336 0.001
R5628 S.n5042 S.n5041 0.001
R5629 S.n4848 S.n4847 0.001
R5630 S.n4679 S.n4678 0.001
R5631 S.n4439 S.n4438 0.001
R5632 S.n4248 S.n4247 0.001
R5633 S.n3995 S.n3994 0.001
R5634 S.n3662 S.n3661 0.001
R5635 S.n3521 S.n3520 0.001
R5636 S.n3294 S.n3293 0.001
R5637 S.n3035 S.n3034 0.001
R5638 S.n2795 S.n2794 0.001
R5639 S.n2526 S.n2525 0.001
R5640 S.n2270 S.n2269 0.001
R5641 S.n2005 S.n2004 0.001
R5642 S.n1674 S.n1673 0.001
R5643 S.n1461 S.n1460 0.001
R5644 S.n1151 S.n1150 0.001
R5645 S.n470 S.n469 0.001
R5646 S.n266 S.n265 0.001
R5647 S.n777 S.n776 0.001
R5648 S.n3059 S.n3058 0.001
R5649 S.n2699 S.n2698 0.001
R5650 S.n2379 S.n2378 0.001
R5651 S.n2177 S.n2176 0.001
R5652 S.n1858 S.n1857 0.001
R5653 S.n1578 S.n1577 0.001
R5654 S.n1312 S.n1311 0.001
R5655 S.n1050 S.n1049 0.001
R5656 S.n289 S.n288 0.001
R5657 S.n3549 S.n3548 0.001
R5658 S.n3215 S.n3214 0.001
R5659 S.n2912 S.n2911 0.001
R5660 S.n2716 S.n2715 0.001
R5661 S.n2403 S.n2402 0.001
R5662 S.n2191 S.n2190 0.001
R5663 S.n1882 S.n1881 0.001
R5664 S.n1595 S.n1594 0.001
R5665 S.n1336 S.n1335 0.001
R5666 S.n1067 S.n1066 0.001
R5667 S.n1088 S.n1087 0.001
R5668 S.n828 S.n827 0.001
R5669 S.n304 S.n303 0.001
R5670 S.n516 S.n515 0.001
R5671 S.n1374 S.n1373 0.001
R5672 S.n1919 S.n1918 0.001
R5673 S.n2440 S.n2439 0.001
R5674 S.n2949 S.n2948 0.001
R5675 S.n3435 S.n3434 0.001
R5676 S.n4022 S.n4021 0.001
R5677 S.n3602 S.n3601 0.001
R5678 S.n3234 S.n3233 0.001
R5679 S.n2735 S.n2734 0.001
R5680 S.n2210 S.n2209 0.001
R5681 S.n1614 S.n1613 0.001
R5682 S.n867 S.n866 0.001
R5683 S.n430 S.n429 0.001
R5684 S.n548 S.n547 0.001
R5685 S.n4470 S.n4469 0.001
R5686 S.n4212 S.n4211 0.001
R5687 S.n3940 S.n3939 0.001
R5688 S.n3626 S.n3625 0.001
R5689 S.n3466 S.n3465 0.001
R5690 S.n3258 S.n3257 0.001
R5691 S.n2980 S.n2979 0.001
R5692 S.n2759 S.n2758 0.001
R5693 S.n2471 S.n2470 0.001
R5694 S.n2234 S.n2233 0.001
R5695 S.n1950 S.n1949 0.001
R5696 S.n1638 S.n1637 0.001
R5697 S.n1405 S.n1404 0.001
R5698 S.n1115 S.n1114 0.001
R5699 S.n895 S.n894 0.001
R5700 S.n450 S.n449 0.001
R5701 S.n1134 S.n1133 0.001
R5702 S.n1432 S.n1431 0.001
R5703 S.n1652 S.n1651 0.001
R5704 S.n1977 S.n1976 0.001
R5705 S.n2248 S.n2247 0.001
R5706 S.n2498 S.n2497 0.001
R5707 S.n2773 S.n2772 0.001
R5708 S.n3007 S.n3006 0.001
R5709 S.n3272 S.n3271 0.001
R5710 S.n3493 S.n3492 0.001
R5711 S.n3640 S.n3639 0.001
R5712 S.n3967 S.n3966 0.001
R5713 S.n4226 S.n4225 0.001
R5714 S.n4411 S.n4410 0.001
R5715 S.n4657 S.n4656 0.001
R5716 S.n4876 S.n4875 0.001
R5717 S.n574 S.n573 0.001
R5718 S.n799 S.n798 0.001
R5719 S.n414 S.n413 0.001
R5720 S.n397 S.n396 0.001
R5721 S.n222 S.n221 0.001
R5722 S.n718 S.n717 0.001
R5723 S.n2029 S.n2028 0.001
R5724 S.n1542 S.n1541 0.001
R5725 S.n1251 S.n1250 0.001
R5726 S.n1014 S.n1013 0.001
R5727 S.n245 S.n244 0.001
R5728 S.n2554 S.n2553 0.001
R5729 S.n2155 S.n2154 0.001
R5730 S.n1821 S.n1820 0.001
R5731 S.n1559 S.n1558 0.001
R5732 S.n1275 S.n1274 0.001
R5733 S.n1031 S.n1030 0.001
R5734 S.n740 S.n739 0.001
R5735 S.n381 S.n380 0.001
R5736 S.n364 S.n363 0.001
R5737 S.n178 S.n177 0.001
R5738 S.n948 S.n947 0.001
R5739 S.n201 S.n200 0.001
R5740 S.n1489 S.n1488 0.001
R5741 S.n995 S.n994 0.001
R5742 S.n681 S.n680 0.001
R5743 S.n348 S.n347 0.001
R5744 S.n331 S.n330 0.001
R5745 S.n487 S.n486 0.001
R5746 S.n1196 S.n1195 0.001
R5747 S.n967 S.n966 0.001
R5748 S.n1739 S.n1738 0.001
R5749 S.n1511 S.n1510 0.001
R5750 S.n2068 S.n2067 0.001
R5751 S.n2050 S.n2049 0.001
R5752 S.n2594 S.n2593 0.001
R5753 S.n2576 S.n2575 0.001
R5754 S.n3098 S.n3097 0.001
R5755 S.n3080 S.n3079 0.001
R5756 S.n3775 S.n3774 0.001
R5757 S.n3571 S.n3570 0.001
R5758 S.n4061 S.n4060 0.001
R5759 S.n4043 S.n4042 0.001
R5760 S.n4503 S.n4502 0.001
R5761 S.n4485 S.n4484 0.001
R5762 S.n4892 S.n4891 0.001
R5763 S.n5081 S.n5080 0.001
R5764 S.n5352 S.n5351 0.001
R5765 S.n1168 S.n1167 0.001
R5766 S.n1762 S.n1761 0.001
R5767 S.n5374 S.n5373 0.001
R5768 S.n5102 S.n5101 0.001
R5769 S.n4915 S.n4914 0.001
R5770 S.n4540 S.n4539 0.001
R5771 S.n4526 S.n4525 0.001
R5772 S.n4098 S.n4097 0.001
R5773 S.n4084 S.n4083 0.001
R5774 S.n3812 S.n3811 0.001
R5775 S.n3798 S.n3797 0.001
R5776 S.n3135 S.n3134 0.001
R5777 S.n3121 S.n3120 0.001
R5778 S.n2631 S.n2630 0.001
R5779 S.n2617 S.n2616 0.001
R5780 S.n2105 S.n2104 0.001
R5781 S.n2091 S.n2090 0.001
R5782 S.n1694 S.n1693 0.001
R5783 S.n1706 S.n1705 0.001
R5784 S.n2122 S.n2121 0.001
R5785 S.n5389 S.n5388 0.001
R5786 S.n5117 S.n5116 0.001
R5787 S.n4931 S.n4930 0.001
R5788 S.n4698 S.n4697 0.001
R5789 S.n4557 S.n4556 0.001
R5790 S.n4268 S.n4267 0.001
R5791 S.n4115 S.n4114 0.001
R5792 S.n3682 S.n3681 0.001
R5793 S.n3829 S.n3828 0.001
R5794 S.n3314 S.n3313 0.001
R5795 S.n3152 S.n3151 0.001
R5796 S.n2815 S.n2814 0.001
R5797 S.n2648 S.n2647 0.001
R5798 S.n2311 S.n2310 0.001
R5799 S.n2287 S.n2286 0.001
R5800 S.n2663 S.n2662 0.001
R5801 S.n5404 S.n5403 0.001
R5802 S.n5133 S.n5132 0.001
R5803 S.n4946 S.n4945 0.001
R5804 S.n4714 S.n4713 0.001
R5805 S.n4572 S.n4571 0.001
R5806 S.n4284 S.n4283 0.001
R5807 S.n4130 S.n4129 0.001
R5808 S.n3698 S.n3697 0.001
R5809 S.n3844 S.n3843 0.001
R5810 S.n3330 S.n3329 0.001
R5811 S.n3167 S.n3166 0.001
R5812 S.n2852 S.n2851 0.001
R5813 S.n2828 S.n2827 0.001
R5814 S.n3182 S.n3181 0.001
R5815 S.n5419 S.n5418 0.001
R5816 S.n5149 S.n5148 0.001
R5817 S.n4961 S.n4960 0.001
R5818 S.n4730 S.n4729 0.001
R5819 S.n4587 S.n4586 0.001
R5820 S.n4300 S.n4299 0.001
R5821 S.n4145 S.n4144 0.001
R5822 S.n3714 S.n3713 0.001
R5823 S.n3859 S.n3858 0.001
R5824 S.n3367 S.n3366 0.001
R5825 S.n3343 S.n3342 0.001
R5826 S.n3874 S.n3873 0.001
R5827 S.n5434 S.n5433 0.001
R5828 S.n5165 S.n5164 0.001
R5829 S.n4976 S.n4975 0.001
R5830 S.n4746 S.n4745 0.001
R5831 S.n4602 S.n4601 0.001
R5832 S.n4316 S.n4315 0.001
R5833 S.n4160 S.n4159 0.001
R5834 S.n3730 S.n3729 0.001
R5835 S.n3742 S.n3741 0.001
R5836 S.n4175 S.n4174 0.001
R5837 S.n5449 S.n5448 0.001
R5838 S.n5181 S.n5180 0.001
R5839 S.n4991 S.n4990 0.001
R5840 S.n4762 S.n4761 0.001
R5841 S.n4617 S.n4616 0.001
R5842 S.n4353 S.n4352 0.001
R5843 S.n4329 S.n4328 0.001
R5844 S.n4632 S.n4631 0.001
R5845 S.n5464 S.n5463 0.001
R5846 S.n5197 S.n5196 0.001
R5847 S.n5006 S.n5005 0.001
R5848 S.n4802 S.n4801 0.001
R5849 S.n4773 S.n4772 0.001
R5850 S.n5224 S.n5223 0.001
R5851 S.n5478 S.n5477 0.001
R5852 S.n5022 S.n5021 0.001
R5853 S.n48 S.n46 0.001
R5854 S.n4191 S.n4190 0.001
R5855 S.n3587 S.n3586 0.001
R5856 S.n3201 S.n3200 0.001
R5857 S.n2684 S.n2683 0.001
R5858 S.n2141 S.n2140 0.001
R5859 S.n1527 S.n1526 0.001
R5860 S.n981 S.n980 0.001
R5861 S.n319 S.n318 0.001
R5862 S.t62 S.n5329 0.001
R5863 S.t62 S.n5326 0.001
R5864 S.n5326 S.n5323 0.001
R5865 S.t44 S.n5077 0.001
R5866 S.t44 S.n5074 0.001
R5867 S.n5074 S.n5071 0.001
R5868 S.n5239 S.t79 0.001
R5869 S.n5260 S.n5241 0.001
R5870 S.t48 S.n641 0.001
R5871 S.t48 S.n644 0.001
R5872 S.t48 S.n614 0.001
R5873 S.t48 S.n611 0.001
R5874 S.n611 S.n608 0.001
R5875 S.t25 S.n939 0.001
R5876 S.t25 S.n936 0.001
R5877 S.n936 S.n933 0.001
R5878 S.t62 S.n5345 0.001
R5879 S.t62 S.n5348 0.001
R5880 S.t44 S.n5053 0.001
R5881 S.t44 S.n5050 0.001
R5882 S.n5050 S.n5047 0.001
R5883 S.t79 S.n4863 0.001
R5884 S.t79 S.n4860 0.001
R5885 S.n4860 S.n4857 0.001
R5886 S.t31 S.n4690 0.001
R5887 S.t31 S.n4687 0.001
R5888 S.n4687 S.n4684 0.001
R5889 S.t50 S.n4454 0.001
R5890 S.t50 S.n4451 0.001
R5891 S.n4451 S.n4448 0.001
R5892 S.t66 S.n4259 0.001
R5893 S.t66 S.n4256 0.001
R5894 S.n4256 S.n4253 0.001
R5895 S.t23 S.n4010 0.001
R5896 S.t23 S.n4007 0.001
R5897 S.n4007 S.n4004 0.001
R5898 S.t53 S.n3673 0.001
R5899 S.t53 S.n3670 0.001
R5900 S.n3670 S.n3667 0.001
R5901 S.t129 S.n3536 0.001
R5902 S.t129 S.n3533 0.001
R5903 S.n3533 S.n3530 0.001
R5904 S.t95 S.n3305 0.001
R5905 S.t95 S.n3302 0.001
R5906 S.n3302 S.n3299 0.001
R5907 S.t14 S.n3050 0.001
R5908 S.t14 S.n3047 0.001
R5909 S.n3047 S.n3044 0.001
R5910 S.t168 S.n2806 0.001
R5911 S.t168 S.n2803 0.001
R5912 S.n2803 S.n2800 0.001
R5913 S.t154 S.n2541 0.001
R5914 S.t154 S.n2538 0.001
R5915 S.n2538 S.n2535 0.001
R5916 S.t8 S.n2281 0.001
R5917 S.t8 S.n2278 0.001
R5918 S.n2278 S.n2275 0.001
R5919 S.t164 S.n2020 0.001
R5920 S.t164 S.n2017 0.001
R5921 S.n2017 S.n2014 0.001
R5922 S.t42 S.n1685 0.001
R5923 S.t42 S.n1682 0.001
R5924 S.n1682 S.n1679 0.001
R5925 S.t55 S.n1476 0.001
R5926 S.t55 S.n1473 0.001
R5927 S.n1473 S.n1470 0.001
R5928 S.t151 S.n1162 0.001
R5929 S.t151 S.n1159 0.001
R5930 S.n1159 S.n1156 0.001
R5931 S.t12 S.n481 0.001
R5932 S.t12 S.n478 0.001
R5933 S.n478 S.n475 0.001
R5934 S.t48 S.n277 0.001
R5935 S.t48 S.n274 0.001
R5936 S.n274 S.n271 0.001
R5937 S.t25 S.n790 0.001
R5938 S.t25 S.n787 0.001
R5939 S.n787 S.n784 0.001
R5940 S.t14 S.n3073 0.001
R5941 S.t14 S.n3076 0.001
R5942 S.t168 S.n2710 0.001
R5943 S.t168 S.n2707 0.001
R5944 S.n2707 S.n2704 0.001
R5945 S.t154 S.n2394 0.001
R5946 S.t154 S.n2391 0.001
R5947 S.n2391 S.n2388 0.001
R5948 S.t8 S.n2185 0.001
R5949 S.t8 S.n2169 0.001
R5950 S.t164 S.n1873 0.001
R5951 S.t164 S.n1870 0.001
R5952 S.n1870 S.n1867 0.001
R5953 S.t42 S.n1589 0.001
R5954 S.t42 S.n1586 0.001
R5955 S.n1586 S.n1583 0.001
R5956 S.t55 S.n1327 0.001
R5957 S.t55 S.n1324 0.001
R5958 S.n1324 S.n1321 0.001
R5959 S.t151 S.n1061 0.001
R5960 S.t151 S.n1058 0.001
R5961 S.n1058 S.n1055 0.001
R5962 S.t48 S.n300 0.001
R5963 S.t48 S.n297 0.001
R5964 S.n297 S.n294 0.001
R5965 S.t129 S.n3564 0.001
R5966 S.t129 S.n3567 0.001
R5967 S.t95 S.n3226 0.001
R5968 S.t95 S.n3223 0.001
R5969 S.n3223 S.n3220 0.001
R5970 S.t14 S.n2932 0.001
R5971 S.t14 S.n2929 0.001
R5972 S.n2929 S.n2926 0.001
R5973 S.t168 S.n2727 0.001
R5974 S.t168 S.n2724 0.001
R5975 S.n2724 S.n2721 0.001
R5976 S.t154 S.n2423 0.001
R5977 S.t154 S.n2420 0.001
R5978 S.n2420 S.n2417 0.001
R5979 S.t8 S.n2202 0.001
R5980 S.t8 S.n2199 0.001
R5981 S.n2199 S.n2196 0.001
R5982 S.t164 S.n1902 0.001
R5983 S.t164 S.n1899 0.001
R5984 S.n1899 S.n1896 0.001
R5985 S.t42 S.n1606 0.001
R5986 S.t42 S.n1603 0.001
R5987 S.n1603 S.n1600 0.001
R5988 S.t55 S.n1356 0.001
R5989 S.t55 S.n1353 0.001
R5990 S.n1353 S.n1350 0.001
R5991 S.t151 S.n1080 0.001
R5992 S.t151 S.n1077 0.001
R5993 S.n1077 S.n1074 0.001
R5994 S.t151 S.n1102 0.001
R5995 S.t151 S.n1099 0.001
R5996 S.n1099 S.n1096 0.001
R5997 S.t25 S.n852 0.001
R5998 S.t25 S.n849 0.001
R5999 S.n849 S.n846 0.001
R6000 S.n502 S.t12 0.001
R6001 S.n510 S.n505 0.001
R6002 S.t48 S.n531 0.001
R6003 S.t48 S.n528 0.001
R6004 S.n528 S.n525 0.001
R6005 S.t55 S.n1389 0.001
R6006 S.t55 S.n1386 0.001
R6007 S.n1386 S.n1383 0.001
R6008 S.t164 S.n1934 0.001
R6009 S.t164 S.n1931 0.001
R6010 S.n1931 S.n1928 0.001
R6011 S.t154 S.n2455 0.001
R6012 S.t154 S.n2452 0.001
R6013 S.n2452 S.n2449 0.001
R6014 S.t14 S.n2964 0.001
R6015 S.t14 S.n2961 0.001
R6016 S.n2961 S.n2958 0.001
R6017 S.t129 S.n3450 0.001
R6018 S.t129 S.n3447 0.001
R6019 S.n3447 S.n3444 0.001
R6020 S.t23 S.n4036 0.001
R6021 S.t23 S.n4039 0.001
R6022 S.t53 S.n3613 0.001
R6023 S.t53 S.n3610 0.001
R6024 S.n3610 S.n3607 0.001
R6025 S.t95 S.n3245 0.001
R6026 S.t95 S.n3242 0.001
R6027 S.n3242 S.n3239 0.001
R6028 S.t168 S.n2746 0.001
R6029 S.t168 S.n2743 0.001
R6030 S.n2743 S.n2740 0.001
R6031 S.t8 S.n2221 0.001
R6032 S.t8 S.n2218 0.001
R6033 S.n2218 S.n2215 0.001
R6034 S.t42 S.n1625 0.001
R6035 S.t42 S.n1622 0.001
R6036 S.n1622 S.n1619 0.001
R6037 S.t25 S.n886 0.001
R6038 S.t25 S.n883 0.001
R6039 S.n883 S.n880 0.001
R6040 S.t12 S.n445 0.001
R6041 S.t12 S.n442 0.001
R6042 S.n442 S.n439 0.001
R6043 S.t48 S.n564 0.001
R6044 S.t48 S.n561 0.001
R6045 S.n561 S.n558 0.001
R6046 S.t50 S.n4478 0.001
R6047 S.t50 S.n4481 0.001
R6048 S.t66 S.n4220 0.001
R6049 S.t66 S.n4217 0.001
R6050 S.n4217 S.n4214 0.001
R6051 S.t23 S.n3958 0.001
R6052 S.t23 S.n3955 0.001
R6053 S.n3955 S.n3952 0.001
R6054 S.t53 S.n3634 0.001
R6055 S.t53 S.n3631 0.001
R6056 S.n3631 S.n3628 0.001
R6057 S.t129 S.n3484 0.001
R6058 S.t129 S.n3481 0.001
R6059 S.n3481 S.n3478 0.001
R6060 S.t95 S.n3266 0.001
R6061 S.t95 S.n3263 0.001
R6062 S.n3263 S.n3260 0.001
R6063 S.t14 S.n2998 0.001
R6064 S.t14 S.n2995 0.001
R6065 S.n2995 S.n2992 0.001
R6066 S.t168 S.n2767 0.001
R6067 S.t168 S.n2764 0.001
R6068 S.n2764 S.n2761 0.001
R6069 S.t154 S.n2489 0.001
R6070 S.t154 S.n2486 0.001
R6071 S.n2486 S.n2483 0.001
R6072 S.t8 S.n2242 0.001
R6073 S.t8 S.n2239 0.001
R6074 S.n2239 S.n2236 0.001
R6075 S.t164 S.n1968 0.001
R6076 S.t164 S.n1965 0.001
R6077 S.n1965 S.n1962 0.001
R6078 S.t42 S.n1646 0.001
R6079 S.t42 S.n1643 0.001
R6080 S.n1643 S.n1640 0.001
R6081 S.t55 S.n1423 0.001
R6082 S.t55 S.n1420 0.001
R6083 S.n1420 S.n1417 0.001
R6084 S.t151 S.n1123 0.001
R6085 S.t151 S.n1120 0.001
R6086 S.n1120 S.n1117 0.001
R6087 S.t25 S.n914 0.001
R6088 S.t25 S.n911 0.001
R6089 S.n911 S.n908 0.001
R6090 S.t12 S.n464 0.001
R6091 S.t12 S.n461 0.001
R6092 S.n461 S.n458 0.001
R6093 S.t151 S.n1143 0.001
R6094 S.t151 S.n1140 0.001
R6095 S.n1140 S.n1137 0.001
R6096 S.t55 S.n1444 0.001
R6097 S.t55 S.n1441 0.001
R6098 S.n1441 S.n1438 0.001
R6099 S.t42 S.n1666 0.001
R6100 S.t42 S.n1663 0.001
R6101 S.n1663 S.n1660 0.001
R6102 S.t164 S.n1988 0.001
R6103 S.t164 S.n1985 0.001
R6104 S.n1985 S.n1982 0.001
R6105 S.t8 S.n2262 0.001
R6106 S.t8 S.n2259 0.001
R6107 S.n2259 S.n2256 0.001
R6108 S.t154 S.n2509 0.001
R6109 S.t154 S.n2506 0.001
R6110 S.n2506 S.n2503 0.001
R6111 S.t168 S.n2787 0.001
R6112 S.t168 S.n2784 0.001
R6113 S.n2784 S.n2781 0.001
R6114 S.t14 S.n3018 0.001
R6115 S.t14 S.n3015 0.001
R6116 S.n3015 S.n3012 0.001
R6117 S.t95 S.n3286 0.001
R6118 S.t95 S.n3283 0.001
R6119 S.n3283 S.n3280 0.001
R6120 S.t129 S.n3504 0.001
R6121 S.t129 S.n3501 0.001
R6122 S.n3501 S.n3498 0.001
R6123 S.t53 S.n3654 0.001
R6124 S.t53 S.n3651 0.001
R6125 S.n3651 S.n3648 0.001
R6126 S.t23 S.n3978 0.001
R6127 S.t23 S.n3975 0.001
R6128 S.n3975 S.n3972 0.001
R6129 S.t66 S.n4240 0.001
R6130 S.t66 S.n4237 0.001
R6131 S.n4237 S.n4234 0.001
R6132 S.t50 S.n4422 0.001
R6133 S.t50 S.n4419 0.001
R6134 S.n4419 S.n4416 0.001
R6135 S.t31 S.n4671 0.001
R6136 S.t31 S.n4668 0.001
R6137 S.n4668 S.n4665 0.001
R6138 S.t79 S.n4884 0.001
R6139 S.t79 S.n4887 0.001
R6140 S.t48 S.n593 0.001
R6141 S.t48 S.n590 0.001
R6142 S.n590 S.n587 0.001
R6143 S.t25 S.n818 0.001
R6144 S.t25 S.n815 0.001
R6145 S.n815 S.n812 0.001
R6146 S.t12 S.n425 0.001
R6147 S.t12 S.n422 0.001
R6148 S.n422 S.n419 0.001
R6149 S.t12 S.n408 0.001
R6150 S.t12 S.n405 0.001
R6151 S.n405 S.n402 0.001
R6152 S.t48 S.n233 0.001
R6153 S.t48 S.n230 0.001
R6154 S.n230 S.n227 0.001
R6155 S.t25 S.n731 0.001
R6156 S.t25 S.n728 0.001
R6157 S.n728 S.n725 0.001
R6158 S.t164 S.n2043 0.001
R6159 S.t164 S.n2046 0.001
R6160 S.t42 S.n1553 0.001
R6161 S.t42 S.n1550 0.001
R6162 S.n1550 S.n1547 0.001
R6163 S.t55 S.n1266 0.001
R6164 S.t55 S.n1263 0.001
R6165 S.n1263 S.n1260 0.001
R6166 S.t151 S.n1025 0.001
R6167 S.t151 S.n1022 0.001
R6168 S.n1022 S.n1019 0.001
R6169 S.t48 S.n256 0.001
R6170 S.t48 S.n253 0.001
R6171 S.n253 S.n250 0.001
R6172 S.t154 S.n2569 0.001
R6173 S.t154 S.n2572 0.001
R6174 S.t8 S.n2166 0.001
R6175 S.t8 S.n2163 0.001
R6176 S.n2163 S.n2160 0.001
R6177 S.t164 S.n1841 0.001
R6178 S.t164 S.n1838 0.001
R6179 S.n1838 S.n1835 0.001
R6180 S.t42 S.n1570 0.001
R6181 S.t42 S.n1567 0.001
R6182 S.n1567 S.n1564 0.001
R6183 S.t55 S.n1295 0.001
R6184 S.t55 S.n1292 0.001
R6185 S.n1292 S.n1289 0.001
R6186 S.t151 S.n1042 0.001
R6187 S.t151 S.n1039 0.001
R6188 S.n1039 S.n1036 0.001
R6189 S.t25 S.n760 0.001
R6190 S.t25 S.n757 0.001
R6191 S.n757 S.n754 0.001
R6192 S.t12 S.n392 0.001
R6193 S.t12 S.n389 0.001
R6194 S.n389 S.n386 0.001
R6195 S.t12 S.n375 0.001
R6196 S.t12 S.n372 0.001
R6197 S.n372 S.n369 0.001
R6198 S.t48 S.n189 0.001
R6199 S.n189 S.n186 0.001
R6200 S.t25 S.n960 0.001
R6201 S.t25 S.n963 0.001
R6202 S.t48 S.n212 0.001
R6203 S.t48 S.n209 0.001
R6204 S.n209 S.n206 0.001
R6205 S.t55 S.n1504 0.001
R6206 S.t55 S.n1507 0.001
R6207 S.t151 S.n1006 0.001
R6208 S.t151 S.n1003 0.001
R6209 S.n1003 S.n1000 0.001
R6210 S.t25 S.n701 0.001
R6211 S.t25 S.n698 0.001
R6212 S.n698 S.n695 0.001
R6213 S.t12 S.n359 0.001
R6214 S.t12 S.n356 0.001
R6215 S.n356 S.n353 0.001
R6216 S.t12 S.n342 0.001
R6217 S.t12 S.n339 0.001
R6218 S.n339 S.n336 0.001
R6219 S.n647 S.t48 0.001
R6220 S.n668 S.n649 0.001
R6221 S.t12 S.n496 0.001
R6222 S.t12 S.n499 0.001
R6223 S.t25 S.n1205 0.001
R6224 S.t25 S.n1208 0.001
R6225 S.n1182 S.t151 0.001
R6226 S.n1192 S.n1185 0.001
R6227 S.t55 S.n1751 0.001
R6228 S.t55 S.n1754 0.001
R6229 S.n1724 S.t42 0.001
R6230 S.n1734 S.n1727 0.001
R6231 S.t164 S.n2080 0.001
R6232 S.t164 S.n2083 0.001
R6233 S.n2063 S.n2056 0.001
R6234 S.t154 S.n2606 0.001
R6235 S.t154 S.n2609 0.001
R6236 S.n2589 S.n2582 0.001
R6237 S.t14 S.n3110 0.001
R6238 S.t14 S.n3113 0.001
R6239 S.n3093 S.n3086 0.001
R6240 S.t129 S.n3787 0.001
R6241 S.t129 S.n3790 0.001
R6242 S.n3760 S.t53 0.001
R6243 S.n3770 S.n3763 0.001
R6244 S.t23 S.n4073 0.001
R6245 S.t23 S.n4076 0.001
R6246 S.n4056 S.n4049 0.001
R6247 S.t50 S.n4515 0.001
R6248 S.t50 S.n4518 0.001
R6249 S.n4498 S.n4491 0.001
R6250 S.t79 S.n4904 0.001
R6251 S.t79 S.n4907 0.001
R6252 S.t44 S.n5091 0.001
R6253 S.t44 S.n5094 0.001
R6254 S.t62 S.n5363 0.001
R6255 S.t62 S.n5366 0.001
R6256 S.n5359 S.n5358 0.001
R6257 S.n5087 S.n5086 0.001
R6258 S.n4900 S.n4899 0.001
R6259 S.n4497 S.n4496 0.001
R6260 S.n4511 S.n4510 0.001
R6261 S.n4055 S.n4054 0.001
R6262 S.n4069 S.n4068 0.001
R6263 S.n3769 S.n3768 0.001
R6264 S.n3783 S.n3782 0.001
R6265 S.n3092 S.n3091 0.001
R6266 S.n3106 S.n3105 0.001
R6267 S.n2588 S.n2587 0.001
R6268 S.n2602 S.n2601 0.001
R6269 S.n2062 S.n2061 0.001
R6270 S.n2076 S.n2075 0.001
R6271 S.n1733 S.n1732 0.001
R6272 S.n1747 S.n1746 0.001
R6273 S.n1191 S.n1190 0.001
R6274 S.n1211 S.t25 0.001
R6275 S.n1229 S.n1213 0.001
R6276 S.t151 S.n1176 0.001
R6277 S.t151 S.n1179 0.001
R6278 S.t55 S.n1766 0.001
R6279 S.t55 S.n1769 0.001
R6280 S.t62 S.n5378 0.001
R6281 S.t62 S.n5381 0.001
R6282 S.t44 S.n5106 0.001
R6283 S.t44 S.n5109 0.001
R6284 S.t79 S.n4920 0.001
R6285 S.t79 S.n4923 0.001
R6286 S.n4541 S.n4534 0.001
R6287 S.t50 S.n4546 0.001
R6288 S.t50 S.n4549 0.001
R6289 S.n4099 S.n4092 0.001
R6290 S.t23 S.n4104 0.001
R6291 S.t23 S.n4107 0.001
R6292 S.n3813 S.n3806 0.001
R6293 S.t129 S.n3818 0.001
R6294 S.t129 S.n3821 0.001
R6295 S.n3136 S.n3129 0.001
R6296 S.t14 S.n3141 0.001
R6297 S.t14 S.n3144 0.001
R6298 S.n2632 S.n2625 0.001
R6299 S.t154 S.n2637 0.001
R6300 S.t154 S.n2640 0.001
R6301 S.n2106 S.n2099 0.001
R6302 S.t164 S.n2111 0.001
R6303 S.t164 S.n2114 0.001
R6304 S.t42 S.n1698 0.001
R6305 S.t42 S.n1701 0.001
R6306 S.n1772 S.t55 0.001
R6307 S.n1808 S.n1774 0.001
R6308 S.t42 S.n1718 0.001
R6309 S.t42 S.n1721 0.001
R6310 S.t164 S.n2316 0.001
R6311 S.t164 S.n2319 0.001
R6312 S.t62 S.n5393 0.001
R6313 S.t62 S.n5396 0.001
R6314 S.t44 S.n5122 0.001
R6315 S.t44 S.n5125 0.001
R6316 S.t79 S.n4935 0.001
R6317 S.t79 S.n4938 0.001
R6318 S.t31 S.n4703 0.001
R6319 S.t31 S.n4706 0.001
R6320 S.t50 S.n4561 0.001
R6321 S.t50 S.n4564 0.001
R6322 S.t66 S.n4273 0.001
R6323 S.t66 S.n4276 0.001
R6324 S.t23 S.n4119 0.001
R6325 S.t23 S.n4122 0.001
R6326 S.t53 S.n3687 0.001
R6327 S.t53 S.n3690 0.001
R6328 S.t129 S.n3833 0.001
R6329 S.t129 S.n3836 0.001
R6330 S.t95 S.n3319 0.001
R6331 S.t95 S.n3322 0.001
R6332 S.t14 S.n3156 0.001
R6333 S.t14 S.n3159 0.001
R6334 S.t168 S.n2820 0.001
R6335 S.t168 S.n2823 0.001
R6336 S.t154 S.n2652 0.001
R6337 S.t154 S.n2655 0.001
R6338 S.n2305 S.t8 0.001
R6339 S.n2312 S.n2305 0.001
R6340 S.n2322 S.t164 0.001
R6341 S.n2358 S.n2324 0.001
R6342 S.t8 S.n2299 0.001
R6343 S.t8 S.n2302 0.001
R6344 S.t154 S.n2857 0.001
R6345 S.t154 S.n2860 0.001
R6346 S.t62 S.n5408 0.001
R6347 S.t62 S.n5411 0.001
R6348 S.t44 S.n5138 0.001
R6349 S.t44 S.n5141 0.001
R6350 S.t79 S.n4950 0.001
R6351 S.t79 S.n4953 0.001
R6352 S.t31 S.n4719 0.001
R6353 S.t31 S.n4722 0.001
R6354 S.t50 S.n4576 0.001
R6355 S.t50 S.n4579 0.001
R6356 S.t66 S.n4289 0.001
R6357 S.t66 S.n4292 0.001
R6358 S.t23 S.n4134 0.001
R6359 S.t23 S.n4137 0.001
R6360 S.t53 S.n3703 0.001
R6361 S.t53 S.n3706 0.001
R6362 S.t129 S.n3848 0.001
R6363 S.t129 S.n3851 0.001
R6364 S.t95 S.n3335 0.001
R6365 S.t95 S.n3338 0.001
R6366 S.t14 S.n3171 0.001
R6367 S.t14 S.n3174 0.001
R6368 S.n2846 S.t168 0.001
R6369 S.n2853 S.n2846 0.001
R6370 S.n2863 S.t154 0.001
R6371 S.n2899 S.n2865 0.001
R6372 S.t168 S.n2840 0.001
R6373 S.t168 S.n2843 0.001
R6374 S.t14 S.n3372 0.001
R6375 S.t14 S.n3375 0.001
R6376 S.t62 S.n5423 0.001
R6377 S.t62 S.n5426 0.001
R6378 S.t44 S.n5154 0.001
R6379 S.t44 S.n5157 0.001
R6380 S.t79 S.n4965 0.001
R6381 S.t79 S.n4968 0.001
R6382 S.t31 S.n4735 0.001
R6383 S.t31 S.n4738 0.001
R6384 S.t50 S.n4591 0.001
R6385 S.t50 S.n4594 0.001
R6386 S.t66 S.n4305 0.001
R6387 S.t66 S.n4308 0.001
R6388 S.t23 S.n4149 0.001
R6389 S.t23 S.n4152 0.001
R6390 S.t53 S.n3719 0.001
R6391 S.t53 S.n3722 0.001
R6392 S.t129 S.n3863 0.001
R6393 S.t129 S.n3866 0.001
R6394 S.n3361 S.t95 0.001
R6395 S.n3368 S.n3361 0.001
R6396 S.n3378 S.t14 0.001
R6397 S.n3414 S.n3380 0.001
R6398 S.t95 S.n3358 0.001
R6399 S.n3355 S.n3346 0.001
R6400 S.t129 S.n3878 0.001
R6401 S.t129 S.n3881 0.001
R6402 S.t62 S.n5438 0.001
R6403 S.t62 S.n5441 0.001
R6404 S.t44 S.n5170 0.001
R6405 S.t44 S.n5173 0.001
R6406 S.t79 S.n4980 0.001
R6407 S.t79 S.n4983 0.001
R6408 S.t31 S.n4751 0.001
R6409 S.t31 S.n4754 0.001
R6410 S.t50 S.n4606 0.001
R6411 S.t50 S.n4609 0.001
R6412 S.t66 S.n4321 0.001
R6413 S.t66 S.n4324 0.001
R6414 S.t23 S.n4164 0.001
R6415 S.t23 S.n4167 0.001
R6416 S.t53 S.n3734 0.001
R6417 S.t53 S.n3737 0.001
R6418 S.n3884 S.t129 0.001
R6419 S.n3920 S.n3886 0.001
R6420 S.t53 S.n3754 0.001
R6421 S.t53 S.n3757 0.001
R6422 S.t23 S.n4358 0.001
R6423 S.t23 S.n4361 0.001
R6424 S.t62 S.n5453 0.001
R6425 S.t62 S.n5456 0.001
R6426 S.t44 S.n5186 0.001
R6427 S.t44 S.n5189 0.001
R6428 S.t79 S.n4995 0.001
R6429 S.t79 S.n4998 0.001
R6430 S.t31 S.n4767 0.001
R6431 S.t31 S.n4770 0.001
R6432 S.t50 S.n4621 0.001
R6433 S.t50 S.n4624 0.001
R6434 S.n4347 S.t66 0.001
R6435 S.n4354 S.n4347 0.001
R6436 S.n4364 S.t23 0.001
R6437 S.n4398 S.n4366 0.001
R6438 S.t66 S.n4341 0.001
R6439 S.t66 S.n4344 0.001
R6440 S.t50 S.n4807 0.001
R6441 S.t50 S.n4810 0.001
R6442 S.t62 S.n5468 0.001
R6443 S.t62 S.n5471 0.001
R6444 S.t44 S.n5202 0.001
R6445 S.t44 S.n5205 0.001
R6446 S.t79 S.n5010 0.001
R6447 S.t79 S.n5013 0.001
R6448 S.n4796 S.t31 0.001
R6449 S.n4803 S.n4796 0.001
R6450 S.n4813 S.t50 0.001
R6451 S.n4831 S.n4815 0.001
R6452 S.t31 S.n4790 0.001
R6453 S.t31 S.n4793 0.001
R6454 S.t79 S.n5233 0.001
R6455 S.t79 S.n5236 0.001
R6456 S.t62 S.n5486 0.001
R6457 S.t62 S.n5489 0.001
R6458 S.n5208 S.t44 0.001
R6459 S.n5216 S.n5211 0.001
R6460 S.n5492 S.t62 0.001
R6461 S.n5498 S.n5494 0.001
R6462 S.n36 S.n35 0.001
R6463 S.n40 S.n39 0.001
R6464 S.n665 S.n664 0.001
R6465 S.n1224 S.n1223 0.001
R6466 S.n1787 S.n1786 0.001
R6467 S.n2337 S.n2336 0.001
R6468 S.n2878 S.n2877 0.001
R6469 S.n3393 S.n3392 0.001
R6470 S.n3899 S.n3898 0.001
R6471 S.n4377 S.n4376 0.001
R6472 S.n4825 S.n4824 0.001
R6473 S.n5260 S.n5239 0.001
R6474 S.n5345 S.n5342 0.001
R6475 S.n4884 S.n4881 0.001
R6476 S.n4478 S.n4475 0.001
R6477 S.n510 S.n502 0.001
R6478 S.n4036 S.n4033 0.001
R6479 S.n3564 S.n3561 0.001
R6480 S.n2185 S.n2182 0.001
R6481 S.n3073 S.n3070 0.001
R6482 S.n2569 S.n2566 0.001
R6483 S.n2043 S.n2040 0.001
R6484 S.n1504 S.n1501 0.001
R6485 S.n186 S.n181 0.001
R6486 S.n960 S.n957 0.001
R6487 S.n641 S.n638 0.001
R6488 S.n5498 S.n5492 0.001
R6489 S.n668 S.n647 0.001
R6490 S.n5363 S.n5360 0.001
R6491 S.n5091 S.n5088 0.001
R6492 S.n4904 S.n4901 0.001
R6493 S.n4498 S.n4488 0.001
R6494 S.n4515 S.n4512 0.001
R6495 S.n4056 S.n4046 0.001
R6496 S.n4073 S.n4070 0.001
R6497 S.n3770 S.n3760 0.001
R6498 S.n3787 S.n3784 0.001
R6499 S.n3093 S.n3083 0.001
R6500 S.n3110 S.n3107 0.001
R6501 S.n2589 S.n2579 0.001
R6502 S.n2606 S.n2603 0.001
R6503 S.n2063 S.n2053 0.001
R6504 S.n2080 S.n2077 0.001
R6505 S.n1734 S.n1724 0.001
R6506 S.n1751 S.n1748 0.001
R6507 S.n1192 S.n1182 0.001
R6508 S.n1205 S.n1202 0.001
R6509 S.n496 S.n493 0.001
R6510 S.n1229 S.n1211 0.001
R6511 S.n5378 S.n5375 0.001
R6512 S.n5106 S.n5103 0.001
R6513 S.n4920 S.n4917 0.001
R6514 S.n4541 S.n4537 0.001
R6515 S.n4546 S.n4543 0.001
R6516 S.n4099 S.n4095 0.001
R6517 S.n4104 S.n4101 0.001
R6518 S.n3813 S.n3809 0.001
R6519 S.n3818 S.n3815 0.001
R6520 S.n3136 S.n3132 0.001
R6521 S.n3141 S.n3138 0.001
R6522 S.n2632 S.n2628 0.001
R6523 S.n2637 S.n2634 0.001
R6524 S.n2106 S.n2102 0.001
R6525 S.n2111 S.n2108 0.001
R6526 S.n1698 S.n1695 0.001
R6527 S.n1766 S.n1763 0.001
R6528 S.n1176 S.n1173 0.001
R6529 S.n1808 S.n1772 0.001
R6530 S.n1718 S.n1715 0.001
R6531 S.n2316 S.n2313 0.001
R6532 S.n2312 S.n2308 0.001
R6533 S.n2652 S.n2649 0.001
R6534 S.n2820 S.n2817 0.001
R6535 S.n3156 S.n3153 0.001
R6536 S.n3319 S.n3316 0.001
R6537 S.n3833 S.n3830 0.001
R6538 S.n3687 S.n3684 0.001
R6539 S.n4119 S.n4116 0.001
R6540 S.n4273 S.n4270 0.001
R6541 S.n4561 S.n4558 0.001
R6542 S.n4703 S.n4700 0.001
R6543 S.n4935 S.n4932 0.001
R6544 S.n5122 S.n5119 0.001
R6545 S.n5393 S.n5390 0.001
R6546 S.n2358 S.n2322 0.001
R6547 S.n2299 S.n2296 0.001
R6548 S.n2857 S.n2854 0.001
R6549 S.n2853 S.n2849 0.001
R6550 S.n3171 S.n3168 0.001
R6551 S.n3335 S.n3332 0.001
R6552 S.n3848 S.n3845 0.001
R6553 S.n3703 S.n3700 0.001
R6554 S.n4134 S.n4131 0.001
R6555 S.n4289 S.n4286 0.001
R6556 S.n4576 S.n4573 0.001
R6557 S.n4719 S.n4716 0.001
R6558 S.n4950 S.n4947 0.001
R6559 S.n5138 S.n5135 0.001
R6560 S.n5408 S.n5405 0.001
R6561 S.n2899 S.n2863 0.001
R6562 S.n2840 S.n2837 0.001
R6563 S.n3372 S.n3369 0.001
R6564 S.n3368 S.n3364 0.001
R6565 S.n3863 S.n3860 0.001
R6566 S.n3719 S.n3716 0.001
R6567 S.n4149 S.n4146 0.001
R6568 S.n4305 S.n4302 0.001
R6569 S.n4591 S.n4588 0.001
R6570 S.n4735 S.n4732 0.001
R6571 S.n4965 S.n4962 0.001
R6572 S.n5154 S.n5151 0.001
R6573 S.n5423 S.n5420 0.001
R6574 S.n3414 S.n3378 0.001
R6575 S.n3358 S.n3355 0.001
R6576 S.n3878 S.n3875 0.001
R6577 S.n3734 S.n3731 0.001
R6578 S.n4164 S.n4161 0.001
R6579 S.n4321 S.n4318 0.001
R6580 S.n4606 S.n4603 0.001
R6581 S.n4751 S.n4748 0.001
R6582 S.n4980 S.n4977 0.001
R6583 S.n5170 S.n5167 0.001
R6584 S.n5438 S.n5435 0.001
R6585 S.n3920 S.n3884 0.001
R6586 S.n3754 S.n3751 0.001
R6587 S.n4358 S.n4355 0.001
R6588 S.n4354 S.n4350 0.001
R6589 S.n4621 S.n4618 0.001
R6590 S.n4767 S.n4764 0.001
R6591 S.n4995 S.n4992 0.001
R6592 S.n5186 S.n5183 0.001
R6593 S.n5453 S.n5450 0.001
R6594 S.n4398 S.n4364 0.001
R6595 S.n4341 S.n4338 0.001
R6596 S.n4807 S.n4804 0.001
R6597 S.n4803 S.n4799 0.001
R6598 S.n5010 S.n5007 0.001
R6599 S.n5202 S.n5199 0.001
R6600 S.n5468 S.n5465 0.001
R6601 S.n4831 S.n4813 0.001
R6602 S.n4790 S.n4787 0.001
R6603 S.n5233 S.n5230 0.001
R6604 S.n5216 S.n5208 0.001
R6605 S.n5486 S.n5483 0.001
C0 DNW S 2936.40fF
C1 DNW G 6.22fF
C2 DNW D 355.65fF
C3 S G 1404.82fF
C4 S D 2210.20fF
C5 G D 1015.90fF
C6 D VSUBS -45.13fF
C7 G VSUBS -129.60fF
C8 S VSUBS 184.25fF $ **FLOATING
C9 DNW VSUBS 6933.01fF $ **FLOATING
C10 S.n0 VSUBS 0.95fF $ **FLOATING
C11 S.n1 VSUBS 0.34fF $ **FLOATING
C12 S.n2 VSUBS 0.33fF $ **FLOATING
C13 S.n3 VSUBS 2.61fF $ **FLOATING
C14 S.n4 VSUBS 8.88fF $ **FLOATING
C15 S.n5 VSUBS 8.88fF $ **FLOATING
C16 S.n6 VSUBS 5.33fF $ **FLOATING
C17 S.n7 VSUBS 2.15fF $ **FLOATING
C18 S.n8 VSUBS 0.95fF $ **FLOATING
C19 S.n9 VSUBS 0.34fF $ **FLOATING
C20 S.n10 VSUBS 0.33fF $ **FLOATING
C21 S.n11 VSUBS 2.61fF $ **FLOATING
C22 S.n12 VSUBS 8.88fF $ **FLOATING
C23 S.n13 VSUBS 8.88fF $ **FLOATING
C24 S.n14 VSUBS 5.33fF $ **FLOATING
C25 S.n15 VSUBS 2.15fF $ **FLOATING
C26 S.n16 VSUBS 0.95fF $ **FLOATING
C27 S.n17 VSUBS 0.34fF $ **FLOATING
C28 S.n18 VSUBS 0.33fF $ **FLOATING
C29 S.n19 VSUBS 9.27fF $ **FLOATING
C30 S.n20 VSUBS 2.61fF $ **FLOATING
C31 S.n21 VSUBS 8.88fF $ **FLOATING
C32 S.n22 VSUBS 8.88fF $ **FLOATING
C33 S.n23 VSUBS 5.33fF $ **FLOATING
C34 S.n24 VSUBS 2.15fF $ **FLOATING
C35 S.n25 VSUBS 13.46fF $ **FLOATING
C36 S.n26 VSUBS 13.46fF $ **FLOATING
C37 S.n27 VSUBS 5.28fF $ **FLOATING
C38 S.n28 VSUBS 2.02fF $ **FLOATING
C39 S.n29 VSUBS 16.23fF $ **FLOATING
C40 S.n30 VSUBS 2.61fF $ **FLOATING
C41 S.n31 VSUBS 0.34fF $ **FLOATING
C42 S.n32 VSUBS 0.30fF $ **FLOATING
C43 S.n33 VSUBS 0.95fF $ **FLOATING
C44 S.t892 VSUBS 0.02fF
C45 S.n34 VSUBS 1.29fF $ **FLOATING
C46 S.n35 VSUBS 38.81fF $ **FLOATING
C47 S.n36 VSUBS 2.20fF $ **FLOATING
C48 S.n37 VSUBS 0.35fF $ **FLOATING
C49 S.n38 VSUBS 0.62fF $ **FLOATING
C50 S.n39 VSUBS 0.52fF $ **FLOATING
C51 S.n40 VSUBS 3.63fF $ **FLOATING
C52 S.n41 VSUBS 4.20fF $ **FLOATING
C53 S.n42 VSUBS 4.17fF $ **FLOATING
C54 S.n43 VSUBS 4.17fF $ **FLOATING
C55 S.n44 VSUBS 4.17fF $ **FLOATING
C56 S.n45 VSUBS 4.64fF $ **FLOATING
C57 S.n46 VSUBS 4.25fF $ **FLOATING
C58 S.n47 VSUBS 4.23fF $ **FLOATING
C59 S.n48 VSUBS 85.89fF $ **FLOATING
C60 S.n49 VSUBS 2.17fF $ **FLOATING
C61 S.n50 VSUBS 12.76fF $ **FLOATING
C62 S.n51 VSUBS 1.87fF $ **FLOATING
C63 S.n52 VSUBS 9.30fF $ **FLOATING
C64 S.n53 VSUBS 0.25fF $ **FLOATING
C65 S.t540 VSUBS 0.02fF
C66 S.n54 VSUBS 0.44fF $ **FLOATING
C67 S.n55 VSUBS 8.88fF $ **FLOATING
C68 S.n56 VSUBS 8.88fF $ **FLOATING
C69 S.n57 VSUBS 5.40fF $ **FLOATING
C70 S.n58 VSUBS 1.94fF $ **FLOATING
C71 S.t768 VSUBS 0.02fF
C72 S.n59 VSUBS 0.88fF $ **FLOATING
C73 S.t555 VSUBS 0.02fF
C74 S.n60 VSUBS 0.88fF $ **FLOATING
C75 S.n61 VSUBS 9.33fF $ **FLOATING
C76 S.n62 VSUBS 3.25fF $ **FLOATING
C77 S.n63 VSUBS 0.38fF $ **FLOATING
C78 S.n64 VSUBS 0.30fF $ **FLOATING
C79 S.n65 VSUBS 0.99fF $ **FLOATING
C80 S.n66 VSUBS 0.02fF $ **FLOATING
C81 S.t1124 VSUBS 0.02fF
C82 S.n67 VSUBS 0.37fF $ **FLOATING
C83 S.n68 VSUBS 8.88fF $ **FLOATING
C84 S.n69 VSUBS 8.88fF $ **FLOATING
C85 S.n70 VSUBS 5.40fF $ **FLOATING
C86 S.n71 VSUBS 1.94fF $ **FLOATING
C87 S.t341 VSUBS 0.02fF
C88 S.n72 VSUBS 0.88fF $ **FLOATING
C89 S.t725 VSUBS 0.02fF
C90 S.n73 VSUBS 0.88fF $ **FLOATING
C91 S.n74 VSUBS 3.25fF $ **FLOATING
C92 S.n75 VSUBS 0.38fF $ **FLOATING
C93 S.n76 VSUBS 0.30fF $ **FLOATING
C94 S.n77 VSUBS 0.99fF $ **FLOATING
C95 S.n78 VSUBS 0.02fF $ **FLOATING
C96 S.t695 VSUBS 0.02fF
C97 S.n79 VSUBS 0.37fF $ **FLOATING
C98 S.n80 VSUBS 8.88fF $ **FLOATING
C99 S.n81 VSUBS 8.88fF $ **FLOATING
C100 S.n82 VSUBS 5.40fF $ **FLOATING
C101 S.n83 VSUBS 1.94fF $ **FLOATING
C102 S.t1086 VSUBS 0.02fF
C103 S.n84 VSUBS 0.88fF $ **FLOATING
C104 S.t304 VSUBS 0.02fF
C105 S.n85 VSUBS 0.88fF $ **FLOATING
C106 S.n86 VSUBS 3.25fF $ **FLOATING
C107 S.n87 VSUBS 0.38fF $ **FLOATING
C108 S.n88 VSUBS 0.30fF $ **FLOATING
C109 S.n89 VSUBS 0.99fF $ **FLOATING
C110 S.n90 VSUBS 0.02fF $ **FLOATING
C111 S.t279 VSUBS 0.02fF
C112 S.n91 VSUBS 0.37fF $ **FLOATING
C113 S.n92 VSUBS 0.30fF $ **FLOATING
C114 S.n93 VSUBS 8.88fF $ **FLOATING
C115 S.n94 VSUBS 8.88fF $ **FLOATING
C116 S.n95 VSUBS 5.16fF $ **FLOATING
C117 S.n96 VSUBS 0.99fF $ **FLOATING
C118 S.n97 VSUBS 0.35fF $ **FLOATING
C119 S.t78 VSUBS 0.02fF
C120 S.n98 VSUBS 0.88fF $ **FLOATING
C121 S.t478 VSUBS 0.02fF
C122 S.n99 VSUBS 0.88fF $ **FLOATING
C123 S.n100 VSUBS 3.35fF $ **FLOATING
C124 S.n101 VSUBS 0.27fF $ **FLOATING
C125 S.n102 VSUBS 1.04fF $ **FLOATING
C126 S.n103 VSUBS 1.13fF $ **FLOATING
C127 S.n104 VSUBS 0.42fF $ **FLOATING
C128 S.n105 VSUBS 0.02fF $ **FLOATING
C129 S.t1105 VSUBS 0.02fF
C130 S.n106 VSUBS 0.37fF $ **FLOATING
C131 S.n107 VSUBS 0.37fF $ **FLOATING
C132 S.n108 VSUBS 0.82fF $ **FLOATING
C133 S.t442 VSUBS 0.02fF
C134 S.n109 VSUBS 0.88fF $ **FLOATING
C135 S.t818 VSUBS 0.02fF
C136 S.n110 VSUBS 0.88fF $ **FLOATING
C137 S.n111 VSUBS 2.61fF $ **FLOATING
C138 S.n112 VSUBS 8.88fF $ **FLOATING
C139 S.n113 VSUBS 8.88fF $ **FLOATING
C140 S.n114 VSUBS 5.69fF $ **FLOATING
C141 S.n115 VSUBS 1.75fF $ **FLOATING
C142 S.n116 VSUBS 1.12fF $ **FLOATING
C143 S.n117 VSUBS 0.00fF $ **FLOATING
C144 S.n118 VSUBS 0.39fF $ **FLOATING
C145 S.n119 VSUBS 0.02fF $ **FLOATING
C146 S.t335 VSUBS 0.02fF
C147 S.n120 VSUBS 0.37fF $ **FLOATING
C148 S.n121 VSUBS 8.88fF $ **FLOATING
C149 S.n122 VSUBS 8.88fF $ **FLOATING
C150 S.n123 VSUBS 5.47fF $ **FLOATING
C151 S.n124 VSUBS 1.60fF $ **FLOATING
C152 S.t781 VSUBS 0.02fF
C153 S.n125 VSUBS 0.88fF $ **FLOATING
C154 S.t30 VSUBS 0.02fF
C155 S.n126 VSUBS 0.88fF $ **FLOATING
C156 S.n127 VSUBS 2.61fF $ **FLOATING
C157 S.n128 VSUBS 1.50fF $ **FLOATING
C158 S.n129 VSUBS 0.02fF $ **FLOATING
C159 S.t681 VSUBS 0.02fF
C160 S.n130 VSUBS 0.37fF $ **FLOATING
C161 S.n131 VSUBS 20.57fF $ **FLOATING
C162 S.n132 VSUBS 20.57fF $ **FLOATING
C163 S.n133 VSUBS 5.72fF $ **FLOATING
C164 S.n134 VSUBS 1.94fF $ **FLOATING
C165 S.t237 VSUBS 0.02fF
C166 S.n135 VSUBS 0.88fF $ **FLOATING
C167 S.t402 VSUBS 0.02fF
C168 S.n136 VSUBS 0.88fF $ **FLOATING
C169 S.n137 VSUBS 1.61fF $ **FLOATING
C170 S.n138 VSUBS 0.02fF $ **FLOATING
C171 S.t942 VSUBS 0.02fF
C172 S.n139 VSUBS 0.37fF $ **FLOATING
C173 S.t150 VSUBS 0.02fF
C174 S.n140 VSUBS 0.88fF $ **FLOATING
C175 S.n141 VSUBS 0.02fF $ **FLOATING
C176 S.t123 VSUBS 0.02fF
C177 S.n142 VSUBS 0.37fF $ **FLOATING
C178 S.t934 VSUBS 0.02fF
C179 S.n143 VSUBS 0.88fF $ **FLOATING
C180 S.t388 VSUBS 0.02fF
C181 S.n144 VSUBS 0.88fF $ **FLOATING
C182 S.n145 VSUBS 0.02fF $ **FLOATING
C183 S.t359 VSUBS 0.02fF
C184 S.n146 VSUBS 0.37fF $ **FLOATING
C185 S.t1110 VSUBS 0.02fF
C186 S.n147 VSUBS 0.88fF $ **FLOATING
C187 S.t1063 VSUBS 0.02fF
C188 S.n148 VSUBS 0.88fF $ **FLOATING
C189 S.n149 VSUBS 0.02fF $ **FLOATING
C190 S.t1036 VSUBS 0.02fF
C191 S.n150 VSUBS 0.37fF $ **FLOATING
C192 S.t684 VSUBS 0.02fF
C193 S.n151 VSUBS 0.88fF $ **FLOATING
C194 S.t119 VSUBS 0.02fF
C195 S.n152 VSUBS 0.88fF $ **FLOATING
C196 S.n153 VSUBS 0.02fF $ **FLOATING
C197 S.t765 VSUBS 0.02fF
C198 S.n154 VSUBS 0.37fF $ **FLOATING
C199 S.t857 VSUBS 0.02fF
C200 S.n155 VSUBS 0.88fF $ **FLOATING
C201 S.t2 VSUBS 114.16fF
C202 S.n156 VSUBS 3.25fF $ **FLOATING
C203 S.n157 VSUBS 9.33fF $ **FLOATING
C204 S.n158 VSUBS 9.27fF $ **FLOATING
C205 S.n159 VSUBS 9.33fF $ **FLOATING
C206 S.n160 VSUBS 9.27fF $ **FLOATING
C207 S.n161 VSUBS 9.27fF $ **FLOATING
C208 S.n162 VSUBS 9.27fF $ **FLOATING
C209 S.n163 VSUBS 9.33fF $ **FLOATING
C210 S.n164 VSUBS 11.41fF $ **FLOATING
C211 S.n165 VSUBS 1.17fF $ **FLOATING
C212 S.n166 VSUBS 0.38fF $ **FLOATING
C213 S.n167 VSUBS 1.19fF $ **FLOATING
C214 S.n168 VSUBS 0.36fF $ **FLOATING
C215 S.n169 VSUBS 0.64fF $ **FLOATING
C216 S.n170 VSUBS 0.43fF $ **FLOATING
C217 S.n171 VSUBS 1.60fF $ **FLOATING
C218 S.n172 VSUBS 0.49fF $ **FLOATING
C219 S.n173 VSUBS 0.45fF $ **FLOATING
C220 S.n174 VSUBS 0.45fF $ **FLOATING
C221 S.n175 VSUBS 1.82fF $ **FLOATING
C222 S.n176 VSUBS 0.12fF $ **FLOATING
C223 S.t436 VSUBS 0.02fF
C224 S.n177 VSUBS 0.14fF $ **FLOATING
C225 S.t814 VSUBS 0.02fF
C226 S.n179 VSUBS 0.12fF $ **FLOATING
C227 S.n180 VSUBS 0.14fF $ **FLOATING
C228 S.t791 VSUBS 0.02fF
C229 S.n182 VSUBS 0.24fF $ **FLOATING
C230 S.n183 VSUBS 0.35fF $ **FLOATING
C231 S.n184 VSUBS 0.60fF $ **FLOATING
C232 S.n185 VSUBS 2.46fF $ **FLOATING
C233 S.n186 VSUBS 2.00fF $ **FLOATING
C234 S.t912 VSUBS 0.02fF
C235 S.n187 VSUBS 0.24fF $ **FLOATING
C236 S.n188 VSUBS 0.90fF $ **FLOATING
C237 S.n189 VSUBS 0.05fF $ **FLOATING
C238 S.n190 VSUBS 0.18fF $ **FLOATING
C239 S.n191 VSUBS 0.09fF $ **FLOATING
C240 S.n192 VSUBS 0.93fF $ **FLOATING
C241 S.n193 VSUBS 0.46fF $ **FLOATING
C242 S.n194 VSUBS 0.76fF $ **FLOATING
C243 S.n195 VSUBS 0.21fF $ **FLOATING
C244 S.n196 VSUBS 0.35fF $ **FLOATING
C245 S.n197 VSUBS 0.53fF $ **FLOATING
C246 S.n198 VSUBS 1.60fF $ **FLOATING
C247 S.n199 VSUBS 0.12fF $ **FLOATING
C248 S.t247 VSUBS 0.02fF
C249 S.n200 VSUBS 0.14fF $ **FLOATING
C250 S.t608 VSUBS 0.02fF
C251 S.n202 VSUBS 0.24fF $ **FLOATING
C252 S.n203 VSUBS 0.35fF $ **FLOATING
C253 S.n204 VSUBS 0.60fF $ **FLOATING
C254 S.n205 VSUBS 2.45fF $ **FLOATING
C255 S.n206 VSUBS 1.94fF $ **FLOATING
C256 S.t743 VSUBS 0.02fF
C257 S.n207 VSUBS 0.24fF $ **FLOATING
C258 S.n208 VSUBS 0.90fF $ **FLOATING
C259 S.n209 VSUBS 0.05fF $ **FLOATING
C260 S.t626 VSUBS 0.02fF
C261 S.n210 VSUBS 0.12fF $ **FLOATING
C262 S.n211 VSUBS 0.14fF $ **FLOATING
C263 S.n213 VSUBS 0.64fF $ **FLOATING
C264 S.n214 VSUBS 0.43fF $ **FLOATING
C265 S.n215 VSUBS 1.60fF $ **FLOATING
C266 S.n216 VSUBS 0.49fF $ **FLOATING
C267 S.n217 VSUBS 0.45fF $ **FLOATING
C268 S.n218 VSUBS 0.45fF $ **FLOATING
C269 S.n219 VSUBS 1.82fF $ **FLOATING
C270 S.n220 VSUBS 0.12fF $ **FLOATING
C271 S.t596 VSUBS 0.02fF
C272 S.n221 VSUBS 0.14fF $ **FLOATING
C273 S.t955 VSUBS 0.02fF
C274 S.n223 VSUBS 0.24fF $ **FLOATING
C275 S.n224 VSUBS 0.35fF $ **FLOATING
C276 S.n225 VSUBS 0.60fF $ **FLOATING
C277 S.n226 VSUBS 2.46fF $ **FLOATING
C278 S.n227 VSUBS 2.00fF $ **FLOATING
C279 S.t1078 VSUBS 0.02fF
C280 S.n228 VSUBS 0.24fF $ **FLOATING
C281 S.n229 VSUBS 0.90fF $ **FLOATING
C282 S.n230 VSUBS 0.05fF $ **FLOATING
C283 S.t976 VSUBS 0.02fF
C284 S.n231 VSUBS 0.12fF $ **FLOATING
C285 S.n232 VSUBS 0.14fF $ **FLOATING
C286 S.n234 VSUBS 0.18fF $ **FLOATING
C287 S.n235 VSUBS 0.09fF $ **FLOATING
C288 S.n236 VSUBS 0.93fF $ **FLOATING
C289 S.n237 VSUBS 0.46fF $ **FLOATING
C290 S.n238 VSUBS 0.76fF $ **FLOATING
C291 S.n239 VSUBS 0.21fF $ **FLOATING
C292 S.n240 VSUBS 0.35fF $ **FLOATING
C293 S.n241 VSUBS 0.53fF $ **FLOATING
C294 S.n242 VSUBS 1.60fF $ **FLOATING
C295 S.n243 VSUBS 0.12fF $ **FLOATING
C296 S.t944 VSUBS 0.02fF
C297 S.n244 VSUBS 0.14fF $ **FLOATING
C298 S.t193 VSUBS 0.02fF
C299 S.n246 VSUBS 0.24fF $ **FLOATING
C300 S.n247 VSUBS 0.35fF $ **FLOATING
C301 S.n248 VSUBS 0.60fF $ **FLOATING
C302 S.n249 VSUBS 2.45fF $ **FLOATING
C303 S.n250 VSUBS 1.94fF $ **FLOATING
C304 S.t310 VSUBS 0.02fF
C305 S.n251 VSUBS 0.24fF $ **FLOATING
C306 S.n252 VSUBS 0.90fF $ **FLOATING
C307 S.n253 VSUBS 0.05fF $ **FLOATING
C308 S.t216 VSUBS 0.02fF
C309 S.n254 VSUBS 0.12fF $ **FLOATING
C310 S.n255 VSUBS 0.14fF $ **FLOATING
C311 S.n257 VSUBS 0.64fF $ **FLOATING
C312 S.n258 VSUBS 0.43fF $ **FLOATING
C313 S.n259 VSUBS 1.60fF $ **FLOATING
C314 S.n260 VSUBS 0.49fF $ **FLOATING
C315 S.n261 VSUBS 0.45fF $ **FLOATING
C316 S.n262 VSUBS 0.45fF $ **FLOATING
C317 S.n263 VSUBS 1.82fF $ **FLOATING
C318 S.n264 VSUBS 0.12fF $ **FLOATING
C319 S.t186 VSUBS 0.02fF
C320 S.n265 VSUBS 0.14fF $ **FLOATING
C321 S.t544 VSUBS 0.02fF
C322 S.n267 VSUBS 0.24fF $ **FLOATING
C323 S.n268 VSUBS 0.35fF $ **FLOATING
C324 S.n269 VSUBS 0.60fF $ **FLOATING
C325 S.n270 VSUBS 2.46fF $ **FLOATING
C326 S.n271 VSUBS 2.00fF $ **FLOATING
C327 S.t657 VSUBS 0.02fF
C328 S.n272 VSUBS 0.24fF $ **FLOATING
C329 S.n273 VSUBS 0.90fF $ **FLOATING
C330 S.n274 VSUBS 0.05fF $ **FLOATING
C331 S.t567 VSUBS 0.02fF
C332 S.n275 VSUBS 0.12fF $ **FLOATING
C333 S.n276 VSUBS 0.14fF $ **FLOATING
C334 S.n278 VSUBS 0.18fF $ **FLOATING
C335 S.n279 VSUBS 0.09fF $ **FLOATING
C336 S.n280 VSUBS 0.93fF $ **FLOATING
C337 S.n281 VSUBS 0.46fF $ **FLOATING
C338 S.n282 VSUBS 0.76fF $ **FLOATING
C339 S.n283 VSUBS 0.21fF $ **FLOATING
C340 S.n284 VSUBS 0.35fF $ **FLOATING
C341 S.n285 VSUBS 0.53fF $ **FLOATING
C342 S.n286 VSUBS 1.60fF $ **FLOATING
C343 S.n287 VSUBS 0.12fF $ **FLOATING
C344 S.t865 VSUBS 0.02fF
C345 S.n288 VSUBS 0.14fF $ **FLOATING
C346 S.t774 VSUBS 0.02fF
C347 S.n290 VSUBS 0.24fF $ **FLOATING
C348 S.n291 VSUBS 0.35fF $ **FLOATING
C349 S.n292 VSUBS 0.60fF $ **FLOATING
C350 S.n293 VSUBS 2.45fF $ **FLOATING
C351 S.n294 VSUBS 1.94fF $ **FLOATING
C352 S.t3 VSUBS 0.02fF
C353 S.n295 VSUBS 0.24fF $ **FLOATING
C354 S.n296 VSUBS 0.90fF $ **FLOATING
C355 S.n297 VSUBS 0.05fF $ **FLOATING
C356 S.t962 VSUBS 0.02fF
C357 S.n298 VSUBS 0.12fF $ **FLOATING
C358 S.n299 VSUBS 0.14fF $ **FLOATING
C359 S.n301 VSUBS 1.87fF $ **FLOATING
C360 S.n302 VSUBS 0.12fF $ **FLOATING
C361 S.t105 VSUBS 0.02fF
C362 S.n303 VSUBS 0.14fF $ **FLOATING
C363 S.t630 VSUBS 0.02fF
C364 S.n305 VSUBS 1.20fF $ **FLOATING
C365 S.n306 VSUBS 2.27fF $ **FLOATING
C366 S.n307 VSUBS 0.60fF $ **FLOATING
C367 S.n308 VSUBS 0.35fF $ **FLOATING
C368 S.n309 VSUBS 0.62fF $ **FLOATING
C369 S.n310 VSUBS 1.14fF $ **FLOATING
C370 S.n311 VSUBS 2.15fF $ **FLOATING
C371 S.n312 VSUBS 0.59fF $ **FLOATING
C372 S.n313 VSUBS 0.01fF $ **FLOATING
C373 S.n314 VSUBS 0.96fF $ **FLOATING
C374 S.t6 VSUBS 14.53fF
C375 S.n315 VSUBS 14.40fF $ **FLOATING
C376 S.n317 VSUBS 0.37fF $ **FLOATING
C377 S.n318 VSUBS 0.23fF $ **FLOATING
C378 S.n319 VSUBS 2.85fF $ **FLOATING
C379 S.n320 VSUBS 2.43fF $ **FLOATING
C380 S.n321 VSUBS 4.25fF $ **FLOATING
C381 S.n322 VSUBS 0.25fF $ **FLOATING
C382 S.n323 VSUBS 0.01fF $ **FLOATING
C383 S.t274 VSUBS 0.02fF
C384 S.n324 VSUBS 0.25fF $ **FLOATING
C385 S.t771 VSUBS 0.02fF
C386 S.n325 VSUBS 0.94fF $ **FLOATING
C387 S.n326 VSUBS 0.70fF $ **FLOATING
C388 S.n327 VSUBS 1.87fF $ **FLOATING
C389 S.n328 VSUBS 1.76fF $ **FLOATING
C390 S.n329 VSUBS 0.12fF $ **FLOATING
C391 S.t673 VSUBS 0.02fF
C392 S.n330 VSUBS 0.14fF $ **FLOATING
C393 S.t980 VSUBS 0.02fF
C394 S.n332 VSUBS 0.24fF $ **FLOATING
C395 S.n333 VSUBS 0.35fF $ **FLOATING
C396 S.n334 VSUBS 0.60fF $ **FLOATING
C397 S.n335 VSUBS 2.71fF $ **FLOATING
C398 S.n336 VSUBS 2.03fF $ **FLOATING
C399 S.t1113 VSUBS 0.02fF
C400 S.n337 VSUBS 0.24fF $ **FLOATING
C401 S.n338 VSUBS 0.90fF $ **FLOATING
C402 S.n339 VSUBS 0.05fF $ **FLOATING
C403 S.t1000 VSUBS 0.02fF
C404 S.n340 VSUBS 0.12fF $ **FLOATING
C405 S.n341 VSUBS 0.14fF $ **FLOATING
C406 S.n343 VSUBS 1.23fF $ **FLOATING
C407 S.n344 VSUBS 1.27fF $ **FLOATING
C408 S.n345 VSUBS 1.86fF $ **FLOATING
C409 S.n346 VSUBS 0.12fF $ **FLOATING
C410 S.t518 VSUBS 0.02fF
C411 S.n347 VSUBS 0.14fF $ **FLOATING
C412 S.t874 VSUBS 0.02fF
C413 S.n349 VSUBS 0.24fF $ **FLOATING
C414 S.n350 VSUBS 0.35fF $ **FLOATING
C415 S.n351 VSUBS 0.60fF $ **FLOATING
C416 S.n352 VSUBS 2.72fF $ **FLOATING
C417 S.n353 VSUBS 2.14fF $ **FLOATING
C418 S.t987 VSUBS 0.02fF
C419 S.n354 VSUBS 0.24fF $ **FLOATING
C420 S.n355 VSUBS 0.90fF $ **FLOATING
C421 S.n356 VSUBS 0.05fF $ **FLOATING
C422 S.t292 VSUBS 0.02fF
C423 S.n357 VSUBS 0.12fF $ **FLOATING
C424 S.n358 VSUBS 0.14fF $ **FLOATING
C425 S.n360 VSUBS 1.87fF $ **FLOATING
C426 S.n361 VSUBS 1.78fF $ **FLOATING
C427 S.n362 VSUBS 0.12fF $ **FLOATING
C428 S.t860 VSUBS 0.02fF
C429 S.n363 VSUBS 0.14fF $ **FLOATING
C430 S.t102 VSUBS 0.02fF
C431 S.n365 VSUBS 0.24fF $ **FLOATING
C432 S.n366 VSUBS 0.35fF $ **FLOATING
C433 S.n367 VSUBS 0.60fF $ **FLOATING
C434 S.n368 VSUBS 2.70fF $ **FLOATING
C435 S.n369 VSUBS 2.03fF $ **FLOATING
C436 S.t226 VSUBS 0.02fF
C437 S.n370 VSUBS 0.24fF $ **FLOATING
C438 S.n371 VSUBS 0.90fF $ **FLOATING
C439 S.n372 VSUBS 0.05fF $ **FLOATING
C440 S.t125 VSUBS 0.02fF
C441 S.n373 VSUBS 0.12fF $ **FLOATING
C442 S.n374 VSUBS 0.14fF $ **FLOATING
C443 S.n376 VSUBS 1.23fF $ **FLOATING
C444 S.n377 VSUBS 1.27fF $ **FLOATING
C445 S.n378 VSUBS 1.86fF $ **FLOATING
C446 S.n379 VSUBS 0.12fF $ **FLOATING
C447 S.t87 VSUBS 0.02fF
C448 S.n380 VSUBS 0.14fF $ **FLOATING
C449 S.t462 VSUBS 0.02fF
C450 S.n382 VSUBS 0.24fF $ **FLOATING
C451 S.n383 VSUBS 0.35fF $ **FLOATING
C452 S.n384 VSUBS 0.60fF $ **FLOATING
C453 S.n385 VSUBS 2.72fF $ **FLOATING
C454 S.n386 VSUBS 2.14fF $ **FLOATING
C455 S.t578 VSUBS 0.02fF
C456 S.n387 VSUBS 0.24fF $ **FLOATING
C457 S.n388 VSUBS 0.90fF $ **FLOATING
C458 S.n389 VSUBS 0.05fF $ **FLOATING
C459 S.t483 VSUBS 0.02fF
C460 S.n390 VSUBS 0.12fF $ **FLOATING
C461 S.n391 VSUBS 0.14fF $ **FLOATING
C462 S.n393 VSUBS 1.87fF $ **FLOATING
C463 S.n394 VSUBS 1.78fF $ **FLOATING
C464 S.n395 VSUBS 0.12fF $ **FLOATING
C465 S.t451 VSUBS 0.02fF
C466 S.n396 VSUBS 0.14fF $ **FLOATING
C467 S.t799 VSUBS 0.02fF
C468 S.n398 VSUBS 0.24fF $ **FLOATING
C469 S.n399 VSUBS 0.35fF $ **FLOATING
C470 S.n400 VSUBS 0.60fF $ **FLOATING
C471 S.n401 VSUBS 2.70fF $ **FLOATING
C472 S.n402 VSUBS 2.03fF $ **FLOATING
C473 S.t921 VSUBS 0.02fF
C474 S.n403 VSUBS 0.24fF $ **FLOATING
C475 S.n404 VSUBS 0.90fF $ **FLOATING
C476 S.n405 VSUBS 0.05fF $ **FLOATING
C477 S.t826 VSUBS 0.02fF
C478 S.n406 VSUBS 0.12fF $ **FLOATING
C479 S.n407 VSUBS 0.14fF $ **FLOATING
C480 S.n409 VSUBS 1.23fF $ **FLOATING
C481 S.n410 VSUBS 1.27fF $ **FLOATING
C482 S.n411 VSUBS 1.86fF $ **FLOATING
C483 S.n412 VSUBS 0.12fF $ **FLOATING
C484 S.t848 VSUBS 0.02fF
C485 S.n413 VSUBS 0.14fF $ **FLOATING
C486 S.t7 VSUBS 0.02fF
C487 S.n415 VSUBS 0.24fF $ **FLOATING
C488 S.n416 VSUBS 0.35fF $ **FLOATING
C489 S.n417 VSUBS 0.60fF $ **FLOATING
C490 S.n418 VSUBS 2.72fF $ **FLOATING
C491 S.n419 VSUBS 2.14fF $ **FLOATING
C492 S.t163 VSUBS 0.02fF
C493 S.n420 VSUBS 0.24fF $ **FLOATING
C494 S.n421 VSUBS 0.90fF $ **FLOATING
C495 S.n422 VSUBS 0.05fF $ **FLOATING
C496 S.t40 VSUBS 0.02fF
C497 S.n423 VSUBS 0.12fF $ **FLOATING
C498 S.n424 VSUBS 0.14fF $ **FLOATING
C499 S.n426 VSUBS 2.58fF $ **FLOATING
C500 S.n427 VSUBS 1.86fF $ **FLOATING
C501 S.n428 VSUBS 0.12fF $ **FLOATING
C502 S.t464 VSUBS 0.02fF
C503 S.n429 VSUBS 0.14fF $ **FLOATING
C504 S.t369 VSUBS 0.02fF
C505 S.n431 VSUBS 0.24fF $ **FLOATING
C506 S.n432 VSUBS 0.35fF $ **FLOATING
C507 S.n433 VSUBS 0.60fF $ **FLOATING
C508 S.n434 VSUBS 0.89fF $ **FLOATING
C509 S.n435 VSUBS 0.76fF $ **FLOATING
C510 S.n436 VSUBS 0.96fF $ **FLOATING
C511 S.n437 VSUBS 0.09fF $ **FLOATING
C512 S.n438 VSUBS 0.32fF $ **FLOATING
C513 S.n439 VSUBS 2.13fF $ **FLOATING
C514 S.t735 VSUBS 0.02fF
C515 S.n440 VSUBS 0.24fF $ **FLOATING
C516 S.n441 VSUBS 0.90fF $ **FLOATING
C517 S.n442 VSUBS 0.05fF $ **FLOATING
C518 S.t841 VSUBS 0.02fF
C519 S.n443 VSUBS 0.12fF $ **FLOATING
C520 S.n444 VSUBS 0.14fF $ **FLOATING
C521 S.n446 VSUBS 2.27fF $ **FLOATING
C522 S.n447 VSUBS 1.86fF $ **FLOATING
C523 S.n448 VSUBS 0.12fF $ **FLOATING
C524 S.t802 VSUBS 0.02fF
C525 S.n449 VSUBS 0.14fF $ **FLOATING
C526 S.t701 VSUBS 0.02fF
C527 S.n451 VSUBS 0.24fF $ **FLOATING
C528 S.n452 VSUBS 0.35fF $ **FLOATING
C529 S.n453 VSUBS 0.60fF $ **FLOATING
C530 S.n454 VSUBS 0.76fF $ **FLOATING
C531 S.n455 VSUBS 0.48fF $ **FLOATING
C532 S.n456 VSUBS 0.09fF $ **FLOATING
C533 S.n457 VSUBS 0.32fF $ **FLOATING
C534 S.n458 VSUBS 2.00fF $ **FLOATING
C535 S.t1068 VSUBS 0.02fF
C536 S.n459 VSUBS 0.24fF $ **FLOATING
C537 S.n460 VSUBS 0.90fF $ **FLOATING
C538 S.n461 VSUBS 0.05fF $ **FLOATING
C539 S.t61 VSUBS 0.02fF
C540 S.n462 VSUBS 0.12fF $ **FLOATING
C541 S.n463 VSUBS 0.14fF $ **FLOATING
C542 S.n465 VSUBS 1.87fF $ **FLOATING
C543 S.n466 VSUBS 1.14fF $ **FLOATING
C544 S.n467 VSUBS 0.22fF $ **FLOATING
C545 S.n468 VSUBS 0.12fF $ **FLOATING
C546 S.t13 VSUBS 0.02fF
C547 S.n469 VSUBS 0.14fF $ **FLOATING
C548 S.t1045 VSUBS 0.02fF
C549 S.n471 VSUBS 0.24fF $ **FLOATING
C550 S.n472 VSUBS 0.35fF $ **FLOATING
C551 S.n473 VSUBS 0.60fF $ **FLOATING
C552 S.n474 VSUBS 2.70fF $ **FLOATING
C553 S.n475 VSUBS 1.86fF $ **FLOATING
C554 S.t308 VSUBS 0.02fF
C555 S.n476 VSUBS 0.24fF $ **FLOATING
C556 S.n477 VSUBS 0.90fF $ **FLOATING
C557 S.n478 VSUBS 0.05fF $ **FLOATING
C558 S.t427 VSUBS 0.02fF
C559 S.n479 VSUBS 0.12fF $ **FLOATING
C560 S.n480 VSUBS 0.14fF $ **FLOATING
C561 S.n482 VSUBS 14.09fF $ **FLOATING
C562 S.n483 VSUBS 2.69fF $ **FLOATING
C563 S.n484 VSUBS 1.94fF $ **FLOATING
C564 S.n485 VSUBS 0.12fF $ **FLOATING
C565 S.t146 VSUBS 0.02fF
C566 S.n486 VSUBS 0.14fF $ **FLOATING
C567 S.t825 VSUBS 0.02fF
C568 S.n488 VSUBS 0.24fF $ **FLOATING
C569 S.n489 VSUBS 0.35fF $ **FLOATING
C570 S.n490 VSUBS 0.60fF $ **FLOATING
C571 S.n491 VSUBS 1.55fF $ **FLOATING
C572 S.n492 VSUBS 0.28fF $ **FLOATING
C573 S.n493 VSUBS 2.08fF $ **FLOATING
C574 S.t769 VSUBS 0.02fF
C575 S.n494 VSUBS 0.12fF $ **FLOATING
C576 S.n495 VSUBS 0.14fF $ **FLOATING
C577 S.t321 VSUBS 0.02fF
C578 S.n497 VSUBS 0.24fF $ **FLOATING
C579 S.n498 VSUBS 0.90fF $ **FLOATING
C580 S.n499 VSUBS 0.05fF $ **FLOATING
C581 S.t12 VSUBS 32.33fF
C582 S.t503 VSUBS 0.02fF
C583 S.n500 VSUBS 0.12fF $ **FLOATING
C584 S.n501 VSUBS 0.14fF $ **FLOATING
C585 S.t397 VSUBS 0.02fF
C586 S.n503 VSUBS 0.24fF $ **FLOATING
C587 S.n504 VSUBS 0.90fF $ **FLOATING
C588 S.n505 VSUBS 0.05fF $ **FLOATING
C589 S.t1130 VSUBS 0.02fF
C590 S.n506 VSUBS 0.24fF $ **FLOATING
C591 S.n507 VSUBS 0.35fF $ **FLOATING
C592 S.n508 VSUBS 0.60fF $ **FLOATING
C593 S.n509 VSUBS 2.21fF $ **FLOATING
C594 S.n510 VSUBS 2.66fF $ **FLOATING
C595 S.n511 VSUBS 2.62fF $ **FLOATING
C596 S.n512 VSUBS 2.34fF $ **FLOATING
C597 S.n513 VSUBS 1.84fF $ **FLOATING
C598 S.n514 VSUBS 0.12fF $ **FLOATING
C599 S.t90 VSUBS 0.02fF
C600 S.n515 VSUBS 0.14fF $ **FLOATING
C601 S.t1119 VSUBS 0.02fF
C602 S.n517 VSUBS 0.24fF $ **FLOATING
C603 S.n518 VSUBS 0.35fF $ **FLOATING
C604 S.n519 VSUBS 0.60fF $ **FLOATING
C605 S.n520 VSUBS 0.40fF $ **FLOATING
C606 S.n521 VSUBS 0.66fF $ **FLOATING
C607 S.n522 VSUBS 0.54fF $ **FLOATING
C608 S.n523 VSUBS 0.32fF $ **FLOATING
C609 S.n524 VSUBS 1.06fF $ **FLOATING
C610 S.n525 VSUBS 2.10fF $ **FLOATING
C611 S.t381 VSUBS 0.02fF
C612 S.n526 VSUBS 0.24fF $ **FLOATING
C613 S.n527 VSUBS 0.90fF $ **FLOATING
C614 S.n528 VSUBS 0.05fF $ **FLOATING
C615 S.t487 VSUBS 0.02fF
C616 S.n529 VSUBS 0.12fF $ **FLOATING
C617 S.n530 VSUBS 0.14fF $ **FLOATING
C618 S.n532 VSUBS 0.03fF $ **FLOATING
C619 S.n533 VSUBS 0.03fF $ **FLOATING
C620 S.n534 VSUBS 0.10fF $ **FLOATING
C621 S.n535 VSUBS 0.36fF $ **FLOATING
C622 S.n536 VSUBS 0.37fF $ **FLOATING
C623 S.n537 VSUBS 0.10fF $ **FLOATING
C624 S.n538 VSUBS 0.12fF $ **FLOATING
C625 S.n539 VSUBS 0.03fF $ **FLOATING
C626 S.n540 VSUBS 0.07fF $ **FLOATING
C627 S.n541 VSUBS 1.39fF $ **FLOATING
C628 S.n542 VSUBS 0.04fF $ **FLOATING
C629 S.n543 VSUBS 0.48fF $ **FLOATING
C630 S.n544 VSUBS 0.37fF $ **FLOATING
C631 S.n545 VSUBS 1.60fF $ **FLOATING
C632 S.n546 VSUBS 0.12fF $ **FLOATING
C633 S.t452 VSUBS 0.02fF
C634 S.n547 VSUBS 0.14fF $ **FLOATING
C635 S.t350 VSUBS 0.02fF
C636 S.n549 VSUBS 0.24fF $ **FLOATING
C637 S.n550 VSUBS 0.35fF $ **FLOATING
C638 S.n551 VSUBS 0.60fF $ **FLOATING
C639 S.n552 VSUBS 0.35fF $ **FLOATING
C640 S.n553 VSUBS 0.53fF $ **FLOATING
C641 S.n554 VSUBS 0.38fF $ **FLOATING
C642 S.n555 VSUBS 0.18fF $ **FLOATING
C643 S.n556 VSUBS 0.25fF $ **FLOATING
C644 S.n557 VSUBS 0.09fF $ **FLOATING
C645 S.n558 VSUBS 1.94fF $ **FLOATING
C646 S.t722 VSUBS 0.02fF
C647 S.n559 VSUBS 0.24fF $ **FLOATING
C648 S.n560 VSUBS 0.90fF $ **FLOATING
C649 S.n561 VSUBS 0.05fF $ **FLOATING
C650 S.t829 VSUBS 0.02fF
C651 S.n562 VSUBS 0.12fF $ **FLOATING
C652 S.n563 VSUBS 0.14fF $ **FLOATING
C653 S.n565 VSUBS 1.48fF $ **FLOATING
C654 S.n566 VSUBS 0.25fF $ **FLOATING
C655 S.n567 VSUBS 0.09fF $ **FLOATING
C656 S.n568 VSUBS 0.77fF $ **FLOATING
C657 S.n569 VSUBS 0.21fF $ **FLOATING
C658 S.n570 VSUBS 1.71fF $ **FLOATING
C659 S.n571 VSUBS 0.44fF $ **FLOATING
C660 S.n572 VSUBS 0.12fF $ **FLOATING
C661 S.t794 VSUBS 0.02fF
C662 S.n573 VSUBS 0.14fF $ **FLOATING
C663 S.t689 VSUBS 0.02fF
C664 S.n575 VSUBS 0.24fF $ **FLOATING
C665 S.n576 VSUBS 0.35fF $ **FLOATING
C666 S.n577 VSUBS 0.60fF $ **FLOATING
C667 S.n578 VSUBS 0.82fF $ **FLOATING
C668 S.n579 VSUBS 0.29fF $ **FLOATING
C669 S.n580 VSUBS 0.25fF $ **FLOATING
C670 S.n581 VSUBS 0.31fF $ **FLOATING
C671 S.n582 VSUBS 0.22fF $ **FLOATING
C672 S.n583 VSUBS 0.60fF $ **FLOATING
C673 S.n584 VSUBS 0.27fF $ **FLOATING
C674 S.n585 VSUBS 0.14fF $ **FLOATING
C675 S.n586 VSUBS 1.72fF $ **FLOATING
C676 S.n587 VSUBS 1.91fF $ **FLOATING
C677 S.t1059 VSUBS 0.02fF
C678 S.n588 VSUBS 0.24fF $ **FLOATING
C679 S.n589 VSUBS 0.90fF $ **FLOATING
C680 S.n590 VSUBS 0.05fF $ **FLOATING
C681 S.t49 VSUBS 0.02fF
C682 S.n591 VSUBS 0.12fF $ **FLOATING
C683 S.n592 VSUBS 0.14fF $ **FLOATING
C684 S.n594 VSUBS 0.19fF $ **FLOATING
C685 S.n595 VSUBS 0.09fF $ **FLOATING
C686 S.n596 VSUBS 0.67fF $ **FLOATING
C687 S.n597 VSUBS 0.28fF $ **FLOATING
C688 S.n598 VSUBS 1.72fF $ **FLOATING
C689 S.n599 VSUBS 0.21fF $ **FLOATING
C690 S.n600 VSUBS 1.82fF $ **FLOATING
C691 S.n601 VSUBS 0.12fF $ **FLOATING
C692 S.t1136 VSUBS 0.02fF
C693 S.n602 VSUBS 0.14fF $ **FLOATING
C694 S.t1034 VSUBS 0.02fF
C695 S.n604 VSUBS 0.24fF $ **FLOATING
C696 S.n605 VSUBS 0.35fF $ **FLOATING
C697 S.n606 VSUBS 0.60fF $ **FLOATING
C698 S.n607 VSUBS 2.46fF $ **FLOATING
C699 S.n608 VSUBS 1.84fF $ **FLOATING
C700 S.t300 VSUBS 0.02fF
C701 S.n609 VSUBS 0.24fF $ **FLOATING
C702 S.n610 VSUBS 0.90fF $ **FLOATING
C703 S.n611 VSUBS 0.05fF $ **FLOATING
C704 S.t416 VSUBS 0.02fF
C705 S.n612 VSUBS 0.12fF $ **FLOATING
C706 S.n613 VSUBS 0.14fF $ **FLOATING
C707 S.n615 VSUBS 0.06fF $ **FLOATING
C708 S.n616 VSUBS 0.20fF $ **FLOATING
C709 S.n617 VSUBS 0.09fF $ **FLOATING
C710 S.n618 VSUBS 0.20fF $ **FLOATING
C711 S.n619 VSUBS 0.09fF $ **FLOATING
C712 S.n620 VSUBS 0.30fF $ **FLOATING
C713 S.n621 VSUBS 0.99fF $ **FLOATING
C714 S.n622 VSUBS 0.44fF $ **FLOATING
C715 S.n623 VSUBS 2.05fF $ **FLOATING
C716 S.n624 VSUBS 0.12fF $ **FLOATING
C717 S.t1137 VSUBS 0.02fF
C718 S.n625 VSUBS 0.14fF $ **FLOATING
C719 S.t390 VSUBS 0.02fF
C720 S.n627 VSUBS 0.24fF $ **FLOATING
C721 S.n628 VSUBS 0.35fF $ **FLOATING
C722 S.n629 VSUBS 0.60fF $ **FLOATING
C723 S.n630 VSUBS 0.43fF $ **FLOATING
C724 S.n631 VSUBS 0.78fF $ **FLOATING
C725 S.n632 VSUBS 0.18fF $ **FLOATING
C726 S.n633 VSUBS 0.95fF $ **FLOATING
C727 S.n634 VSUBS 0.39fF $ **FLOATING
C728 S.n635 VSUBS 0.44fF $ **FLOATING
C729 S.n636 VSUBS 0.25fF $ **FLOATING
C730 S.n637 VSUBS 0.09fF $ **FLOATING
C731 S.n638 VSUBS 1.79fF $ **FLOATING
C732 S.t420 VSUBS 0.02fF
C733 S.n639 VSUBS 0.12fF $ **FLOATING
C734 S.n640 VSUBS 0.14fF $ **FLOATING
C735 S.t517 VSUBS 0.02fF
C736 S.n642 VSUBS 0.24fF $ **FLOATING
C737 S.n643 VSUBS 0.90fF $ **FLOATING
C738 S.n644 VSUBS 0.05fF $ **FLOATING
C739 S.t48 VSUBS 31.95fF
C740 S.t754 VSUBS 0.02fF
C741 S.n645 VSUBS 0.01fF $ **FLOATING
C742 S.n646 VSUBS 0.25fF $ **FLOATING
C743 S.t400 VSUBS 0.02fF
C744 S.n648 VSUBS 1.18fF $ **FLOATING
C745 S.n649 VSUBS 0.05fF $ **FLOATING
C746 S.t254 VSUBS 0.02fF
C747 S.n650 VSUBS 0.63fF $ **FLOATING
C748 S.n651 VSUBS 0.60fF $ **FLOATING
C749 S.n652 VSUBS 8.88fF $ **FLOATING
C750 S.n653 VSUBS 20.14fF $ **FLOATING
C751 S.n654 VSUBS 8.88fF $ **FLOATING
C752 S.n655 VSUBS 20.14fF $ **FLOATING
C753 S.n656 VSUBS 0.59fF $ **FLOATING
C754 S.n657 VSUBS 0.21fF $ **FLOATING
C755 S.n658 VSUBS 0.87fF $ **FLOATING
C756 S.n659 VSUBS 0.87fF $ **FLOATING
C757 S.n660 VSUBS 2.55fF $ **FLOATING
C758 S.n661 VSUBS 0.28fF $ **FLOATING
C759 S.t162 VSUBS 14.53fF
C760 S.n662 VSUBS 15.80fF $ **FLOATING
C761 S.n663 VSUBS 0.21fF $ **FLOATING
C762 S.n664 VSUBS 1.40fF $ **FLOATING
C763 S.n665 VSUBS 4.20fF $ **FLOATING
C764 S.n666 VSUBS 1.12fF $ **FLOATING
C765 S.n667 VSUBS 1.78fF $ **FLOATING
C766 S.n668 VSUBS 4.18fF $ **FLOATING
C767 S.n669 VSUBS 0.24fF $ **FLOATING
C768 S.n670 VSUBS 1.48fF $ **FLOATING
C769 S.n671 VSUBS 1.29fF $ **FLOATING
C770 S.n672 VSUBS 0.27fF $ **FLOATING
C771 S.n673 VSUBS 1.86fF $ **FLOATING
C772 S.n674 VSUBS 0.25fF $ **FLOATING
C773 S.n675 VSUBS 0.09fF $ **FLOATING
C774 S.n676 VSUBS 0.21fF $ **FLOATING
C775 S.n677 VSUBS 0.79fF $ **FLOATING
C776 S.n678 VSUBS 0.44fF $ **FLOATING
C777 S.n679 VSUBS 0.12fF $ **FLOATING
C778 S.t176 VSUBS 0.02fF
C779 S.n680 VSUBS 0.14fF $ **FLOATING
C780 S.t419 VSUBS 0.02fF
C781 S.n682 VSUBS 0.24fF $ **FLOATING
C782 S.n683 VSUBS 0.35fF $ **FLOATING
C783 S.n684 VSUBS 0.60fF $ **FLOATING
C784 S.n685 VSUBS 0.02fF $ **FLOATING
C785 S.n686 VSUBS 0.01fF $ **FLOATING
C786 S.n687 VSUBS 0.02fF $ **FLOATING
C787 S.n688 VSUBS 0.08fF $ **FLOATING
C788 S.n689 VSUBS 0.06fF $ **FLOATING
C789 S.n690 VSUBS 0.03fF $ **FLOATING
C790 S.n691 VSUBS 0.03fF $ **FLOATING
C791 S.n692 VSUBS 0.99fF $ **FLOATING
C792 S.n693 VSUBS 0.36fF $ **FLOATING
C793 S.n694 VSUBS 1.83fF $ **FLOATING
C794 S.n695 VSUBS 1.96fF $ **FLOATING
C795 S.t651 VSUBS 0.02fF
C796 S.n696 VSUBS 0.24fF $ **FLOATING
C797 S.n697 VSUBS 0.90fF $ **FLOATING
C798 S.n698 VSUBS 0.05fF $ **FLOATING
C799 S.t560 VSUBS 0.02fF
C800 S.n699 VSUBS 0.12fF $ **FLOATING
C801 S.n700 VSUBS 0.14fF $ **FLOATING
C802 S.n702 VSUBS 1.87fF $ **FLOATING
C803 S.n703 VSUBS 0.06fF $ **FLOATING
C804 S.n704 VSUBS 0.03fF $ **FLOATING
C805 S.n705 VSUBS 0.03fF $ **FLOATING
C806 S.n706 VSUBS 0.98fF $ **FLOATING
C807 S.n707 VSUBS 0.02fF $ **FLOATING
C808 S.n708 VSUBS 0.01fF $ **FLOATING
C809 S.n709 VSUBS 0.02fF $ **FLOATING
C810 S.n710 VSUBS 0.08fF $ **FLOATING
C811 S.n711 VSUBS 0.35fF $ **FLOATING
C812 S.n712 VSUBS 1.84fF $ **FLOATING
C813 S.t233 VSUBS 0.02fF
C814 S.n713 VSUBS 0.24fF $ **FLOATING
C815 S.n714 VSUBS 0.35fF $ **FLOATING
C816 S.n715 VSUBS 0.60fF $ **FLOATING
C817 S.n716 VSUBS 0.12fF $ **FLOATING
C818 S.t1115 VSUBS 0.02fF
C819 S.n717 VSUBS 0.14fF $ **FLOATING
C820 S.n719 VSUBS 0.94fF $ **FLOATING
C821 S.n720 VSUBS 0.58fF $ **FLOATING
C822 S.n721 VSUBS 0.25fF $ **FLOATING
C823 S.n722 VSUBS 0.69fF $ **FLOATING
C824 S.n723 VSUBS 0.22fF $ **FLOATING
C825 S.n724 VSUBS 0.09fF $ **FLOATING
C826 S.n725 VSUBS 1.86fF $ **FLOATING
C827 S.t501 VSUBS 0.02fF
C828 S.n726 VSUBS 0.24fF $ **FLOATING
C829 S.n727 VSUBS 0.90fF $ **FLOATING
C830 S.n728 VSUBS 0.05fF $ **FLOATING
C831 S.t391 VSUBS 0.02fF
C832 S.n729 VSUBS 0.12fF $ **FLOATING
C833 S.n730 VSUBS 0.14fF $ **FLOATING
C834 S.n732 VSUBS 1.86fF $ **FLOATING
C835 S.n733 VSUBS 0.25fF $ **FLOATING
C836 S.n734 VSUBS 0.09fF $ **FLOATING
C837 S.n735 VSUBS 0.21fF $ **FLOATING
C838 S.n736 VSUBS 0.79fF $ **FLOATING
C839 S.n737 VSUBS 0.44fF $ **FLOATING
C840 S.n738 VSUBS 0.12fF $ **FLOATING
C841 S.t346 VSUBS 0.02fF
C842 S.n739 VSUBS 0.14fF $ **FLOATING
C843 S.t582 VSUBS 0.02fF
C844 S.n741 VSUBS 0.24fF $ **FLOATING
C845 S.n742 VSUBS 0.35fF $ **FLOATING
C846 S.n743 VSUBS 0.60fF $ **FLOATING
C847 S.n744 VSUBS 0.02fF $ **FLOATING
C848 S.n745 VSUBS 0.01fF $ **FLOATING
C849 S.n746 VSUBS 0.02fF $ **FLOATING
C850 S.n747 VSUBS 0.08fF $ **FLOATING
C851 S.n748 VSUBS 0.06fF $ **FLOATING
C852 S.n749 VSUBS 0.03fF $ **FLOATING
C853 S.n750 VSUBS 0.03fF $ **FLOATING
C854 S.n751 VSUBS 0.99fF $ **FLOATING
C855 S.n752 VSUBS 0.36fF $ **FLOATING
C856 S.n753 VSUBS 1.83fF $ **FLOATING
C857 S.n754 VSUBS 1.96fF $ **FLOATING
C858 S.t839 VSUBS 0.02fF
C859 S.n755 VSUBS 0.24fF $ **FLOATING
C860 S.n756 VSUBS 0.90fF $ **FLOATING
C861 S.n757 VSUBS 0.05fF $ **FLOATING
C862 S.t730 VSUBS 0.02fF
C863 S.n758 VSUBS 0.12fF $ **FLOATING
C864 S.n759 VSUBS 0.14fF $ **FLOATING
C865 S.n761 VSUBS 1.87fF $ **FLOATING
C866 S.n762 VSUBS 0.06fF $ **FLOATING
C867 S.n763 VSUBS 0.03fF $ **FLOATING
C868 S.n764 VSUBS 0.03fF $ **FLOATING
C869 S.n765 VSUBS 0.98fF $ **FLOATING
C870 S.n766 VSUBS 0.02fF $ **FLOATING
C871 S.n767 VSUBS 0.01fF $ **FLOATING
C872 S.n768 VSUBS 0.02fF $ **FLOATING
C873 S.n769 VSUBS 0.08fF $ **FLOATING
C874 S.n770 VSUBS 0.35fF $ **FLOATING
C875 S.n771 VSUBS 1.84fF $ **FLOATING
C876 S.t927 VSUBS 0.02fF
C877 S.n772 VSUBS 0.24fF $ **FLOATING
C878 S.n773 VSUBS 0.35fF $ **FLOATING
C879 S.n774 VSUBS 0.60fF $ **FLOATING
C880 S.n775 VSUBS 0.12fF $ **FLOATING
C881 S.t685 VSUBS 0.02fF
C882 S.n776 VSUBS 0.14fF $ **FLOATING
C883 S.n778 VSUBS 0.94fF $ **FLOATING
C884 S.n779 VSUBS 0.58fF $ **FLOATING
C885 S.n780 VSUBS 0.25fF $ **FLOATING
C886 S.n781 VSUBS 0.69fF $ **FLOATING
C887 S.n782 VSUBS 0.22fF $ **FLOATING
C888 S.n783 VSUBS 0.09fF $ **FLOATING
C889 S.n784 VSUBS 1.86fF $ **FLOATING
C890 S.t59 VSUBS 0.02fF
C891 S.n785 VSUBS 0.24fF $ **FLOATING
C892 S.n786 VSUBS 0.90fF $ **FLOATING
C893 S.n787 VSUBS 0.05fF $ **FLOATING
C894 S.t1065 VSUBS 0.02fF
C895 S.n788 VSUBS 0.12fF $ **FLOATING
C896 S.n789 VSUBS 0.14fF $ **FLOATING
C897 S.n791 VSUBS 1.86fF $ **FLOATING
C898 S.n792 VSUBS 0.25fF $ **FLOATING
C899 S.n793 VSUBS 0.09fF $ **FLOATING
C900 S.n794 VSUBS 0.21fF $ **FLOATING
C901 S.n795 VSUBS 0.79fF $ **FLOATING
C902 S.n796 VSUBS 0.44fF $ **FLOATING
C903 S.n797 VSUBS 0.12fF $ **FLOATING
C904 S.t1030 VSUBS 0.02fF
C905 S.n798 VSUBS 0.14fF $ **FLOATING
C906 S.t167 VSUBS 0.02fF
C907 S.n800 VSUBS 0.24fF $ **FLOATING
C908 S.n801 VSUBS 0.35fF $ **FLOATING
C909 S.n802 VSUBS 0.60fF $ **FLOATING
C910 S.n803 VSUBS 0.02fF $ **FLOATING
C911 S.n804 VSUBS 0.01fF $ **FLOATING
C912 S.n805 VSUBS 0.02fF $ **FLOATING
C913 S.n806 VSUBS 0.08fF $ **FLOATING
C914 S.n807 VSUBS 0.03fF $ **FLOATING
C915 S.n808 VSUBS 0.03fF $ **FLOATING
C916 S.n809 VSUBS 1.01fF $ **FLOATING
C917 S.n810 VSUBS 0.36fF $ **FLOATING
C918 S.n811 VSUBS 1.83fF $ **FLOATING
C919 S.n812 VSUBS 1.96fF $ **FLOATING
C920 S.t425 VSUBS 0.02fF
C921 S.n813 VSUBS 0.24fF $ **FLOATING
C922 S.n814 VSUBS 0.90fF $ **FLOATING
C923 S.n815 VSUBS 0.05fF $ **FLOATING
C924 S.t305 VSUBS 0.02fF
C925 S.n816 VSUBS 0.12fF $ **FLOATING
C926 S.n817 VSUBS 0.14fF $ **FLOATING
C927 S.n819 VSUBS 0.25fF $ **FLOATING
C928 S.n820 VSUBS 0.09fF $ **FLOATING
C929 S.n821 VSUBS 0.69fF $ **FLOATING
C930 S.n822 VSUBS 0.22fF $ **FLOATING
C931 S.n823 VSUBS 0.94fF $ **FLOATING
C932 S.n824 VSUBS 0.58fF $ **FLOATING
C933 S.n825 VSUBS 1.87fF $ **FLOATING
C934 S.n826 VSUBS 0.12fF $ **FLOATING
C935 S.t117 VSUBS 0.02fF
C936 S.n827 VSUBS 0.14fF $ **FLOATING
C937 S.t417 VSUBS 0.02fF
C938 S.n829 VSUBS 0.24fF $ **FLOATING
C939 S.n830 VSUBS 0.35fF $ **FLOATING
C940 S.n831 VSUBS 0.60fF $ **FLOATING
C941 S.n832 VSUBS 0.18fF $ **FLOATING
C942 S.n833 VSUBS 0.21fF $ **FLOATING
C943 S.n834 VSUBS 0.47fF $ **FLOATING
C944 S.n835 VSUBS 0.33fF $ **FLOATING
C945 S.n836 VSUBS 0.01fF $ **FLOATING
C946 S.n837 VSUBS 0.01fF $ **FLOATING
C947 S.n838 VSUBS 0.01fF $ **FLOATING
C948 S.n839 VSUBS 0.07fF $ **FLOATING
C949 S.n840 VSUBS 0.07fF $ **FLOATING
C950 S.n841 VSUBS 0.04fF $ **FLOATING
C951 S.n842 VSUBS 0.05fF $ **FLOATING
C952 S.n843 VSUBS 0.41fF $ **FLOATING
C953 S.n844 VSUBS 0.57fF $ **FLOATING
C954 S.n845 VSUBS 0.19fF $ **FLOATING
C955 S.n846 VSUBS 1.94fF $ **FLOATING
C956 S.t410 VSUBS 0.02fF
C957 S.n847 VSUBS 0.24fF $ **FLOATING
C958 S.n848 VSUBS 0.90fF $ **FLOATING
C959 S.n849 VSUBS 0.05fF $ **FLOATING
C960 S.t712 VSUBS 0.02fF
C961 S.n850 VSUBS 0.12fF $ **FLOATING
C962 S.n851 VSUBS 0.14fF $ **FLOATING
C963 S.n853 VSUBS 0.04fF $ **FLOATING
C964 S.n854 VSUBS 0.03fF $ **FLOATING
C965 S.n855 VSUBS 0.03fF $ **FLOATING
C966 S.n856 VSUBS 0.10fF $ **FLOATING
C967 S.n857 VSUBS 0.36fF $ **FLOATING
C968 S.n858 VSUBS 0.37fF $ **FLOATING
C969 S.n859 VSUBS 0.10fF $ **FLOATING
C970 S.n860 VSUBS 0.12fF $ **FLOATING
C971 S.n861 VSUBS 0.07fF $ **FLOATING
C972 S.n862 VSUBS 0.12fF $ **FLOATING
C973 S.n863 VSUBS 0.18fF $ **FLOATING
C974 S.n864 VSUBS 1.86fF $ **FLOATING
C975 S.n865 VSUBS 0.12fF $ **FLOATING
C976 S.t473 VSUBS 0.02fF
C977 S.n866 VSUBS 0.14fF $ **FLOATING
C978 S.t757 VSUBS 0.02fF
C979 S.n868 VSUBS 0.24fF $ **FLOATING
C980 S.n869 VSUBS 0.35fF $ **FLOATING
C981 S.n870 VSUBS 0.60fF $ **FLOATING
C982 S.n871 VSUBS 0.41fF $ **FLOATING
C983 S.n872 VSUBS 0.20fF $ **FLOATING
C984 S.n873 VSUBS 0.16fF $ **FLOATING
C985 S.n874 VSUBS 0.28fF $ **FLOATING
C986 S.n875 VSUBS 0.21fF $ **FLOATING
C987 S.n876 VSUBS 0.78fF $ **FLOATING
C988 S.n877 VSUBS 0.31fF $ **FLOATING
C989 S.n878 VSUBS 0.22fF $ **FLOATING
C990 S.n879 VSUBS 0.38fF $ **FLOATING
C991 S.n880 VSUBS 3.57fF $ **FLOATING
C992 S.t750 VSUBS 0.02fF
C993 S.n881 VSUBS 0.24fF $ **FLOATING
C994 S.n882 VSUBS 0.90fF $ **FLOATING
C995 S.n883 VSUBS 0.05fF $ **FLOATING
C996 S.t854 VSUBS 0.02fF
C997 S.n884 VSUBS 0.12fF $ **FLOATING
C998 S.n885 VSUBS 0.14fF $ **FLOATING
C999 S.n887 VSUBS 0.25fF $ **FLOATING
C1000 S.n888 VSUBS 0.09fF $ **FLOATING
C1001 S.n889 VSUBS 0.21fF $ **FLOATING
C1002 S.n890 VSUBS 1.27fF $ **FLOATING
C1003 S.n891 VSUBS 0.52fF $ **FLOATING
C1004 S.n892 VSUBS 1.86fF $ **FLOATING
C1005 S.n893 VSUBS 0.12fF $ **FLOATING
C1006 S.t815 VSUBS 0.02fF
C1007 S.n894 VSUBS 0.14fF $ **FLOATING
C1008 S.t1098 VSUBS 0.02fF
C1009 S.n896 VSUBS 0.24fF $ **FLOATING
C1010 S.n897 VSUBS 0.35fF $ **FLOATING
C1011 S.n898 VSUBS 0.60fF $ **FLOATING
C1012 S.n899 VSUBS 0.41fF $ **FLOATING
C1013 S.n900 VSUBS 0.20fF $ **FLOATING
C1014 S.n901 VSUBS 0.16fF $ **FLOATING
C1015 S.n902 VSUBS 0.28fF $ **FLOATING
C1016 S.n903 VSUBS 0.21fF $ **FLOATING
C1017 S.n904 VSUBS 0.30fF $ **FLOATING
C1018 S.n905 VSUBS 0.36fF $ **FLOATING
C1019 S.n906 VSUBS 0.22fF $ **FLOATING
C1020 S.n907 VSUBS 0.38fF $ **FLOATING
C1021 S.n908 VSUBS 2.39fF $ **FLOATING
C1022 S.t1089 VSUBS 0.02fF
C1023 S.n909 VSUBS 0.24fF $ **FLOATING
C1024 S.n910 VSUBS 0.90fF $ **FLOATING
C1025 S.n911 VSUBS 0.05fF $ **FLOATING
C1026 S.t77 VSUBS 0.02fF
C1027 S.n912 VSUBS 0.12fF $ **FLOATING
C1028 S.n913 VSUBS 0.14fF $ **FLOATING
C1029 S.n915 VSUBS 1.87fF $ **FLOATING
C1030 S.n916 VSUBS 2.64fF $ **FLOATING
C1031 S.t327 VSUBS 0.02fF
C1032 S.n917 VSUBS 0.24fF $ **FLOATING
C1033 S.n918 VSUBS 0.35fF $ **FLOATING
C1034 S.n919 VSUBS 0.60fF $ **FLOATING
C1035 S.n920 VSUBS 0.12fF $ **FLOATING
C1036 S.t26 VSUBS 0.02fF
C1037 S.n921 VSUBS 0.14fF $ **FLOATING
C1038 S.n923 VSUBS 0.69fF $ **FLOATING
C1039 S.n924 VSUBS 0.22fF $ **FLOATING
C1040 S.n925 VSUBS 0.25fF $ **FLOATING
C1041 S.n926 VSUBS 0.09fF $ **FLOATING
C1042 S.n927 VSUBS 0.22fF $ **FLOATING
C1043 S.n928 VSUBS 0.69fF $ **FLOATING
C1044 S.n929 VSUBS 1.14fF $ **FLOATING
C1045 S.n930 VSUBS 0.22fF $ **FLOATING
C1046 S.n931 VSUBS 0.25fF $ **FLOATING
C1047 S.n932 VSUBS 0.09fF $ **FLOATING
C1048 S.n933 VSUBS 1.86fF $ **FLOATING
C1049 S.t320 VSUBS 0.02fF
C1050 S.n934 VSUBS 0.24fF $ **FLOATING
C1051 S.n935 VSUBS 0.90fF $ **FLOATING
C1052 S.n936 VSUBS 0.05fF $ **FLOATING
C1053 S.t437 VSUBS 0.02fF
C1054 S.n937 VSUBS 0.12fF $ **FLOATING
C1055 S.n938 VSUBS 0.14fF $ **FLOATING
C1056 S.n940 VSUBS 14.09fF $ **FLOATING
C1057 S.n941 VSUBS 1.70fF $ **FLOATING
C1058 S.n942 VSUBS 3.02fF $ **FLOATING
C1059 S.t1118 VSUBS 0.02fF
C1060 S.n943 VSUBS 0.24fF $ **FLOATING
C1061 S.n944 VSUBS 0.35fF $ **FLOATING
C1062 S.n945 VSUBS 0.60fF $ **FLOATING
C1063 S.n946 VSUBS 0.12fF $ **FLOATING
C1064 S.t885 VSUBS 0.02fF
C1065 S.n947 VSUBS 0.14fF $ **FLOATING
C1066 S.n949 VSUBS 0.28fF $ **FLOATING
C1067 S.n950 VSUBS 0.74fF $ **FLOATING
C1068 S.n951 VSUBS 0.59fF $ **FLOATING
C1069 S.n952 VSUBS 0.20fF $ **FLOATING
C1070 S.n953 VSUBS 0.20fF $ **FLOATING
C1071 S.n954 VSUBS 0.06fF $ **FLOATING
C1072 S.n955 VSUBS 0.09fF $ **FLOATING
C1073 S.n956 VSUBS 0.09fF $ **FLOATING
C1074 S.n957 VSUBS 1.97fF $ **FLOATING
C1075 S.t157 VSUBS 0.02fF
C1076 S.n958 VSUBS 0.12fF $ **FLOATING
C1077 S.n959 VSUBS 0.14fF $ **FLOATING
C1078 S.t250 VSUBS 0.02fF
C1079 S.n961 VSUBS 0.24fF $ **FLOATING
C1080 S.n962 VSUBS 0.90fF $ **FLOATING
C1081 S.n963 VSUBS 0.05fF $ **FLOATING
C1082 S.n964 VSUBS 1.86fF $ **FLOATING
C1083 S.n965 VSUBS 0.12fF $ **FLOATING
C1084 S.t648 VSUBS 0.02fF
C1085 S.n966 VSUBS 0.14fF $ **FLOATING
C1086 S.t739 VSUBS 0.02fF
C1087 S.n968 VSUBS 1.20fF $ **FLOATING
C1088 S.n969 VSUBS 0.60fF $ **FLOATING
C1089 S.n970 VSUBS 0.35fF $ **FLOATING
C1090 S.n971 VSUBS 0.62fF $ **FLOATING
C1091 S.n972 VSUBS 1.14fF $ **FLOATING
C1092 S.n973 VSUBS 2.15fF $ **FLOATING
C1093 S.n974 VSUBS 0.59fF $ **FLOATING
C1094 S.n975 VSUBS 0.01fF $ **FLOATING
C1095 S.n976 VSUBS 0.96fF $ **FLOATING
C1096 S.t127 VSUBS 14.53fF
C1097 S.n977 VSUBS 14.40fF $ **FLOATING
C1098 S.n979 VSUBS 0.37fF $ **FLOATING
C1099 S.n980 VSUBS 0.23fF $ **FLOATING
C1100 S.n981 VSUBS 2.87fF $ **FLOATING
C1101 S.n982 VSUBS 2.43fF $ **FLOATING
C1102 S.n983 VSUBS 1.94fF $ **FLOATING
C1103 S.n984 VSUBS 3.89fF $ **FLOATING
C1104 S.n985 VSUBS 0.25fF $ **FLOATING
C1105 S.n986 VSUBS 0.01fF $ **FLOATING
C1106 S.t386 VSUBS 0.02fF
C1107 S.n987 VSUBS 0.25fF $ **FLOATING
C1108 S.t393 VSUBS 0.02fF
C1109 S.n988 VSUBS 0.94fF $ **FLOATING
C1110 S.n989 VSUBS 0.70fF $ **FLOATING
C1111 S.n990 VSUBS 0.77fF $ **FLOATING
C1112 S.n991 VSUBS 1.91fF $ **FLOATING
C1113 S.n992 VSUBS 1.86fF $ **FLOATING
C1114 S.n993 VSUBS 0.12fF $ **FLOATING
C1115 S.t784 VSUBS 0.02fF
C1116 S.n994 VSUBS 0.14fF $ **FLOATING
C1117 S.t1074 VSUBS 0.02fF
C1118 S.n996 VSUBS 0.24fF $ **FLOATING
C1119 S.n997 VSUBS 0.35fF $ **FLOATING
C1120 S.n998 VSUBS 0.60fF $ **FLOATING
C1121 S.n999 VSUBS 1.50fF $ **FLOATING
C1122 S.n1000 VSUBS 2.96fF $ **FLOATING
C1123 S.t734 VSUBS 0.02fF
C1124 S.n1001 VSUBS 0.24fF $ **FLOATING
C1125 S.n1002 VSUBS 0.90fF $ **FLOATING
C1126 S.n1003 VSUBS 0.05fF $ **FLOATING
C1127 S.t1104 VSUBS 0.02fF
C1128 S.n1004 VSUBS 0.12fF $ **FLOATING
C1129 S.n1005 VSUBS 0.14fF $ **FLOATING
C1130 S.n1007 VSUBS 1.87fF $ **FLOATING
C1131 S.n1008 VSUBS 1.86fF $ **FLOATING
C1132 S.t963 VSUBS 0.02fF
C1133 S.n1009 VSUBS 0.24fF $ **FLOATING
C1134 S.n1010 VSUBS 0.35fF $ **FLOATING
C1135 S.n1011 VSUBS 0.60fF $ **FLOATING
C1136 S.n1012 VSUBS 0.12fF $ **FLOATING
C1137 S.t602 VSUBS 0.02fF
C1138 S.n1013 VSUBS 0.14fF $ **FLOATING
C1139 S.n1015 VSUBS 1.14fF $ **FLOATING
C1140 S.n1016 VSUBS 0.22fF $ **FLOATING
C1141 S.n1017 VSUBS 0.25fF $ **FLOATING
C1142 S.n1018 VSUBS 0.09fF $ **FLOATING
C1143 S.n1019 VSUBS 1.86fF $ **FLOATING
C1144 S.t613 VSUBS 0.02fF
C1145 S.n1020 VSUBS 0.24fF $ **FLOATING
C1146 S.n1021 VSUBS 0.90fF $ **FLOATING
C1147 S.n1022 VSUBS 0.05fF $ **FLOATING
C1148 S.t408 VSUBS 0.02fF
C1149 S.n1023 VSUBS 0.12fF $ **FLOATING
C1150 S.n1024 VSUBS 0.14fF $ **FLOATING
C1151 S.n1026 VSUBS 0.77fF $ **FLOATING
C1152 S.n1027 VSUBS 1.92fF $ **FLOATING
C1153 S.n1028 VSUBS 1.86fF $ **FLOATING
C1154 S.n1029 VSUBS 0.12fF $ **FLOATING
C1155 S.t950 VSUBS 0.02fF
C1156 S.n1030 VSUBS 0.14fF $ **FLOATING
C1157 S.t204 VSUBS 0.02fF
C1158 S.n1032 VSUBS 0.24fF $ **FLOATING
C1159 S.n1033 VSUBS 0.35fF $ **FLOATING
C1160 S.n1034 VSUBS 0.60fF $ **FLOATING
C1161 S.n1035 VSUBS 1.82fF $ **FLOATING
C1162 S.n1036 VSUBS 2.96fF $ **FLOATING
C1163 S.t960 VSUBS 0.02fF
C1164 S.n1037 VSUBS 0.24fF $ **FLOATING
C1165 S.n1038 VSUBS 0.90fF $ **FLOATING
C1166 S.n1039 VSUBS 0.05fF $ **FLOATING
C1167 S.t221 VSUBS 0.02fF
C1168 S.n1040 VSUBS 0.12fF $ **FLOATING
C1169 S.n1041 VSUBS 0.14fF $ **FLOATING
C1170 S.n1043 VSUBS 1.87fF $ **FLOATING
C1171 S.n1044 VSUBS 1.86fF $ **FLOATING
C1172 S.t550 VSUBS 0.02fF
C1173 S.n1045 VSUBS 0.24fF $ **FLOATING
C1174 S.n1046 VSUBS 0.35fF $ **FLOATING
C1175 S.n1047 VSUBS 0.60fF $ **FLOATING
C1176 S.n1048 VSUBS 0.12fF $ **FLOATING
C1177 S.t189 VSUBS 0.02fF
C1178 S.n1049 VSUBS 0.14fF $ **FLOATING
C1179 S.n1051 VSUBS 1.14fF $ **FLOATING
C1180 S.n1052 VSUBS 0.22fF $ **FLOATING
C1181 S.n1053 VSUBS 0.25fF $ **FLOATING
C1182 S.n1054 VSUBS 0.09fF $ **FLOATING
C1183 S.n1055 VSUBS 1.86fF $ **FLOATING
C1184 S.t200 VSUBS 0.02fF
C1185 S.n1056 VSUBS 0.24fF $ **FLOATING
C1186 S.n1057 VSUBS 0.90fF $ **FLOATING
C1187 S.n1058 VSUBS 0.05fF $ **FLOATING
C1188 S.t570 VSUBS 0.02fF
C1189 S.n1059 VSUBS 0.12fF $ **FLOATING
C1190 S.n1060 VSUBS 0.14fF $ **FLOATING
C1191 S.n1062 VSUBS 0.77fF $ **FLOATING
C1192 S.n1063 VSUBS 1.92fF $ **FLOATING
C1193 S.n1064 VSUBS 1.86fF $ **FLOATING
C1194 S.n1065 VSUBS 0.12fF $ **FLOATING
C1195 S.t543 VSUBS 0.02fF
C1196 S.n1066 VSUBS 0.14fF $ **FLOATING
C1197 S.t895 VSUBS 0.02fF
C1198 S.n1068 VSUBS 0.24fF $ **FLOATING
C1199 S.n1069 VSUBS 0.35fF $ **FLOATING
C1200 S.n1070 VSUBS 0.60fF $ **FLOATING
C1201 S.n1071 VSUBS 0.06fF $ **FLOATING
C1202 S.n1072 VSUBS 0.89fF $ **FLOATING
C1203 S.n1073 VSUBS 1.09fF $ **FLOATING
C1204 S.n1074 VSUBS 2.94fF $ **FLOATING
C1205 S.t546 VSUBS 0.02fF
C1206 S.n1075 VSUBS 0.24fF $ **FLOATING
C1207 S.n1076 VSUBS 0.90fF $ **FLOATING
C1208 S.n1077 VSUBS 0.05fF $ **FLOATING
C1209 S.t917 VSUBS 0.02fF
C1210 S.n1078 VSUBS 0.12fF $ **FLOATING
C1211 S.n1079 VSUBS 0.14fF $ **FLOATING
C1212 S.n1081 VSUBS 0.25fF $ **FLOATING
C1213 S.n1082 VSUBS 0.09fF $ **FLOATING
C1214 S.n1083 VSUBS 1.14fF $ **FLOATING
C1215 S.n1084 VSUBS 0.22fF $ **FLOATING
C1216 S.n1085 VSUBS 1.87fF $ **FLOATING
C1217 S.n1086 VSUBS 0.12fF $ **FLOATING
C1218 S.t937 VSUBS 0.02fF
C1219 S.n1087 VSUBS 0.14fF $ **FLOATING
C1220 S.t128 VSUBS 0.02fF
C1221 S.n1089 VSUBS 0.24fF $ **FLOATING
C1222 S.n1090 VSUBS 0.35fF $ **FLOATING
C1223 S.n1091 VSUBS 0.60fF $ **FLOATING
C1224 S.n1092 VSUBS 1.09fF $ **FLOATING
C1225 S.n1093 VSUBS 0.67fF $ **FLOATING
C1226 S.n1094 VSUBS 0.54fF $ **FLOATING
C1227 S.n1095 VSUBS 0.31fF $ **FLOATING
C1228 S.n1096 VSUBS 1.81fF $ **FLOATING
C1229 S.t893 VSUBS 0.02fF
C1230 S.n1097 VSUBS 0.24fF $ **FLOATING
C1231 S.n1098 VSUBS 0.90fF $ **FLOATING
C1232 S.n1099 VSUBS 0.05fF $ **FLOATING
C1233 S.t159 VSUBS 0.02fF
C1234 S.n1100 VSUBS 0.12fF $ **FLOATING
C1235 S.n1101 VSUBS 0.14fF $ **FLOATING
C1236 S.n1103 VSUBS 1.86fF $ **FLOATING
C1237 S.n1104 VSUBS 0.47fF $ **FLOATING
C1238 S.n1105 VSUBS 0.09fF $ **FLOATING
C1239 S.n1106 VSUBS 0.32fF $ **FLOATING
C1240 S.n1107 VSUBS 0.30fF $ **FLOATING
C1241 S.n1108 VSUBS 0.76fF $ **FLOATING
C1242 S.n1109 VSUBS 0.58fF $ **FLOATING
C1243 S.t628 VSUBS 0.02fF
C1244 S.n1110 VSUBS 0.24fF $ **FLOATING
C1245 S.n1111 VSUBS 0.35fF $ **FLOATING
C1246 S.n1112 VSUBS 0.60fF $ **FLOATING
C1247 S.n1113 VSUBS 0.12fF $ **FLOATING
C1248 S.t727 VSUBS 0.02fF
C1249 S.n1114 VSUBS 0.14fF $ **FLOATING
C1250 S.n1116 VSUBS 2.58fF $ **FLOATING
C1251 S.n1117 VSUBS 2.13fF $ **FLOATING
C1252 S.t1138 VSUBS 0.02fF
C1253 S.n1118 VSUBS 0.24fF $ **FLOATING
C1254 S.n1119 VSUBS 0.90fF $ **FLOATING
C1255 S.n1120 VSUBS 0.05fF $ **FLOATING
C1256 S.t1109 VSUBS 0.02fF
C1257 S.n1121 VSUBS 0.12fF $ **FLOATING
C1258 S.n1122 VSUBS 0.14fF $ **FLOATING
C1259 S.n1124 VSUBS 1.86fF $ **FLOATING
C1260 S.n1125 VSUBS 0.47fF $ **FLOATING
C1261 S.n1126 VSUBS 0.35fF $ **FLOATING
C1262 S.n1127 VSUBS 0.30fF $ **FLOATING
C1263 S.n1128 VSUBS 1.26fF $ **FLOATING
C1264 S.t978 VSUBS 0.02fF
C1265 S.n1129 VSUBS 0.24fF $ **FLOATING
C1266 S.n1130 VSUBS 0.35fF $ **FLOATING
C1267 S.n1131 VSUBS 0.60fF $ **FLOATING
C1268 S.n1132 VSUBS 0.12fF $ **FLOATING
C1269 S.t1061 VSUBS 0.02fF
C1270 S.n1133 VSUBS 0.14fF $ **FLOATING
C1271 S.n1135 VSUBS 0.77fF $ **FLOATING
C1272 S.n1136 VSUBS 2.27fF $ **FLOATING
C1273 S.n1137 VSUBS 2.00fF $ **FLOATING
C1274 S.t376 VSUBS 0.02fF
C1275 S.n1138 VSUBS 0.24fF $ **FLOATING
C1276 S.n1139 VSUBS 0.90fF $ **FLOATING
C1277 S.n1140 VSUBS 0.05fF $ **FLOATING
C1278 S.t342 VSUBS 0.02fF
C1279 S.n1141 VSUBS 0.12fF $ **FLOATING
C1280 S.n1142 VSUBS 0.14fF $ **FLOATING
C1281 S.n1144 VSUBS 1.87fF $ **FLOATING
C1282 S.n1145 VSUBS 2.65fF $ **FLOATING
C1283 S.t217 VSUBS 0.02fF
C1284 S.n1146 VSUBS 0.24fF $ **FLOATING
C1285 S.n1147 VSUBS 0.35fF $ **FLOATING
C1286 S.n1148 VSUBS 0.60fF $ **FLOATING
C1287 S.n1149 VSUBS 0.12fF $ **FLOATING
C1288 S.t302 VSUBS 0.02fF
C1289 S.n1150 VSUBS 0.14fF $ **FLOATING
C1290 S.n1152 VSUBS 1.14fF $ **FLOATING
C1291 S.n1153 VSUBS 0.22fF $ **FLOATING
C1292 S.n1154 VSUBS 0.25fF $ **FLOATING
C1293 S.n1155 VSUBS 0.09fF $ **FLOATING
C1294 S.n1156 VSUBS 1.86fF $ **FLOATING
C1295 S.t714 VSUBS 0.02fF
C1296 S.n1157 VSUBS 0.24fF $ **FLOATING
C1297 S.n1158 VSUBS 0.90fF $ **FLOATING
C1298 S.n1159 VSUBS 0.05fF $ **FLOATING
C1299 S.t683 VSUBS 0.02fF
C1300 S.n1160 VSUBS 0.12fF $ **FLOATING
C1301 S.n1161 VSUBS 0.14fF $ **FLOATING
C1302 S.n1163 VSUBS 14.09fF $ **FLOATING
C1303 S.n1164 VSUBS 2.69fF $ **FLOATING
C1304 S.n1165 VSUBS 1.57fF $ **FLOATING
C1305 S.n1166 VSUBS 0.12fF $ **FLOATING
C1306 S.t152 VSUBS 0.02fF
C1307 S.n1167 VSUBS 0.14fF $ **FLOATING
C1308 S.t697 VSUBS 0.02fF
C1309 S.n1169 VSUBS 0.24fF $ **FLOATING
C1310 S.n1170 VSUBS 0.35fF $ **FLOATING
C1311 S.n1171 VSUBS 0.60fF $ **FLOATING
C1312 S.n1172 VSUBS 2.34fF $ **FLOATING
C1313 S.n1173 VSUBS 2.27fF $ **FLOATING
C1314 S.t264 VSUBS 0.02fF
C1315 S.n1174 VSUBS 0.12fF $ **FLOATING
C1316 S.n1175 VSUBS 0.14fF $ **FLOATING
C1317 S.t506 VSUBS 0.02fF
C1318 S.n1177 VSUBS 0.24fF $ **FLOATING
C1319 S.n1178 VSUBS 0.90fF $ **FLOATING
C1320 S.n1179 VSUBS 0.05fF $ **FLOATING
C1321 S.t151 VSUBS 32.33fF
C1322 S.t1027 VSUBS 0.02fF
C1323 S.n1180 VSUBS 0.12fF $ **FLOATING
C1324 S.n1181 VSUBS 0.14fF $ **FLOATING
C1325 S.t1051 VSUBS 0.02fF
C1326 S.n1183 VSUBS 0.24fF $ **FLOATING
C1327 S.n1184 VSUBS 0.90fF $ **FLOATING
C1328 S.n1185 VSUBS 0.05fF $ **FLOATING
C1329 S.t568 VSUBS 0.02fF
C1330 S.n1186 VSUBS 0.24fF $ **FLOATING
C1331 S.n1187 VSUBS 0.35fF $ **FLOATING
C1332 S.n1188 VSUBS 0.60fF $ **FLOATING
C1333 S.n1189 VSUBS 0.31fF $ **FLOATING
C1334 S.n1190 VSUBS 1.53fF $ **FLOATING
C1335 S.n1191 VSUBS 0.15fF $ **FLOATING
C1336 S.n1192 VSUBS 4.92fF $ **FLOATING
C1337 S.n1193 VSUBS 1.86fF $ **FLOATING
C1338 S.n1194 VSUBS 0.12fF $ **FLOATING
C1339 S.t403 VSUBS 0.02fF
C1340 S.n1195 VSUBS 0.14fF $ **FLOATING
C1341 S.t669 VSUBS 0.02fF
C1342 S.n1197 VSUBS 0.24fF $ **FLOATING
C1343 S.n1198 VSUBS 0.35fF $ **FLOATING
C1344 S.n1199 VSUBS 0.60fF $ **FLOATING
C1345 S.n1200 VSUBS 0.70fF $ **FLOATING
C1346 S.n1201 VSUBS 1.26fF $ **FLOATING
C1347 S.n1202 VSUBS 5.90fF $ **FLOATING
C1348 S.t779 VSUBS 0.02fF
C1349 S.n1203 VSUBS 0.12fF $ **FLOATING
C1350 S.n1204 VSUBS 0.14fF $ **FLOATING
C1351 S.t664 VSUBS 0.02fF
C1352 S.n1206 VSUBS 0.24fF $ **FLOATING
C1353 S.n1207 VSUBS 0.90fF $ **FLOATING
C1354 S.n1208 VSUBS 0.05fF $ **FLOATING
C1355 S.t25 VSUBS 31.95fF
C1356 S.t644 VSUBS 0.02fF
C1357 S.n1209 VSUBS 0.01fF $ **FLOATING
C1358 S.n1210 VSUBS 0.25fF $ **FLOATING
C1359 S.t139 VSUBS 0.02fF
C1360 S.n1212 VSUBS 1.18fF $ **FLOATING
C1361 S.n1213 VSUBS 0.05fF $ **FLOATING
C1362 S.t990 VSUBS 0.02fF
C1363 S.n1214 VSUBS 0.63fF $ **FLOATING
C1364 S.n1215 VSUBS 0.60fF $ **FLOATING
C1365 S.n1216 VSUBS 0.59fF $ **FLOATING
C1366 S.n1217 VSUBS 0.21fF $ **FLOATING
C1367 S.n1218 VSUBS 0.59fF $ **FLOATING
C1368 S.n1219 VSUBS 2.55fF $ **FLOATING
C1369 S.n1220 VSUBS 0.28fF $ **FLOATING
C1370 S.t166 VSUBS 14.53fF
C1371 S.n1221 VSUBS 15.80fF $ **FLOATING
C1372 S.n1222 VSUBS 0.76fF $ **FLOATING
C1373 S.n1223 VSUBS 0.27fF $ **FLOATING
C1374 S.n1224 VSUBS 3.96fF $ **FLOATING
C1375 S.n1225 VSUBS 1.49fF $ **FLOATING
C1376 S.n1226 VSUBS 0.35fF $ **FLOATING
C1377 S.n1227 VSUBS 1.28fF $ **FLOATING
C1378 S.n1228 VSUBS 0.15fF $ **FLOATING
C1379 S.n1229 VSUBS 1.64fF $ **FLOATING
C1380 S.n1230 VSUBS 2.61fF $ **FLOATING
C1381 S.n1231 VSUBS 0.24fF $ **FLOATING
C1382 S.n1232 VSUBS 1.48fF $ **FLOATING
C1383 S.n1233 VSUBS 1.29fF $ **FLOATING
C1384 S.n1234 VSUBS 0.27fF $ **FLOATING
C1385 S.n1235 VSUBS 1.87fF $ **FLOATING
C1386 S.n1236 VSUBS 0.06fF $ **FLOATING
C1387 S.n1237 VSUBS 0.03fF $ **FLOATING
C1388 S.n1238 VSUBS 0.03fF $ **FLOATING
C1389 S.n1239 VSUBS 0.98fF $ **FLOATING
C1390 S.n1240 VSUBS 0.02fF $ **FLOATING
C1391 S.n1241 VSUBS 0.01fF $ **FLOATING
C1392 S.n1242 VSUBS 0.02fF $ **FLOATING
C1393 S.n1243 VSUBS 0.08fF $ **FLOATING
C1394 S.n1244 VSUBS 0.36fF $ **FLOATING
C1395 S.n1245 VSUBS 1.83fF $ **FLOATING
C1396 S.t621 VSUBS 0.02fF
C1397 S.n1246 VSUBS 0.24fF $ **FLOATING
C1398 S.n1247 VSUBS 0.35fF $ **FLOATING
C1399 S.n1248 VSUBS 0.60fF $ **FLOATING
C1400 S.n1249 VSUBS 0.12fF $ **FLOATING
C1401 S.t266 VSUBS 0.02fF
C1402 S.n1250 VSUBS 0.14fF $ **FLOATING
C1403 S.n1252 VSUBS 0.69fF $ **FLOATING
C1404 S.n1253 VSUBS 0.22fF $ **FLOATING
C1405 S.n1254 VSUBS 0.22fF $ **FLOATING
C1406 S.n1255 VSUBS 0.69fF $ **FLOATING
C1407 S.n1256 VSUBS 1.14fF $ **FLOATING
C1408 S.n1257 VSUBS 0.22fF $ **FLOATING
C1409 S.n1258 VSUBS 0.25fF $ **FLOATING
C1410 S.n1259 VSUBS 0.09fF $ **FLOATING
C1411 S.n1260 VSUBS 1.86fF $ **FLOATING
C1412 S.t760 VSUBS 0.02fF
C1413 S.n1261 VSUBS 0.24fF $ **FLOATING
C1414 S.n1262 VSUBS 0.90fF $ **FLOATING
C1415 S.n1263 VSUBS 0.05fF $ **FLOATING
C1416 S.t646 VSUBS 0.02fF
C1417 S.n1264 VSUBS 0.12fF $ **FLOATING
C1418 S.n1265 VSUBS 0.14fF $ **FLOATING
C1419 S.n1267 VSUBS 0.25fF $ **FLOATING
C1420 S.n1268 VSUBS 0.09fF $ **FLOATING
C1421 S.n1269 VSUBS 0.21fF $ **FLOATING
C1422 S.n1270 VSUBS 0.91fF $ **FLOATING
C1423 S.n1271 VSUBS 0.44fF $ **FLOATING
C1424 S.n1272 VSUBS 1.86fF $ **FLOATING
C1425 S.n1273 VSUBS 0.12fF $ **FLOATING
C1426 S.t97 VSUBS 0.02fF
C1427 S.n1274 VSUBS 0.14fF $ **FLOATING
C1428 S.t469 VSUBS 0.02fF
C1429 S.n1276 VSUBS 0.24fF $ **FLOATING
C1430 S.n1277 VSUBS 0.35fF $ **FLOATING
C1431 S.n1278 VSUBS 0.60fF $ **FLOATING
C1432 S.n1279 VSUBS 0.02fF $ **FLOATING
C1433 S.n1280 VSUBS 0.01fF $ **FLOATING
C1434 S.n1281 VSUBS 0.02fF $ **FLOATING
C1435 S.n1282 VSUBS 0.08fF $ **FLOATING
C1436 S.n1283 VSUBS 0.06fF $ **FLOATING
C1437 S.n1284 VSUBS 0.03fF $ **FLOATING
C1438 S.n1285 VSUBS 0.03fF $ **FLOATING
C1439 S.n1286 VSUBS 0.99fF $ **FLOATING
C1440 S.n1287 VSUBS 0.35fF $ **FLOATING
C1441 S.n1288 VSUBS 1.85fF $ **FLOATING
C1442 S.n1289 VSUBS 1.97fF $ **FLOATING
C1443 S.t584 VSUBS 0.02fF
C1444 S.n1290 VSUBS 0.24fF $ **FLOATING
C1445 S.n1291 VSUBS 0.90fF $ **FLOATING
C1446 S.n1292 VSUBS 0.05fF $ **FLOATING
C1447 S.t495 VSUBS 0.02fF
C1448 S.n1293 VSUBS 0.12fF $ **FLOATING
C1449 S.n1294 VSUBS 0.14fF $ **FLOATING
C1450 S.n1296 VSUBS 1.87fF $ **FLOATING
C1451 S.n1297 VSUBS 0.06fF $ **FLOATING
C1452 S.n1298 VSUBS 0.03fF $ **FLOATING
C1453 S.n1299 VSUBS 0.03fF $ **FLOATING
C1454 S.n1300 VSUBS 0.98fF $ **FLOATING
C1455 S.n1301 VSUBS 0.02fF $ **FLOATING
C1456 S.n1302 VSUBS 0.01fF $ **FLOATING
C1457 S.n1303 VSUBS 0.02fF $ **FLOATING
C1458 S.n1304 VSUBS 0.08fF $ **FLOATING
C1459 S.n1305 VSUBS 0.36fF $ **FLOATING
C1460 S.n1306 VSUBS 1.83fF $ **FLOATING
C1461 S.t810 VSUBS 0.02fF
C1462 S.n1307 VSUBS 0.24fF $ **FLOATING
C1463 S.n1308 VSUBS 0.35fF $ **FLOATING
C1464 S.n1309 VSUBS 0.60fF $ **FLOATING
C1465 S.n1310 VSUBS 0.12fF $ **FLOATING
C1466 S.t457 VSUBS 0.02fF
C1467 S.n1311 VSUBS 0.14fF $ **FLOATING
C1468 S.n1313 VSUBS 0.69fF $ **FLOATING
C1469 S.n1314 VSUBS 0.22fF $ **FLOATING
C1470 S.n1315 VSUBS 0.22fF $ **FLOATING
C1471 S.n1316 VSUBS 0.69fF $ **FLOATING
C1472 S.n1317 VSUBS 1.14fF $ **FLOATING
C1473 S.n1318 VSUBS 0.22fF $ **FLOATING
C1474 S.n1319 VSUBS 0.25fF $ **FLOATING
C1475 S.n1320 VSUBS 0.09fF $ **FLOATING
C1476 S.n1321 VSUBS 1.86fF $ **FLOATING
C1477 S.t930 VSUBS 0.02fF
C1478 S.n1322 VSUBS 0.24fF $ **FLOATING
C1479 S.n1323 VSUBS 0.90fF $ **FLOATING
C1480 S.n1324 VSUBS 0.05fF $ **FLOATING
C1481 S.t835 VSUBS 0.02fF
C1482 S.n1325 VSUBS 0.12fF $ **FLOATING
C1483 S.n1326 VSUBS 0.14fF $ **FLOATING
C1484 S.n1328 VSUBS 0.25fF $ **FLOATING
C1485 S.n1329 VSUBS 0.09fF $ **FLOATING
C1486 S.n1330 VSUBS 0.21fF $ **FLOATING
C1487 S.n1331 VSUBS 0.91fF $ **FLOATING
C1488 S.n1332 VSUBS 0.44fF $ **FLOATING
C1489 S.n1333 VSUBS 1.86fF $ **FLOATING
C1490 S.n1334 VSUBS 0.12fF $ **FLOATING
C1491 S.t795 VSUBS 0.02fF
C1492 S.n1335 VSUBS 0.14fF $ **FLOATING
C1493 S.t17 VSUBS 0.02fF
C1494 S.n1337 VSUBS 0.24fF $ **FLOATING
C1495 S.n1338 VSUBS 0.35fF $ **FLOATING
C1496 S.n1339 VSUBS 0.60fF $ **FLOATING
C1497 S.n1340 VSUBS 0.02fF $ **FLOATING
C1498 S.n1341 VSUBS 0.01fF $ **FLOATING
C1499 S.n1342 VSUBS 0.02fF $ **FLOATING
C1500 S.n1343 VSUBS 0.08fF $ **FLOATING
C1501 S.n1344 VSUBS 0.06fF $ **FLOATING
C1502 S.n1345 VSUBS 0.03fF $ **FLOATING
C1503 S.n1346 VSUBS 0.03fF $ **FLOATING
C1504 S.n1347 VSUBS 0.99fF $ **FLOATING
C1505 S.n1348 VSUBS 0.35fF $ **FLOATING
C1506 S.n1349 VSUBS 1.81fF $ **FLOATING
C1507 S.n1350 VSUBS 1.97fF $ **FLOATING
C1508 S.t171 VSUBS 0.02fF
C1509 S.n1351 VSUBS 0.24fF $ **FLOATING
C1510 S.n1352 VSUBS 0.90fF $ **FLOATING
C1511 S.n1353 VSUBS 0.05fF $ **FLOATING
C1512 S.t56 VSUBS 0.02fF
C1513 S.n1354 VSUBS 0.12fF $ **FLOATING
C1514 S.n1355 VSUBS 0.14fF $ **FLOATING
C1515 S.n1357 VSUBS 1.87fF $ **FLOATING
C1516 S.n1358 VSUBS 0.63fF $ **FLOATING
C1517 S.n1359 VSUBS 0.07fF $ **FLOATING
C1518 S.n1360 VSUBS 0.04fF $ **FLOATING
C1519 S.n1361 VSUBS 0.05fF $ **FLOATING
C1520 S.n1362 VSUBS 0.86fF $ **FLOATING
C1521 S.n1363 VSUBS 0.01fF $ **FLOATING
C1522 S.n1364 VSUBS 0.01fF $ **FLOATING
C1523 S.n1365 VSUBS 0.01fF $ **FLOATING
C1524 S.n1366 VSUBS 0.07fF $ **FLOATING
C1525 S.n1367 VSUBS 0.68fF $ **FLOATING
C1526 S.n1368 VSUBS 0.13fF $ **FLOATING
C1527 S.t392 VSUBS 0.02fF
C1528 S.n1369 VSUBS 0.24fF $ **FLOATING
C1529 S.n1370 VSUBS 0.35fF $ **FLOATING
C1530 S.n1371 VSUBS 0.60fF $ **FLOATING
C1531 S.n1372 VSUBS 0.12fF $ **FLOATING
C1532 S.t1141 VSUBS 0.02fF
C1533 S.n1373 VSUBS 0.14fF $ **FLOATING
C1534 S.n1375 VSUBS 0.69fF $ **FLOATING
C1535 S.n1376 VSUBS 0.22fF $ **FLOATING
C1536 S.n1377 VSUBS 0.22fF $ **FLOATING
C1537 S.n1378 VSUBS 0.69fF $ **FLOATING
C1538 S.n1379 VSUBS 1.14fF $ **FLOATING
C1539 S.n1380 VSUBS 0.22fF $ **FLOATING
C1540 S.n1381 VSUBS 0.25fF $ **FLOATING
C1541 S.n1382 VSUBS 0.09fF $ **FLOATING
C1542 S.n1383 VSUBS 2.29fF $ **FLOATING
C1543 S.t520 VSUBS 0.02fF
C1544 S.n1384 VSUBS 0.24fF $ **FLOATING
C1545 S.n1385 VSUBS 0.90fF $ **FLOATING
C1546 S.n1386 VSUBS 0.05fF $ **FLOATING
C1547 S.t422 VSUBS 0.02fF
C1548 S.n1387 VSUBS 0.12fF $ **FLOATING
C1549 S.n1388 VSUBS 0.14fF $ **FLOATING
C1550 S.n1390 VSUBS 1.86fF $ **FLOATING
C1551 S.n1391 VSUBS 0.45fF $ **FLOATING
C1552 S.n1392 VSUBS 0.22fF $ **FLOATING
C1553 S.n1393 VSUBS 0.38fF $ **FLOATING
C1554 S.n1394 VSUBS 0.16fF $ **FLOATING
C1555 S.n1395 VSUBS 0.28fF $ **FLOATING
C1556 S.n1396 VSUBS 0.21fF $ **FLOATING
C1557 S.n1397 VSUBS 0.30fF $ **FLOATING
C1558 S.n1398 VSUBS 0.41fF $ **FLOATING
C1559 S.n1399 VSUBS 0.20fF $ **FLOATING
C1560 S.t638 VSUBS 0.02fF
C1561 S.n1400 VSUBS 0.24fF $ **FLOATING
C1562 S.n1401 VSUBS 0.35fF $ **FLOATING
C1563 S.n1402 VSUBS 0.60fF $ **FLOATING
C1564 S.n1403 VSUBS 0.12fF $ **FLOATING
C1565 S.t741 VSUBS 0.02fF
C1566 S.n1404 VSUBS 0.14fF $ **FLOATING
C1567 S.n1406 VSUBS 0.04fF $ **FLOATING
C1568 S.n1407 VSUBS 0.03fF $ **FLOATING
C1569 S.n1408 VSUBS 0.03fF $ **FLOATING
C1570 S.n1409 VSUBS 0.10fF $ **FLOATING
C1571 S.n1410 VSUBS 0.36fF $ **FLOATING
C1572 S.n1411 VSUBS 0.37fF $ **FLOATING
C1573 S.n1412 VSUBS 0.10fF $ **FLOATING
C1574 S.n1413 VSUBS 0.12fF $ **FLOATING
C1575 S.n1414 VSUBS 0.07fF $ **FLOATING
C1576 S.n1415 VSUBS 0.12fF $ **FLOATING
C1577 S.n1416 VSUBS 0.18fF $ **FLOATING
C1578 S.n1417 VSUBS 3.95fF $ **FLOATING
C1579 S.t1012 VSUBS 0.02fF
C1580 S.n1418 VSUBS 0.24fF $ **FLOATING
C1581 S.n1419 VSUBS 0.90fF $ **FLOATING
C1582 S.n1420 VSUBS 0.05fF $ **FLOATING
C1583 S.t821 VSUBS 0.02fF
C1584 S.n1421 VSUBS 0.12fF $ **FLOATING
C1585 S.n1422 VSUBS 0.14fF $ **FLOATING
C1586 S.n1424 VSUBS 0.25fF $ **FLOATING
C1587 S.n1425 VSUBS 0.09fF $ **FLOATING
C1588 S.n1426 VSUBS 0.21fF $ **FLOATING
C1589 S.n1427 VSUBS 1.27fF $ **FLOATING
C1590 S.n1428 VSUBS 0.52fF $ **FLOATING
C1591 S.n1429 VSUBS 1.86fF $ **FLOATING
C1592 S.n1430 VSUBS 0.12fF $ **FLOATING
C1593 S.t1076 VSUBS 0.02fF
C1594 S.n1431 VSUBS 0.14fF $ **FLOATING
C1595 S.t988 VSUBS 0.02fF
C1596 S.n1433 VSUBS 0.24fF $ **FLOATING
C1597 S.n1434 VSUBS 0.35fF $ **FLOATING
C1598 S.n1435 VSUBS 0.60fF $ **FLOATING
C1599 S.n1436 VSUBS 0.70fF $ **FLOATING
C1600 S.n1437 VSUBS 1.56fF $ **FLOATING
C1601 S.n1438 VSUBS 2.42fF $ **FLOATING
C1602 S.t248 VSUBS 0.02fF
C1603 S.n1439 VSUBS 0.24fF $ **FLOATING
C1604 S.n1440 VSUBS 0.90fF $ **FLOATING
C1605 S.n1441 VSUBS 0.05fF $ **FLOATING
C1606 S.t358 VSUBS 0.02fF
C1607 S.n1442 VSUBS 0.12fF $ **FLOATING
C1608 S.n1443 VSUBS 0.14fF $ **FLOATING
C1609 S.n1445 VSUBS 1.87fF $ **FLOATING
C1610 S.n1446 VSUBS 0.06fF $ **FLOATING
C1611 S.n1447 VSUBS 0.03fF $ **FLOATING
C1612 S.n1448 VSUBS 0.03fF $ **FLOATING
C1613 S.n1449 VSUBS 0.98fF $ **FLOATING
C1614 S.n1450 VSUBS 0.02fF $ **FLOATING
C1615 S.n1451 VSUBS 0.01fF $ **FLOATING
C1616 S.n1452 VSUBS 0.02fF $ **FLOATING
C1617 S.n1453 VSUBS 0.08fF $ **FLOATING
C1618 S.n1454 VSUBS 0.36fF $ **FLOATING
C1619 S.n1455 VSUBS 1.83fF $ **FLOATING
C1620 S.t228 VSUBS 0.02fF
C1621 S.n1456 VSUBS 0.24fF $ **FLOATING
C1622 S.n1457 VSUBS 0.35fF $ **FLOATING
C1623 S.n1458 VSUBS 0.60fF $ **FLOATING
C1624 S.n1459 VSUBS 0.12fF $ **FLOATING
C1625 S.t309 VSUBS 0.02fF
C1626 S.n1460 VSUBS 0.14fF $ **FLOATING
C1627 S.n1462 VSUBS 0.69fF $ **FLOATING
C1628 S.n1463 VSUBS 0.22fF $ **FLOATING
C1629 S.n1464 VSUBS 0.22fF $ **FLOATING
C1630 S.n1465 VSUBS 0.69fF $ **FLOATING
C1631 S.n1466 VSUBS 1.14fF $ **FLOATING
C1632 S.n1467 VSUBS 0.22fF $ **FLOATING
C1633 S.n1468 VSUBS 0.25fF $ **FLOATING
C1634 S.n1469 VSUBS 0.09fF $ **FLOATING
C1635 S.n1470 VSUBS 1.86fF $ **FLOATING
C1636 S.t599 VSUBS 0.02fF
C1637 S.n1471 VSUBS 0.24fF $ **FLOATING
C1638 S.n1472 VSUBS 0.90fF $ **FLOATING
C1639 S.n1473 VSUBS 0.05fF $ **FLOATING
C1640 S.t691 VSUBS 0.02fF
C1641 S.n1474 VSUBS 0.12fF $ **FLOATING
C1642 S.n1475 VSUBS 0.14fF $ **FLOATING
C1643 S.n1477 VSUBS 14.09fF $ **FLOATING
C1644 S.n1478 VSUBS 0.06fF $ **FLOATING
C1645 S.n1479 VSUBS 0.20fF $ **FLOATING
C1646 S.n1480 VSUBS 0.09fF $ **FLOATING
C1647 S.n1481 VSUBS 0.20fF $ **FLOATING
C1648 S.n1482 VSUBS 0.09fF $ **FLOATING
C1649 S.n1483 VSUBS 0.30fF $ **FLOATING
C1650 S.n1484 VSUBS 0.69fF $ **FLOATING
C1651 S.n1485 VSUBS 0.44fF $ **FLOATING
C1652 S.n1486 VSUBS 2.30fF $ **FLOATING
C1653 S.n1487 VSUBS 0.12fF $ **FLOATING
C1654 S.t973 VSUBS 0.02fF
C1655 S.n1488 VSUBS 0.14fF $ **FLOATING
C1656 S.t224 VSUBS 0.02fF
C1657 S.n1490 VSUBS 0.24fF $ **FLOATING
C1658 S.n1491 VSUBS 0.35fF $ **FLOATING
C1659 S.n1492 VSUBS 0.60fF $ **FLOATING
C1660 S.n1493 VSUBS 1.88fF $ **FLOATING
C1661 S.n1494 VSUBS 0.17fF $ **FLOATING
C1662 S.n1495 VSUBS 0.76fF $ **FLOATING
C1663 S.n1496 VSUBS 0.31fF $ **FLOATING
C1664 S.n1497 VSUBS 0.25fF $ **FLOATING
C1665 S.n1498 VSUBS 0.29fF $ **FLOATING
C1666 S.n1499 VSUBS 0.46fF $ **FLOATING
C1667 S.n1500 VSUBS 0.16fF $ **FLOATING
C1668 S.n1501 VSUBS 1.90fF $ **FLOATING
C1669 S.t245 VSUBS 0.02fF
C1670 S.n1502 VSUBS 0.12fF $ **FLOATING
C1671 S.n1503 VSUBS 0.14fF $ **FLOATING
C1672 S.t354 VSUBS 0.02fF
C1673 S.n1505 VSUBS 0.24fF $ **FLOATING
C1674 S.n1506 VSUBS 0.90fF $ **FLOATING
C1675 S.n1507 VSUBS 0.05fF $ **FLOATING
C1676 S.n1508 VSUBS 1.86fF $ **FLOATING
C1677 S.n1509 VSUBS 0.12fF $ **FLOATING
C1678 S.t668 VSUBS 0.02fF
C1679 S.n1510 VSUBS 0.14fF $ **FLOATING
C1680 S.t498 VSUBS 0.02fF
C1681 S.n1512 VSUBS 1.20fF $ **FLOATING
C1682 S.n1513 VSUBS 0.36fF $ **FLOATING
C1683 S.n1514 VSUBS 1.21fF $ **FLOATING
C1684 S.n1515 VSUBS 0.60fF $ **FLOATING
C1685 S.n1516 VSUBS 0.35fF $ **FLOATING
C1686 S.n1517 VSUBS 0.62fF $ **FLOATING
C1687 S.n1518 VSUBS 1.14fF $ **FLOATING
C1688 S.n1519 VSUBS 2.15fF $ **FLOATING
C1689 S.n1520 VSUBS 0.59fF $ **FLOATING
C1690 S.n1521 VSUBS 0.01fF $ **FLOATING
C1691 S.n1522 VSUBS 0.96fF $ **FLOATING
C1692 S.t99 VSUBS 14.53fF
C1693 S.n1523 VSUBS 14.40fF $ **FLOATING
C1694 S.n1525 VSUBS 0.37fF $ **FLOATING
C1695 S.n1526 VSUBS 0.23fF $ **FLOATING
C1696 S.n1527 VSUBS 2.76fF $ **FLOATING
C1697 S.n1528 VSUBS 2.43fF $ **FLOATING
C1698 S.n1529 VSUBS 3.96fF $ **FLOATING
C1699 S.n1530 VSUBS 0.25fF $ **FLOATING
C1700 S.n1531 VSUBS 0.01fF $ **FLOATING
C1701 S.t124 VSUBS 0.02fF
C1702 S.n1532 VSUBS 0.25fF $ **FLOATING
C1703 S.t605 VSUBS 0.02fF
C1704 S.n1533 VSUBS 0.94fF $ **FLOATING
C1705 S.n1534 VSUBS 0.70fF $ **FLOATING
C1706 S.n1535 VSUBS 1.87fF $ **FLOATING
C1707 S.n1536 VSUBS 1.86fF $ **FLOATING
C1708 S.t836 VSUBS 0.02fF
C1709 S.n1537 VSUBS 0.24fF $ **FLOATING
C1710 S.n1538 VSUBS 0.35fF $ **FLOATING
C1711 S.n1539 VSUBS 0.60fF $ **FLOATING
C1712 S.n1540 VSUBS 0.12fF $ **FLOATING
C1713 S.t537 VSUBS 0.02fF
C1714 S.n1541 VSUBS 0.14fF $ **FLOATING
C1715 S.n1543 VSUBS 1.14fF $ **FLOATING
C1716 S.n1544 VSUBS 0.22fF $ **FLOATING
C1717 S.n1545 VSUBS 0.25fF $ **FLOATING
C1718 S.n1546 VSUBS 0.09fF $ **FLOATING
C1719 S.n1547 VSUBS 1.86fF $ **FLOATING
C1720 S.t953 VSUBS 0.02fF
C1721 S.n1548 VSUBS 0.24fF $ **FLOATING
C1722 S.n1549 VSUBS 0.90fF $ **FLOATING
C1723 S.n1550 VSUBS 0.05fF $ **FLOATING
C1724 S.t859 VSUBS 0.02fF
C1725 S.n1551 VSUBS 0.12fF $ **FLOATING
C1726 S.n1552 VSUBS 0.14fF $ **FLOATING
C1727 S.n1554 VSUBS 0.77fF $ **FLOATING
C1728 S.n1555 VSUBS 1.92fF $ **FLOATING
C1729 S.n1556 VSUBS 1.86fF $ **FLOATING
C1730 S.n1557 VSUBS 0.12fF $ **FLOATING
C1731 S.t360 VSUBS 0.02fF
C1732 S.n1558 VSUBS 0.14fF $ **FLOATING
C1733 S.t713 VSUBS 0.02fF
C1734 S.n1560 VSUBS 0.24fF $ **FLOATING
C1735 S.n1561 VSUBS 0.35fF $ **FLOATING
C1736 S.n1562 VSUBS 0.60fF $ **FLOATING
C1737 S.n1563 VSUBS 1.82fF $ **FLOATING
C1738 S.n1564 VSUBS 2.96fF $ **FLOATING
C1739 S.t849 VSUBS 0.02fF
C1740 S.n1565 VSUBS 0.24fF $ **FLOATING
C1741 S.n1566 VSUBS 0.90fF $ **FLOATING
C1742 S.n1567 VSUBS 0.05fF $ **FLOATING
C1743 S.t149 VSUBS 0.02fF
C1744 S.n1568 VSUBS 0.12fF $ **FLOATING
C1745 S.n1569 VSUBS 0.14fF $ **FLOATING
C1746 S.n1571 VSUBS 1.87fF $ **FLOATING
C1747 S.n1572 VSUBS 1.86fF $ **FLOATING
C1748 S.t1050 VSUBS 0.02fF
C1749 S.n1573 VSUBS 0.24fF $ **FLOATING
C1750 S.n1574 VSUBS 0.35fF $ **FLOATING
C1751 S.n1575 VSUBS 0.60fF $ **FLOATING
C1752 S.n1576 VSUBS 0.12fF $ **FLOATING
C1753 S.t692 VSUBS 0.02fF
C1754 S.n1577 VSUBS 0.14fF $ **FLOATING
C1755 S.n1579 VSUBS 1.14fF $ **FLOATING
C1756 S.n1580 VSUBS 0.22fF $ **FLOATING
C1757 S.n1581 VSUBS 0.25fF $ **FLOATING
C1758 S.n1582 VSUBS 0.09fF $ **FLOATING
C1759 S.n1583 VSUBS 1.86fF $ **FLOATING
C1760 S.t74 VSUBS 0.02fF
C1761 S.n1584 VSUBS 0.24fF $ **FLOATING
C1762 S.n1585 VSUBS 0.90fF $ **FLOATING
C1763 S.n1586 VSUBS 0.05fF $ **FLOATING
C1764 S.t1079 VSUBS 0.02fF
C1765 S.n1587 VSUBS 0.12fF $ **FLOATING
C1766 S.n1588 VSUBS 0.14fF $ **FLOATING
C1767 S.n1590 VSUBS 0.77fF $ **FLOATING
C1768 S.n1591 VSUBS 1.92fF $ **FLOATING
C1769 S.n1592 VSUBS 1.86fF $ **FLOATING
C1770 S.n1593 VSUBS 0.12fF $ **FLOATING
C1771 S.t1037 VSUBS 0.02fF
C1772 S.n1594 VSUBS 0.14fF $ **FLOATING
C1773 S.t289 VSUBS 0.02fF
C1774 S.n1596 VSUBS 0.24fF $ **FLOATING
C1775 S.n1597 VSUBS 0.35fF $ **FLOATING
C1776 S.n1598 VSUBS 0.60fF $ **FLOATING
C1777 S.n1599 VSUBS 1.82fF $ **FLOATING
C1778 S.n1600 VSUBS 2.96fF $ **FLOATING
C1779 S.t432 VSUBS 0.02fF
C1780 S.n1601 VSUBS 0.24fF $ **FLOATING
C1781 S.n1602 VSUBS 0.90fF $ **FLOATING
C1782 S.n1603 VSUBS 0.05fF $ **FLOATING
C1783 S.t311 VSUBS 0.02fF
C1784 S.n1604 VSUBS 0.12fF $ **FLOATING
C1785 S.n1605 VSUBS 0.14fF $ **FLOATING
C1786 S.n1607 VSUBS 1.87fF $ **FLOATING
C1787 S.n1608 VSUBS 1.73fF $ **FLOATING
C1788 S.t632 VSUBS 0.02fF
C1789 S.n1609 VSUBS 0.24fF $ **FLOATING
C1790 S.n1610 VSUBS 0.35fF $ **FLOATING
C1791 S.n1611 VSUBS 0.60fF $ **FLOATING
C1792 S.n1612 VSUBS 0.12fF $ **FLOATING
C1793 S.t280 VSUBS 0.02fF
C1794 S.n1613 VSUBS 0.14fF $ **FLOATING
C1795 S.n1615 VSUBS 1.14fF $ **FLOATING
C1796 S.n1616 VSUBS 0.22fF $ **FLOATING
C1797 S.n1617 VSUBS 0.25fF $ **FLOATING
C1798 S.n1618 VSUBS 0.09fF $ **FLOATING
C1799 S.n1619 VSUBS 2.41fF $ **FLOATING
C1800 S.t772 VSUBS 0.02fF
C1801 S.n1620 VSUBS 0.24fF $ **FLOATING
C1802 S.n1621 VSUBS 0.90fF $ **FLOATING
C1803 S.n1622 VSUBS 0.05fF $ **FLOATING
C1804 S.t658 VSUBS 0.02fF
C1805 S.n1623 VSUBS 0.12fF $ **FLOATING
C1806 S.n1624 VSUBS 0.14fF $ **FLOATING
C1807 S.n1626 VSUBS 1.86fF $ **FLOATING
C1808 S.n1627 VSUBS 0.47fF $ **FLOATING
C1809 S.n1628 VSUBS 0.09fF $ **FLOATING
C1810 S.n1629 VSUBS 0.32fF $ **FLOATING
C1811 S.n1630 VSUBS 0.30fF $ **FLOATING
C1812 S.n1631 VSUBS 0.76fF $ **FLOATING
C1813 S.n1632 VSUBS 0.58fF $ **FLOATING
C1814 S.t981 VSUBS 0.02fF
C1815 S.n1633 VSUBS 0.24fF $ **FLOATING
C1816 S.n1634 VSUBS 0.35fF $ **FLOATING
C1817 S.n1635 VSUBS 0.60fF $ **FLOATING
C1818 S.n1636 VSUBS 0.12fF $ **FLOATING
C1819 S.t678 VSUBS 0.02fF
C1820 S.n1637 VSUBS 0.14fF $ **FLOATING
C1821 S.n1639 VSUBS 2.58fF $ **FLOATING
C1822 S.n1640 VSUBS 2.13fF $ **FLOATING
C1823 S.t1117 VSUBS 0.02fF
C1824 S.n1641 VSUBS 0.24fF $ **FLOATING
C1825 S.n1642 VSUBS 0.90fF $ **FLOATING
C1826 S.n1643 VSUBS 0.05fF $ **FLOATING
C1827 S.t1004 VSUBS 0.02fF
C1828 S.n1644 VSUBS 0.12fF $ **FLOATING
C1829 S.n1645 VSUBS 0.14fF $ **FLOATING
C1830 S.n1647 VSUBS 0.77fF $ **FLOATING
C1831 S.n1648 VSUBS 2.27fF $ **FLOATING
C1832 S.n1649 VSUBS 1.86fF $ **FLOATING
C1833 S.n1650 VSUBS 0.12fF $ **FLOATING
C1834 S.t1097 VSUBS 0.02fF
C1835 S.n1651 VSUBS 0.14fF $ **FLOATING
C1836 S.t998 VSUBS 0.02fF
C1837 S.n1653 VSUBS 0.24fF $ **FLOATING
C1838 S.n1654 VSUBS 0.35fF $ **FLOATING
C1839 S.n1655 VSUBS 0.60fF $ **FLOATING
C1840 S.n1656 VSUBS 1.37fF $ **FLOATING
C1841 S.n1657 VSUBS 0.70fF $ **FLOATING
C1842 S.n1658 VSUBS 1.13fF $ **FLOATING
C1843 S.n1659 VSUBS 0.35fF $ **FLOATING
C1844 S.n1660 VSUBS 2.00fF $ **FLOATING
C1845 S.t259 VSUBS 0.02fF
C1846 S.n1661 VSUBS 0.24fF $ **FLOATING
C1847 S.n1662 VSUBS 0.90fF $ **FLOATING
C1848 S.n1663 VSUBS 0.05fF $ **FLOATING
C1849 S.t374 VSUBS 0.02fF
C1850 S.n1664 VSUBS 0.12fF $ **FLOATING
C1851 S.n1665 VSUBS 0.14fF $ **FLOATING
C1852 S.n1667 VSUBS 1.87fF $ **FLOATING
C1853 S.n1668 VSUBS 1.86fF $ **FLOATING
C1854 S.t240 VSUBS 0.02fF
C1855 S.n1669 VSUBS 0.24fF $ **FLOATING
C1856 S.n1670 VSUBS 0.35fF $ **FLOATING
C1857 S.n1671 VSUBS 0.60fF $ **FLOATING
C1858 S.n1672 VSUBS 0.12fF $ **FLOATING
C1859 S.t324 VSUBS 0.02fF
C1860 S.n1673 VSUBS 0.14fF $ **FLOATING
C1861 S.n1675 VSUBS 1.14fF $ **FLOATING
C1862 S.n1676 VSUBS 0.22fF $ **FLOATING
C1863 S.n1677 VSUBS 0.25fF $ **FLOATING
C1864 S.n1678 VSUBS 0.09fF $ **FLOATING
C1865 S.n1679 VSUBS 1.86fF $ **FLOATING
C1866 S.t609 VSUBS 0.02fF
C1867 S.n1680 VSUBS 0.24fF $ **FLOATING
C1868 S.n1681 VSUBS 0.90fF $ **FLOATING
C1869 S.n1682 VSUBS 0.05fF $ **FLOATING
C1870 S.t710 VSUBS 0.02fF
C1871 S.n1683 VSUBS 0.12fF $ **FLOATING
C1872 S.n1684 VSUBS 0.14fF $ **FLOATING
C1873 S.n1686 VSUBS 14.09fF $ **FLOATING
C1874 S.n1687 VSUBS 1.86fF $ **FLOATING
C1875 S.n1688 VSUBS 2.65fF $ **FLOATING
C1876 S.t935 VSUBS 0.02fF
C1877 S.n1689 VSUBS 0.24fF $ **FLOATING
C1878 S.n1690 VSUBS 0.35fF $ **FLOATING
C1879 S.n1691 VSUBS 0.60fF $ **FLOATING
C1880 S.n1692 VSUBS 0.12fF $ **FLOATING
C1881 S.t1015 VSUBS 0.02fF
C1882 S.n1693 VSUBS 0.14fF $ **FLOATING
C1883 S.n1695 VSUBS 5.12fF $ **FLOATING
C1884 S.t287 VSUBS 0.02fF
C1885 S.n1696 VSUBS 0.12fF $ **FLOATING
C1886 S.n1697 VSUBS 0.14fF $ **FLOATING
C1887 S.t195 VSUBS 0.02fF
C1888 S.n1699 VSUBS 0.24fF $ **FLOATING
C1889 S.n1700 VSUBS 0.90fF $ **FLOATING
C1890 S.n1701 VSUBS 0.05fF $ **FLOATING
C1891 S.n1702 VSUBS 2.70fF $ **FLOATING
C1892 S.n1703 VSUBS 1.58fF $ **FLOATING
C1893 S.n1704 VSUBS 0.12fF $ **FLOATING
C1894 S.t43 VSUBS 0.02fF
C1895 S.n1705 VSUBS 0.14fF $ **FLOATING
C1896 S.t587 VSUBS 0.02fF
C1897 S.n1707 VSUBS 0.24fF $ **FLOATING
C1898 S.n1708 VSUBS 0.35fF $ **FLOATING
C1899 S.n1709 VSUBS 0.60fF $ **FLOATING
C1900 S.n1710 VSUBS 0.07fF $ **FLOATING
C1901 S.n1711 VSUBS 0.01fF $ **FLOATING
C1902 S.n1712 VSUBS 0.23fF $ **FLOATING
C1903 S.n1713 VSUBS 1.15fF $ **FLOATING
C1904 S.n1714 VSUBS 1.33fF $ **FLOATING
C1905 S.n1715 VSUBS 2.27fF $ **FLOATING
C1906 S.t631 VSUBS 0.02fF
C1907 S.n1716 VSUBS 0.12fF $ **FLOATING
C1908 S.n1717 VSUBS 0.14fF $ **FLOATING
C1909 S.t86 VSUBS 0.02fF
C1910 S.n1719 VSUBS 0.24fF $ **FLOATING
C1911 S.n1720 VSUBS 0.90fF $ **FLOATING
C1912 S.n1721 VSUBS 0.05fF $ **FLOATING
C1913 S.t42 VSUBS 32.33fF
C1914 S.t1048 VSUBS 0.02fF
C1915 S.n1722 VSUBS 0.12fF $ **FLOATING
C1916 S.n1723 VSUBS 0.14fF $ **FLOATING
C1917 S.t954 VSUBS 0.02fF
C1918 S.n1725 VSUBS 0.24fF $ **FLOATING
C1919 S.n1726 VSUBS 0.90fF $ **FLOATING
C1920 S.n1727 VSUBS 0.05fF $ **FLOATING
C1921 S.t590 VSUBS 0.02fF
C1922 S.n1728 VSUBS 0.24fF $ **FLOATING
C1923 S.n1729 VSUBS 0.35fF $ **FLOATING
C1924 S.n1730 VSUBS 0.60fF $ **FLOATING
C1925 S.n1731 VSUBS 0.31fF $ **FLOATING
C1926 S.n1732 VSUBS 1.08fF $ **FLOATING
C1927 S.n1733 VSUBS 0.15fF $ **FLOATING
C1928 S.n1734 VSUBS 2.08fF $ **FLOATING
C1929 S.n1735 VSUBS 2.91fF $ **FLOATING
C1930 S.n1736 VSUBS 1.86fF $ **FLOATING
C1931 S.n1737 VSUBS 0.12fF $ **FLOATING
C1932 S.t656 VSUBS 0.02fF
C1933 S.n1738 VSUBS 0.14fF $ **FLOATING
C1934 S.t576 VSUBS 0.02fF
C1935 S.n1740 VSUBS 0.24fF $ **FLOATING
C1936 S.n1741 VSUBS 0.35fF $ **FLOATING
C1937 S.n1742 VSUBS 0.60fF $ **FLOATING
C1938 S.n1743 VSUBS 0.91fF $ **FLOATING
C1939 S.n1744 VSUBS 0.31fF $ **FLOATING
C1940 S.n1745 VSUBS 0.91fF $ **FLOATING
C1941 S.n1746 VSUBS 1.08fF $ **FLOATING
C1942 S.n1747 VSUBS 0.15fF $ **FLOATING
C1943 S.n1748 VSUBS 4.63fF $ **FLOATING
C1944 S.t1035 VSUBS 0.02fF
C1945 S.n1749 VSUBS 0.12fF $ **FLOATING
C1946 S.n1750 VSUBS 0.14fF $ **FLOATING
C1947 S.t946 VSUBS 0.02fF
C1948 S.n1752 VSUBS 0.24fF $ **FLOATING
C1949 S.n1753 VSUBS 0.90fF $ **FLOATING
C1950 S.n1754 VSUBS 0.05fF $ **FLOATING
C1951 S.n1755 VSUBS 1.86fF $ **FLOATING
C1952 S.n1756 VSUBS 2.64fF $ **FLOATING
C1953 S.t924 VSUBS 0.02fF
C1954 S.n1757 VSUBS 0.24fF $ **FLOATING
C1955 S.n1758 VSUBS 0.35fF $ **FLOATING
C1956 S.n1759 VSUBS 0.60fF $ **FLOATING
C1957 S.n1760 VSUBS 0.12fF $ **FLOATING
C1958 S.t1003 VSUBS 0.02fF
C1959 S.n1761 VSUBS 0.14fF $ **FLOATING
C1960 S.n1763 VSUBS 5.39fF $ **FLOATING
C1961 S.t278 VSUBS 0.02fF
C1962 S.n1764 VSUBS 0.12fF $ **FLOATING
C1963 S.n1765 VSUBS 0.14fF $ **FLOATING
C1964 S.t187 VSUBS 0.02fF
C1965 S.n1767 VSUBS 0.24fF $ **FLOATING
C1966 S.n1768 VSUBS 0.90fF $ **FLOATING
C1967 S.n1769 VSUBS 0.05fF $ **FLOATING
C1968 S.t55 VSUBS 31.95fF
C1969 S.t649 VSUBS 0.02fF
C1970 S.n1770 VSUBS 0.01fF $ **FLOATING
C1971 S.n1771 VSUBS 0.25fF $ **FLOATING
C1972 S.t234 VSUBS 0.02fF
C1973 S.n1773 VSUBS 1.18fF $ **FLOATING
C1974 S.n1774 VSUBS 0.05fF $ **FLOATING
C1975 S.t111 VSUBS 0.02fF
C1976 S.n1775 VSUBS 0.63fF $ **FLOATING
C1977 S.n1776 VSUBS 0.60fF $ **FLOATING
C1978 S.n1777 VSUBS 8.88fF $ **FLOATING
C1979 S.n1778 VSUBS 8.88fF $ **FLOATING
C1980 S.n1779 VSUBS 0.59fF $ **FLOATING
C1981 S.n1780 VSUBS 0.21fF $ **FLOATING
C1982 S.n1781 VSUBS 0.59fF $ **FLOATING
C1983 S.n1782 VSUBS 2.55fF $ **FLOATING
C1984 S.n1783 VSUBS 0.28fF $ **FLOATING
C1985 S.t16 VSUBS 14.53fF
C1986 S.n1784 VSUBS 15.80fF $ **FLOATING
C1987 S.n1785 VSUBS 0.76fF $ **FLOATING
C1988 S.n1786 VSUBS 0.27fF $ **FLOATING
C1989 S.n1787 VSUBS 3.96fF $ **FLOATING
C1990 S.n1788 VSUBS 1.34fF $ **FLOATING
C1991 S.n1789 VSUBS 0.01fF $ **FLOATING
C1992 S.n1790 VSUBS 0.02fF $ **FLOATING
C1993 S.n1791 VSUBS 0.03fF $ **FLOATING
C1994 S.n1792 VSUBS 0.04fF $ **FLOATING
C1995 S.n1793 VSUBS 0.17fF $ **FLOATING
C1996 S.n1794 VSUBS 0.01fF $ **FLOATING
C1997 S.n1795 VSUBS 0.02fF $ **FLOATING
C1998 S.n1796 VSUBS 0.01fF $ **FLOATING
C1999 S.n1797 VSUBS 0.01fF $ **FLOATING
C2000 S.n1798 VSUBS 0.01fF $ **FLOATING
C2001 S.n1799 VSUBS 0.01fF $ **FLOATING
C2002 S.n1800 VSUBS 0.01fF $ **FLOATING
C2003 S.n1801 VSUBS 0.01fF $ **FLOATING
C2004 S.n1802 VSUBS 0.02fF $ **FLOATING
C2005 S.n1803 VSUBS 0.05fF $ **FLOATING
C2006 S.n1804 VSUBS 0.04fF $ **FLOATING
C2007 S.n1805 VSUBS 0.11fF $ **FLOATING
C2008 S.n1806 VSUBS 0.37fF $ **FLOATING
C2009 S.n1807 VSUBS 0.20fF $ **FLOATING
C2010 S.n1808 VSUBS 4.34fF $ **FLOATING
C2011 S.n1809 VSUBS 0.24fF $ **FLOATING
C2012 S.n1810 VSUBS 1.48fF $ **FLOATING
C2013 S.n1811 VSUBS 1.29fF $ **FLOATING
C2014 S.n1812 VSUBS 0.27fF $ **FLOATING
C2015 S.n1813 VSUBS 0.25fF $ **FLOATING
C2016 S.n1814 VSUBS 0.09fF $ **FLOATING
C2017 S.n1815 VSUBS 0.21fF $ **FLOATING
C2018 S.n1816 VSUBS 0.91fF $ **FLOATING
C2019 S.n1817 VSUBS 0.44fF $ **FLOATING
C2020 S.n1818 VSUBS 1.86fF $ **FLOATING
C2021 S.n1819 VSUBS 0.12fF $ **FLOATING
C2022 S.t1132 VSUBS 0.02fF
C2023 S.n1820 VSUBS 0.14fF $ **FLOATING
C2024 S.t385 VSUBS 0.02fF
C2025 S.n1822 VSUBS 0.24fF $ **FLOATING
C2026 S.n1823 VSUBS 0.35fF $ **FLOATING
C2027 S.n1824 VSUBS 0.60fF $ **FLOATING
C2028 S.n1825 VSUBS 0.02fF $ **FLOATING
C2029 S.n1826 VSUBS 0.01fF $ **FLOATING
C2030 S.n1827 VSUBS 0.02fF $ **FLOATING
C2031 S.n1828 VSUBS 0.08fF $ **FLOATING
C2032 S.n1829 VSUBS 0.06fF $ **FLOATING
C2033 S.n1830 VSUBS 0.03fF $ **FLOATING
C2034 S.n1831 VSUBS 0.03fF $ **FLOATING
C2035 S.n1832 VSUBS 0.99fF $ **FLOATING
C2036 S.n1833 VSUBS 0.35fF $ **FLOATING
C2037 S.n1834 VSUBS 1.85fF $ **FLOATING
C2038 S.n1835 VSUBS 1.97fF $ **FLOATING
C2039 S.t515 VSUBS 0.02fF
C2040 S.n1836 VSUBS 0.24fF $ **FLOATING
C2041 S.n1837 VSUBS 0.90fF $ **FLOATING
C2042 S.n1838 VSUBS 0.05fF $ **FLOATING
C2043 S.t414 VSUBS 0.02fF
C2044 S.n1839 VSUBS 0.12fF $ **FLOATING
C2045 S.n1840 VSUBS 0.14fF $ **FLOATING
C2046 S.n1842 VSUBS 1.87fF $ **FLOATING
C2047 S.n1843 VSUBS 0.06fF $ **FLOATING
C2048 S.n1844 VSUBS 0.03fF $ **FLOATING
C2049 S.n1845 VSUBS 0.03fF $ **FLOATING
C2050 S.n1846 VSUBS 0.98fF $ **FLOATING
C2051 S.n1847 VSUBS 0.02fF $ **FLOATING
C2052 S.n1848 VSUBS 0.01fF $ **FLOATING
C2053 S.n1849 VSUBS 0.02fF $ **FLOATING
C2054 S.n1850 VSUBS 0.08fF $ **FLOATING
C2055 S.n1851 VSUBS 0.36fF $ **FLOATING
C2056 S.n1852 VSUBS 1.83fF $ **FLOATING
C2057 S.t209 VSUBS 0.02fF
C2058 S.n1853 VSUBS 0.24fF $ **FLOATING
C2059 S.n1854 VSUBS 0.35fF $ **FLOATING
C2060 S.n1855 VSUBS 0.60fF $ **FLOATING
C2061 S.n1856 VSUBS 0.12fF $ **FLOATING
C2062 S.t956 VSUBS 0.02fF
C2063 S.n1857 VSUBS 0.14fF $ **FLOATING
C2064 S.n1859 VSUBS 0.69fF $ **FLOATING
C2065 S.n1860 VSUBS 0.22fF $ **FLOATING
C2066 S.n1861 VSUBS 0.22fF $ **FLOATING
C2067 S.n1862 VSUBS 0.69fF $ **FLOATING
C2068 S.n1863 VSUBS 1.14fF $ **FLOATING
C2069 S.n1864 VSUBS 0.22fF $ **FLOATING
C2070 S.n1865 VSUBS 0.25fF $ **FLOATING
C2071 S.n1866 VSUBS 0.09fF $ **FLOATING
C2072 S.n1867 VSUBS 1.86fF $ **FLOATING
C2073 S.t326 VSUBS 0.02fF
C2074 S.n1868 VSUBS 0.24fF $ **FLOATING
C2075 S.n1869 VSUBS 0.90fF $ **FLOATING
C2076 S.n1870 VSUBS 0.05fF $ **FLOATING
C2077 S.t227 VSUBS 0.02fF
C2078 S.n1871 VSUBS 0.12fF $ **FLOATING
C2079 S.n1872 VSUBS 0.14fF $ **FLOATING
C2080 S.n1874 VSUBS 0.25fF $ **FLOATING
C2081 S.n1875 VSUBS 0.09fF $ **FLOATING
C2082 S.n1876 VSUBS 0.21fF $ **FLOATING
C2083 S.n1877 VSUBS 0.91fF $ **FLOATING
C2084 S.n1878 VSUBS 0.44fF $ **FLOATING
C2085 S.n1879 VSUBS 1.86fF $ **FLOATING
C2086 S.n1880 VSUBS 0.12fF $ **FLOATING
C2087 S.t194 VSUBS 0.02fF
C2088 S.n1881 VSUBS 0.14fF $ **FLOATING
C2089 S.t557 VSUBS 0.02fF
C2090 S.n1883 VSUBS 0.24fF $ **FLOATING
C2091 S.n1884 VSUBS 0.35fF $ **FLOATING
C2092 S.n1885 VSUBS 0.60fF $ **FLOATING
C2093 S.n1886 VSUBS 0.02fF $ **FLOATING
C2094 S.n1887 VSUBS 0.01fF $ **FLOATING
C2095 S.n1888 VSUBS 0.02fF $ **FLOATING
C2096 S.n1889 VSUBS 0.08fF $ **FLOATING
C2097 S.n1890 VSUBS 0.06fF $ **FLOATING
C2098 S.n1891 VSUBS 0.03fF $ **FLOATING
C2099 S.n1892 VSUBS 0.03fF $ **FLOATING
C2100 S.n1893 VSUBS 0.99fF $ **FLOATING
C2101 S.n1894 VSUBS 0.35fF $ **FLOATING
C2102 S.n1895 VSUBS 1.85fF $ **FLOATING
C2103 S.n1896 VSUBS 1.97fF $ **FLOATING
C2104 S.t670 VSUBS 0.02fF
C2105 S.n1897 VSUBS 0.24fF $ **FLOATING
C2106 S.n1898 VSUBS 0.90fF $ **FLOATING
C2107 S.n1899 VSUBS 0.05fF $ **FLOATING
C2108 S.t575 VSUBS 0.02fF
C2109 S.n1900 VSUBS 0.12fF $ **FLOATING
C2110 S.n1901 VSUBS 0.14fF $ **FLOATING
C2111 S.n1903 VSUBS 1.87fF $ **FLOATING
C2112 S.n1904 VSUBS 0.07fF $ **FLOATING
C2113 S.n1905 VSUBS 0.04fF $ **FLOATING
C2114 S.n1906 VSUBS 0.05fF $ **FLOATING
C2115 S.n1907 VSUBS 0.86fF $ **FLOATING
C2116 S.n1908 VSUBS 0.01fF $ **FLOATING
C2117 S.n1909 VSUBS 0.01fF $ **FLOATING
C2118 S.n1910 VSUBS 0.01fF $ **FLOATING
C2119 S.n1911 VSUBS 0.07fF $ **FLOATING
C2120 S.n1912 VSUBS 0.68fF $ **FLOATING
C2121 S.n1913 VSUBS 0.71fF $ **FLOATING
C2122 S.t901 VSUBS 0.02fF
C2123 S.n1914 VSUBS 0.24fF $ **FLOATING
C2124 S.n1915 VSUBS 0.35fF $ **FLOATING
C2125 S.n1916 VSUBS 0.60fF $ **FLOATING
C2126 S.n1917 VSUBS 0.12fF $ **FLOATING
C2127 S.t545 VSUBS 0.02fF
C2128 S.n1918 VSUBS 0.14fF $ **FLOATING
C2129 S.n1920 VSUBS 0.69fF $ **FLOATING
C2130 S.n1921 VSUBS 0.22fF $ **FLOATING
C2131 S.n1922 VSUBS 0.22fF $ **FLOATING
C2132 S.n1923 VSUBS 0.69fF $ **FLOATING
C2133 S.n1924 VSUBS 1.14fF $ **FLOATING
C2134 S.n1925 VSUBS 0.22fF $ **FLOATING
C2135 S.n1926 VSUBS 0.25fF $ **FLOATING
C2136 S.n1927 VSUBS 0.09fF $ **FLOATING
C2137 S.n1928 VSUBS 2.29fF $ **FLOATING
C2138 S.t1016 VSUBS 0.02fF
C2139 S.n1929 VSUBS 0.24fF $ **FLOATING
C2140 S.n1930 VSUBS 0.90fF $ **FLOATING
C2141 S.n1931 VSUBS 0.05fF $ **FLOATING
C2142 S.t922 VSUBS 0.02fF
C2143 S.n1932 VSUBS 0.12fF $ **FLOATING
C2144 S.n1933 VSUBS 0.14fF $ **FLOATING
C2145 S.n1935 VSUBS 1.86fF $ **FLOATING
C2146 S.n1936 VSUBS 0.45fF $ **FLOATING
C2147 S.n1937 VSUBS 0.22fF $ **FLOATING
C2148 S.n1938 VSUBS 0.38fF $ **FLOATING
C2149 S.n1939 VSUBS 0.16fF $ **FLOATING
C2150 S.n1940 VSUBS 0.28fF $ **FLOATING
C2151 S.n1941 VSUBS 0.21fF $ **FLOATING
C2152 S.n1942 VSUBS 0.30fF $ **FLOATING
C2153 S.n1943 VSUBS 0.41fF $ **FLOATING
C2154 S.n1944 VSUBS 0.20fF $ **FLOATING
C2155 S.t136 VSUBS 0.02fF
C2156 S.n1945 VSUBS 0.24fF $ **FLOATING
C2157 S.n1946 VSUBS 0.35fF $ **FLOATING
C2158 S.n1947 VSUBS 0.60fF $ **FLOATING
C2159 S.n1948 VSUBS 0.12fF $ **FLOATING
C2160 S.t890 VSUBS 0.02fF
C2161 S.n1949 VSUBS 0.14fF $ **FLOATING
C2162 S.n1951 VSUBS 0.04fF $ **FLOATING
C2163 S.n1952 VSUBS 0.03fF $ **FLOATING
C2164 S.n1953 VSUBS 0.03fF $ **FLOATING
C2165 S.n1954 VSUBS 0.10fF $ **FLOATING
C2166 S.n1955 VSUBS 0.36fF $ **FLOATING
C2167 S.n1956 VSUBS 0.37fF $ **FLOATING
C2168 S.n1957 VSUBS 0.10fF $ **FLOATING
C2169 S.n1958 VSUBS 0.12fF $ **FLOATING
C2170 S.n1959 VSUBS 0.07fF $ **FLOATING
C2171 S.n1960 VSUBS 0.12fF $ **FLOATING
C2172 S.n1961 VSUBS 0.18fF $ **FLOATING
C2173 S.n1962 VSUBS 3.95fF $ **FLOATING
C2174 S.t251 VSUBS 0.02fF
C2175 S.n1963 VSUBS 0.24fF $ **FLOATING
C2176 S.n1964 VSUBS 0.90fF $ **FLOATING
C2177 S.n1965 VSUBS 0.05fF $ **FLOATING
C2178 S.t165 VSUBS 0.02fF
C2179 S.n1966 VSUBS 0.12fF $ **FLOATING
C2180 S.n1967 VSUBS 0.14fF $ **FLOATING
C2181 S.n1969 VSUBS 0.25fF $ **FLOATING
C2182 S.n1970 VSUBS 0.09fF $ **FLOATING
C2183 S.n1971 VSUBS 0.21fF $ **FLOATING
C2184 S.n1972 VSUBS 1.27fF $ **FLOATING
C2185 S.n1973 VSUBS 0.52fF $ **FLOATING
C2186 S.n1974 VSUBS 1.86fF $ **FLOATING
C2187 S.n1975 VSUBS 0.12fF $ **FLOATING
C2188 S.t1107 VSUBS 0.02fF
C2189 S.n1976 VSUBS 0.14fF $ **FLOATING
C2190 S.t1009 VSUBS 0.02fF
C2191 S.n1978 VSUBS 0.24fF $ **FLOATING
C2192 S.n1979 VSUBS 0.35fF $ **FLOATING
C2193 S.n1980 VSUBS 0.60fF $ **FLOATING
C2194 S.n1981 VSUBS 1.56fF $ **FLOATING
C2195 S.n1982 VSUBS 2.42fF $ **FLOATING
C2196 S.t271 VSUBS 0.02fF
C2197 S.n1983 VSUBS 0.24fF $ **FLOATING
C2198 S.n1984 VSUBS 0.90fF $ **FLOATING
C2199 S.n1985 VSUBS 0.05fF $ **FLOATING
C2200 S.t563 VSUBS 0.02fF
C2201 S.n1986 VSUBS 0.12fF $ **FLOATING
C2202 S.n1987 VSUBS 0.14fF $ **FLOATING
C2203 S.n1989 VSUBS 1.87fF $ **FLOATING
C2204 S.n1990 VSUBS 0.06fF $ **FLOATING
C2205 S.n1991 VSUBS 0.03fF $ **FLOATING
C2206 S.n1992 VSUBS 0.03fF $ **FLOATING
C2207 S.n1993 VSUBS 0.98fF $ **FLOATING
C2208 S.n1994 VSUBS 0.02fF $ **FLOATING
C2209 S.n1995 VSUBS 0.01fF $ **FLOATING
C2210 S.n1996 VSUBS 0.02fF $ **FLOATING
C2211 S.n1997 VSUBS 0.08fF $ **FLOATING
C2212 S.n1998 VSUBS 0.36fF $ **FLOATING
C2213 S.n1999 VSUBS 1.83fF $ **FLOATING
C2214 S.t246 VSUBS 0.02fF
C2215 S.n2000 VSUBS 0.24fF $ **FLOATING
C2216 S.n2001 VSUBS 0.35fF $ **FLOATING
C2217 S.n2002 VSUBS 0.60fF $ **FLOATING
C2218 S.n2003 VSUBS 0.12fF $ **FLOATING
C2219 S.t339 VSUBS 0.02fF
C2220 S.n2004 VSUBS 0.14fF $ **FLOATING
C2221 S.n2006 VSUBS 0.69fF $ **FLOATING
C2222 S.n2007 VSUBS 0.22fF $ **FLOATING
C2223 S.n2008 VSUBS 0.22fF $ **FLOATING
C2224 S.n2009 VSUBS 0.69fF $ **FLOATING
C2225 S.n2010 VSUBS 1.14fF $ **FLOATING
C2226 S.n2011 VSUBS 0.22fF $ **FLOATING
C2227 S.n2012 VSUBS 0.25fF $ **FLOATING
C2228 S.n2013 VSUBS 0.09fF $ **FLOATING
C2229 S.n2014 VSUBS 1.86fF $ **FLOATING
C2230 S.t617 VSUBS 0.02fF
C2231 S.n2015 VSUBS 0.24fF $ **FLOATING
C2232 S.n2016 VSUBS 0.90fF $ **FLOATING
C2233 S.n2017 VSUBS 0.05fF $ **FLOATING
C2234 S.t724 VSUBS 0.02fF
C2235 S.n2018 VSUBS 0.12fF $ **FLOATING
C2236 S.n2019 VSUBS 0.14fF $ **FLOATING
C2237 S.n2021 VSUBS 14.09fF $ **FLOATING
C2238 S.n2022 VSUBS 1.70fF $ **FLOATING
C2239 S.n2023 VSUBS 3.01fF $ **FLOATING
C2240 S.t1082 VSUBS 0.02fF
C2241 S.n2024 VSUBS 0.24fF $ **FLOATING
C2242 S.n2025 VSUBS 0.35fF $ **FLOATING
C2243 S.n2026 VSUBS 0.60fF $ **FLOATING
C2244 S.n2027 VSUBS 0.12fF $ **FLOATING
C2245 S.t728 VSUBS 0.02fF
C2246 S.n2028 VSUBS 0.14fF $ **FLOATING
C2247 S.n2030 VSUBS 0.31fF $ **FLOATING
C2248 S.n2031 VSUBS 0.22fF $ **FLOATING
C2249 S.n2032 VSUBS 0.65fF $ **FLOATING
C2250 S.n2033 VSUBS 0.94fF $ **FLOATING
C2251 S.n2034 VSUBS 0.22fF $ **FLOATING
C2252 S.n2035 VSUBS 0.20fF $ **FLOATING
C2253 S.n2036 VSUBS 0.20fF $ **FLOATING
C2254 S.n2037 VSUBS 0.06fF $ **FLOATING
C2255 S.n2038 VSUBS 0.09fF $ **FLOATING
C2256 S.n2039 VSUBS 0.09fF $ **FLOATING
C2257 S.n2040 VSUBS 1.97fF $ **FLOATING
C2258 S.t1114 VSUBS 0.02fF
C2259 S.n2041 VSUBS 0.12fF $ **FLOATING
C2260 S.n2042 VSUBS 0.14fF $ **FLOATING
C2261 S.t100 VSUBS 0.02fF
C2262 S.n2044 VSUBS 0.24fF $ **FLOATING
C2263 S.n2045 VSUBS 0.90fF $ **FLOATING
C2264 S.n2046 VSUBS 0.05fF $ **FLOATING
C2265 S.n2047 VSUBS 1.86fF $ **FLOATING
C2266 S.n2048 VSUBS 0.12fF $ **FLOATING
C2267 S.t688 VSUBS 0.02fF
C2268 S.n2049 VSUBS 0.14fF $ **FLOATING
C2269 S.t1071 VSUBS 0.02fF
C2270 S.n2051 VSUBS 0.12fF $ **FLOATING
C2271 S.n2052 VSUBS 0.14fF $ **FLOATING
C2272 S.t975 VSUBS 0.02fF
C2273 S.n2054 VSUBS 0.24fF $ **FLOATING
C2274 S.n2055 VSUBS 0.90fF $ **FLOATING
C2275 S.n2056 VSUBS 0.05fF $ **FLOATING
C2276 S.t606 VSUBS 0.02fF
C2277 S.n2057 VSUBS 0.24fF $ **FLOATING
C2278 S.n2058 VSUBS 0.35fF $ **FLOATING
C2279 S.n2059 VSUBS 0.60fF $ **FLOATING
C2280 S.n2060 VSUBS 0.31fF $ **FLOATING
C2281 S.n2061 VSUBS 1.08fF $ **FLOATING
C2282 S.n2062 VSUBS 0.15fF $ **FLOATING
C2283 S.n2063 VSUBS 2.08fF $ **FLOATING
C2284 S.n2064 VSUBS 2.91fF $ **FLOATING
C2285 S.n2065 VSUBS 1.86fF $ **FLOATING
C2286 S.n2066 VSUBS 0.12fF $ **FLOATING
C2287 S.t680 VSUBS 0.02fF
C2288 S.n2067 VSUBS 0.14fF $ **FLOATING
C2289 S.t597 VSUBS 0.02fF
C2290 S.n2069 VSUBS 0.24fF $ **FLOATING
C2291 S.n2070 VSUBS 0.35fF $ **FLOATING
C2292 S.n2071 VSUBS 0.60fF $ **FLOATING
C2293 S.n2072 VSUBS 0.91fF $ **FLOATING
C2294 S.n2073 VSUBS 0.31fF $ **FLOATING
C2295 S.n2074 VSUBS 0.91fF $ **FLOATING
C2296 S.n2075 VSUBS 1.08fF $ **FLOATING
C2297 S.n2076 VSUBS 0.15fF $ **FLOATING
C2298 S.n2077 VSUBS 4.90fF $ **FLOATING
C2299 S.t1058 VSUBS 0.02fF
C2300 S.n2078 VSUBS 0.12fF $ **FLOATING
C2301 S.n2079 VSUBS 0.14fF $ **FLOATING
C2302 S.t969 VSUBS 0.02fF
C2303 S.n2081 VSUBS 0.24fF $ **FLOATING
C2304 S.n2082 VSUBS 0.90fF $ **FLOATING
C2305 S.n2083 VSUBS 0.05fF $ **FLOATING
C2306 S.n2084 VSUBS 1.86fF $ **FLOATING
C2307 S.n2085 VSUBS 2.64fF $ **FLOATING
C2308 S.t943 VSUBS 0.02fF
C2309 S.n2086 VSUBS 0.24fF $ **FLOATING
C2310 S.n2087 VSUBS 0.35fF $ **FLOATING
C2311 S.n2088 VSUBS 0.60fF $ **FLOATING
C2312 S.n2089 VSUBS 0.12fF $ **FLOATING
C2313 S.t1025 VSUBS 0.02fF
C2314 S.n2090 VSUBS 0.14fF $ **FLOATING
C2315 S.n2092 VSUBS 1.86fF $ **FLOATING
C2316 S.n2093 VSUBS 2.64fF $ **FLOATING
C2317 S.t951 VSUBS 0.02fF
C2318 S.n2094 VSUBS 0.24fF $ **FLOATING
C2319 S.n2095 VSUBS 0.35fF $ **FLOATING
C2320 S.n2096 VSUBS 0.60fF $ **FLOATING
C2321 S.t215 VSUBS 0.02fF
C2322 S.n2097 VSUBS 0.24fF $ **FLOATING
C2323 S.n2098 VSUBS 0.90fF $ **FLOATING
C2324 S.n2099 VSUBS 0.05fF $ **FLOATING
C2325 S.t307 VSUBS 0.02fF
C2326 S.n2100 VSUBS 0.12fF $ **FLOATING
C2327 S.n2101 VSUBS 0.14fF $ **FLOATING
C2328 S.n2103 VSUBS 0.12fF $ **FLOATING
C2329 S.t1033 VSUBS 0.02fF
C2330 S.n2104 VSUBS 0.14fF $ **FLOATING
C2331 S.n2106 VSUBS 2.27fF $ **FLOATING
C2332 S.n2107 VSUBS 2.91fF $ **FLOATING
C2333 S.n2108 VSUBS 4.83fF $ **FLOATING
C2334 S.t298 VSUBS 0.02fF
C2335 S.n2109 VSUBS 0.12fF $ **FLOATING
C2336 S.n2110 VSUBS 0.14fF $ **FLOATING
C2337 S.t208 VSUBS 0.02fF
C2338 S.n2112 VSUBS 0.24fF $ **FLOATING
C2339 S.n2113 VSUBS 0.90fF $ **FLOATING
C2340 S.n2114 VSUBS 0.05fF $ **FLOATING
C2341 S.n2115 VSUBS 1.86fF $ **FLOATING
C2342 S.n2116 VSUBS 2.64fF $ **FLOATING
C2343 S.t184 VSUBS 0.02fF
C2344 S.n2117 VSUBS 0.24fF $ **FLOATING
C2345 S.n2118 VSUBS 0.35fF $ **FLOATING
C2346 S.n2119 VSUBS 0.60fF $ **FLOATING
C2347 S.n2120 VSUBS 0.12fF $ **FLOATING
C2348 S.t261 VSUBS 0.02fF
C2349 S.n2121 VSUBS 0.14fF $ **FLOATING
C2350 S.n2123 VSUBS 1.86fF $ **FLOATING
C2351 S.n2124 VSUBS 2.65fF $ **FLOATING
C2352 S.t192 VSUBS 0.02fF
C2353 S.n2125 VSUBS 0.24fF $ **FLOATING
C2354 S.n2126 VSUBS 0.35fF $ **FLOATING
C2355 S.n2127 VSUBS 0.60fF $ **FLOATING
C2356 S.t231 VSUBS 0.02fF
C2357 S.n2128 VSUBS 1.20fF $ **FLOATING
C2358 S.n2129 VSUBS 0.60fF $ **FLOATING
C2359 S.n2130 VSUBS 0.35fF $ **FLOATING
C2360 S.n2131 VSUBS 0.62fF $ **FLOATING
C2361 S.n2132 VSUBS 1.14fF $ **FLOATING
C2362 S.n2133 VSUBS 2.15fF $ **FLOATING
C2363 S.n2134 VSUBS 0.59fF $ **FLOATING
C2364 S.n2135 VSUBS 0.01fF $ **FLOATING
C2365 S.n2136 VSUBS 0.96fF $ **FLOATING
C2366 S.t21 VSUBS 14.53fF
C2367 S.n2137 VSUBS 14.40fF $ **FLOATING
C2368 S.n2139 VSUBS 0.37fF $ **FLOATING
C2369 S.n2140 VSUBS 0.23fF $ **FLOATING
C2370 S.n2141 VSUBS 2.87fF $ **FLOATING
C2371 S.n2142 VSUBS 2.43fF $ **FLOATING
C2372 S.n2143 VSUBS 1.94fF $ **FLOATING
C2373 S.n2144 VSUBS 3.89fF $ **FLOATING
C2374 S.n2145 VSUBS 0.25fF $ **FLOATING
C2375 S.n2146 VSUBS 0.01fF $ **FLOATING
C2376 S.t977 VSUBS 0.02fF
C2377 S.n2147 VSUBS 0.25fF $ **FLOATING
C2378 S.t365 VSUBS 0.02fF
C2379 S.n2148 VSUBS 0.94fF $ **FLOATING
C2380 S.n2149 VSUBS 0.70fF $ **FLOATING
C2381 S.n2150 VSUBS 0.77fF $ **FLOATING
C2382 S.n2151 VSUBS 1.91fF $ **FLOATING
C2383 S.n2152 VSUBS 1.86fF $ **FLOATING
C2384 S.n2153 VSUBS 0.12fF $ **FLOATING
C2385 S.t270 VSUBS 0.02fF
C2386 S.n2154 VSUBS 0.14fF $ **FLOATING
C2387 S.t580 VSUBS 0.02fF
C2388 S.n2156 VSUBS 0.24fF $ **FLOATING
C2389 S.n2157 VSUBS 0.35fF $ **FLOATING
C2390 S.n2158 VSUBS 0.60fF $ **FLOATING
C2391 S.n2159 VSUBS 1.50fF $ **FLOATING
C2392 S.n2160 VSUBS 2.96fF $ **FLOATING
C2393 S.t696 VSUBS 0.02fF
C2394 S.n2161 VSUBS 0.24fF $ **FLOATING
C2395 S.n2162 VSUBS 0.90fF $ **FLOATING
C2396 S.n2163 VSUBS 0.05fF $ **FLOATING
C2397 S.t598 VSUBS 0.02fF
C2398 S.n2164 VSUBS 0.12fF $ **FLOATING
C2399 S.n2165 VSUBS 0.14fF $ **FLOATING
C2400 S.t591 VSUBS 0.02fF
C2401 S.n2167 VSUBS 0.24fF $ **FLOATING
C2402 S.n2168 VSUBS 0.90fF $ **FLOATING
C2403 S.n2169 VSUBS 0.05fF $ **FLOATING
C2404 S.n2170 VSUBS 1.87fF $ **FLOATING
C2405 S.n2171 VSUBS 1.86fF $ **FLOATING
C2406 S.t472 VSUBS 0.02fF
C2407 S.n2172 VSUBS 0.24fF $ **FLOATING
C2408 S.n2173 VSUBS 0.35fF $ **FLOATING
C2409 S.n2174 VSUBS 0.60fF $ **FLOATING
C2410 S.n2175 VSUBS 0.12fF $ **FLOATING
C2411 S.t103 VSUBS 0.02fF
C2412 S.n2176 VSUBS 0.14fF $ **FLOATING
C2413 S.n2178 VSUBS 1.14fF $ **FLOATING
C2414 S.n2179 VSUBS 0.22fF $ **FLOATING
C2415 S.n2180 VSUBS 0.25fF $ **FLOATING
C2416 S.n2181 VSUBS 0.09fF $ **FLOATING
C2417 S.n2182 VSUBS 1.86fF $ **FLOATING
C2418 S.t994 VSUBS 0.02fF
C2419 S.n2183 VSUBS 0.12fF $ **FLOATING
C2420 S.n2184 VSUBS 0.14fF $ **FLOATING
C2421 S.n2186 VSUBS 0.77fF $ **FLOATING
C2422 S.n2187 VSUBS 1.92fF $ **FLOATING
C2423 S.n2188 VSUBS 1.86fF $ **FLOATING
C2424 S.n2189 VSUBS 0.12fF $ **FLOATING
C2425 S.t459 VSUBS 0.02fF
C2426 S.n2190 VSUBS 0.14fF $ **FLOATING
C2427 S.t817 VSUBS 0.02fF
C2428 S.n2192 VSUBS 0.24fF $ **FLOATING
C2429 S.n2193 VSUBS 0.35fF $ **FLOATING
C2430 S.n2194 VSUBS 0.60fF $ **FLOATING
C2431 S.n2195 VSUBS 1.82fF $ **FLOATING
C2432 S.n2196 VSUBS 2.96fF $ **FLOATING
C2433 S.t936 VSUBS 0.02fF
C2434 S.n2197 VSUBS 0.24fF $ **FLOATING
C2435 S.n2198 VSUBS 0.90fF $ **FLOATING
C2436 S.n2199 VSUBS 0.05fF $ **FLOATING
C2437 S.t840 VSUBS 0.02fF
C2438 S.n2200 VSUBS 0.12fF $ **FLOATING
C2439 S.n2201 VSUBS 0.14fF $ **FLOATING
C2440 S.n2203 VSUBS 1.87fF $ **FLOATING
C2441 S.n2204 VSUBS 1.73fF $ **FLOATING
C2442 S.t22 VSUBS 0.02fF
C2443 S.n2205 VSUBS 0.24fF $ **FLOATING
C2444 S.n2206 VSUBS 0.35fF $ **FLOATING
C2445 S.n2207 VSUBS 0.60fF $ **FLOATING
C2446 S.n2208 VSUBS 0.12fF $ **FLOATING
C2447 S.t800 VSUBS 0.02fF
C2448 S.n2209 VSUBS 0.14fF $ **FLOATING
C2449 S.n2211 VSUBS 1.14fF $ **FLOATING
C2450 S.n2212 VSUBS 0.22fF $ **FLOATING
C2451 S.n2213 VSUBS 0.25fF $ **FLOATING
C2452 S.n2214 VSUBS 0.09fF $ **FLOATING
C2453 S.n2215 VSUBS 2.41fF $ **FLOATING
C2454 S.t175 VSUBS 0.02fF
C2455 S.n2216 VSUBS 0.24fF $ **FLOATING
C2456 S.n2217 VSUBS 0.90fF $ **FLOATING
C2457 S.n2218 VSUBS 0.05fF $ **FLOATING
C2458 S.t60 VSUBS 0.02fF
C2459 S.n2219 VSUBS 0.12fF $ **FLOATING
C2460 S.n2220 VSUBS 0.14fF $ **FLOATING
C2461 S.n2222 VSUBS 1.86fF $ **FLOATING
C2462 S.n2223 VSUBS 0.47fF $ **FLOATING
C2463 S.n2224 VSUBS 0.09fF $ **FLOATING
C2464 S.n2225 VSUBS 0.32fF $ **FLOATING
C2465 S.n2226 VSUBS 0.30fF $ **FLOATING
C2466 S.n2227 VSUBS 0.76fF $ **FLOATING
C2467 S.n2228 VSUBS 0.58fF $ **FLOATING
C2468 S.t401 VSUBS 0.02fF
C2469 S.n2229 VSUBS 0.24fF $ **FLOATING
C2470 S.n2230 VSUBS 0.35fF $ **FLOATING
C2471 S.n2231 VSUBS 0.60fF $ **FLOATING
C2472 S.n2232 VSUBS 0.12fF $ **FLOATING
C2473 S.t9 VSUBS 0.02fF
C2474 S.n2233 VSUBS 0.14fF $ **FLOATING
C2475 S.n2235 VSUBS 2.58fF $ **FLOATING
C2476 S.n2236 VSUBS 2.13fF $ **FLOATING
C2477 S.t526 VSUBS 0.02fF
C2478 S.n2237 VSUBS 0.24fF $ **FLOATING
C2479 S.n2238 VSUBS 0.90fF $ **FLOATING
C2480 S.n2239 VSUBS 0.05fF $ **FLOATING
C2481 S.t426 VSUBS 0.02fF
C2482 S.n2240 VSUBS 0.12fF $ **FLOATING
C2483 S.n2241 VSUBS 0.14fF $ **FLOATING
C2484 S.n2243 VSUBS 0.77fF $ **FLOATING
C2485 S.n2244 VSUBS 2.27fF $ **FLOATING
C2486 S.n2245 VSUBS 1.86fF $ **FLOATING
C2487 S.n2246 VSUBS 0.12fF $ **FLOATING
C2488 S.t447 VSUBS 0.02fF
C2489 S.n2247 VSUBS 0.14fF $ **FLOATING
C2490 S.t742 VSUBS 0.02fF
C2491 S.n2249 VSUBS 0.24fF $ **FLOATING
C2492 S.n2250 VSUBS 0.35fF $ **FLOATING
C2493 S.n2251 VSUBS 0.60fF $ **FLOATING
C2494 S.n2252 VSUBS 1.37fF $ **FLOATING
C2495 S.n2253 VSUBS 0.70fF $ **FLOATING
C2496 S.n2254 VSUBS 1.13fF $ **FLOATING
C2497 S.n2255 VSUBS 0.35fF $ **FLOATING
C2498 S.n2256 VSUBS 2.00fF $ **FLOATING
C2499 S.t870 VSUBS 0.02fF
C2500 S.n2257 VSUBS 0.24fF $ **FLOATING
C2501 S.n2258 VSUBS 0.90fF $ **FLOATING
C2502 S.n2259 VSUBS 0.05fF $ **FLOATING
C2503 S.t766 VSUBS 0.02fF
C2504 S.n2260 VSUBS 0.12fF $ **FLOATING
C2505 S.n2261 VSUBS 0.14fF $ **FLOATING
C2506 S.n2263 VSUBS 1.87fF $ **FLOATING
C2507 S.n2264 VSUBS 1.86fF $ **FLOATING
C2508 S.t256 VSUBS 0.02fF
C2509 S.n2265 VSUBS 0.24fF $ **FLOATING
C2510 S.n2266 VSUBS 0.35fF $ **FLOATING
C2511 S.n2267 VSUBS 0.60fF $ **FLOATING
C2512 S.n2268 VSUBS 0.12fF $ **FLOATING
C2513 S.t352 VSUBS 0.02fF
C2514 S.n2269 VSUBS 0.14fF $ **FLOATING
C2515 S.n2271 VSUBS 1.14fF $ **FLOATING
C2516 S.n2272 VSUBS 0.22fF $ **FLOATING
C2517 S.n2273 VSUBS 0.25fF $ **FLOATING
C2518 S.n2274 VSUBS 0.09fF $ **FLOATING
C2519 S.n2275 VSUBS 1.86fF $ **FLOATING
C2520 S.t625 VSUBS 0.02fF
C2521 S.n2276 VSUBS 0.24fF $ **FLOATING
C2522 S.n2277 VSUBS 0.90fF $ **FLOATING
C2523 S.n2278 VSUBS 0.05fF $ **FLOATING
C2524 S.t737 VSUBS 0.02fF
C2525 S.n2279 VSUBS 0.12fF $ **FLOATING
C2526 S.n2280 VSUBS 0.14fF $ **FLOATING
C2527 S.n2282 VSUBS 14.09fF $ **FLOATING
C2528 S.n2283 VSUBS 2.70fF $ **FLOATING
C2529 S.n2284 VSUBS 1.58fF $ **FLOATING
C2530 S.n2285 VSUBS 0.12fF $ **FLOATING
C2531 S.t1062 VSUBS 0.02fF
C2532 S.n2286 VSUBS 0.14fF $ **FLOATING
C2533 S.t476 VSUBS 0.02fF
C2534 S.n2288 VSUBS 0.24fF $ **FLOATING
C2535 S.n2289 VSUBS 0.35fF $ **FLOATING
C2536 S.n2290 VSUBS 0.60fF $ **FLOATING
C2537 S.n2291 VSUBS 0.07fF $ **FLOATING
C2538 S.n2292 VSUBS 0.01fF $ **FLOATING
C2539 S.n2293 VSUBS 0.23fF $ **FLOATING
C2540 S.n2294 VSUBS 1.15fF $ **FLOATING
C2541 S.n2295 VSUBS 1.33fF $ **FLOATING
C2542 S.n2296 VSUBS 2.27fF $ **FLOATING
C2543 S.t1001 VSUBS 0.02fF
C2544 S.n2297 VSUBS 0.12fF $ **FLOATING
C2545 S.n2298 VSUBS 0.14fF $ **FLOATING
C2546 S.t1070 VSUBS 0.02fF
C2547 S.n2300 VSUBS 0.24fF $ **FLOATING
C2548 S.n2301 VSUBS 0.90fF $ **FLOATING
C2549 S.n2302 VSUBS 0.05fF $ **FLOATING
C2550 S.t8 VSUBS 32.33fF
C2551 S.t565 VSUBS 0.02fF
C2552 S.n2303 VSUBS 0.24fF $ **FLOATING
C2553 S.n2304 VSUBS 0.90fF $ **FLOATING
C2554 S.n2305 VSUBS 0.05fF $ **FLOATING
C2555 S.t654 VSUBS 0.02fF
C2556 S.n2306 VSUBS 0.12fF $ **FLOATING
C2557 S.n2307 VSUBS 0.14fF $ **FLOATING
C2558 S.n2309 VSUBS 0.12fF $ **FLOATING
C2559 S.t275 VSUBS 0.02fF
C2560 S.n2310 VSUBS 0.14fF $ **FLOATING
C2561 S.n2312 VSUBS 5.11fF $ **FLOATING
C2562 S.n2313 VSUBS 5.38fF $ **FLOATING
C2563 S.t643 VSUBS 0.02fF
C2564 S.n2314 VSUBS 0.12fF $ **FLOATING
C2565 S.n2315 VSUBS 0.14fF $ **FLOATING
C2566 S.t556 VSUBS 0.02fF
C2567 S.n2317 VSUBS 0.24fF $ **FLOATING
C2568 S.n2318 VSUBS 0.90fF $ **FLOATING
C2569 S.n2319 VSUBS 0.05fF $ **FLOATING
C2570 S.t164 VSUBS 31.95fF
C2571 S.t566 VSUBS 0.02fF
C2572 S.n2320 VSUBS 0.01fF $ **FLOATING
C2573 S.n2321 VSUBS 0.25fF $ **FLOATING
C2574 S.t1095 VSUBS 0.02fF
C2575 S.n2323 VSUBS 1.18fF $ **FLOATING
C2576 S.n2324 VSUBS 0.05fF $ **FLOATING
C2577 S.t968 VSUBS 0.02fF
C2578 S.n2325 VSUBS 0.63fF $ **FLOATING
C2579 S.n2326 VSUBS 0.60fF $ **FLOATING
C2580 S.n2327 VSUBS 8.88fF $ **FLOATING
C2581 S.n2328 VSUBS 8.88fF $ **FLOATING
C2582 S.n2329 VSUBS 0.59fF $ **FLOATING
C2583 S.n2330 VSUBS 0.21fF $ **FLOATING
C2584 S.n2331 VSUBS 0.59fF $ **FLOATING
C2585 S.n2332 VSUBS 2.55fF $ **FLOATING
C2586 S.n2333 VSUBS 0.28fF $ **FLOATING
C2587 S.t135 VSUBS 14.53fF
C2588 S.n2334 VSUBS 15.80fF $ **FLOATING
C2589 S.n2335 VSUBS 0.76fF $ **FLOATING
C2590 S.n2336 VSUBS 0.27fF $ **FLOATING
C2591 S.n2337 VSUBS 3.96fF $ **FLOATING
C2592 S.n2338 VSUBS 1.34fF $ **FLOATING
C2593 S.n2339 VSUBS 0.01fF $ **FLOATING
C2594 S.n2340 VSUBS 0.02fF $ **FLOATING
C2595 S.n2341 VSUBS 0.03fF $ **FLOATING
C2596 S.n2342 VSUBS 0.04fF $ **FLOATING
C2597 S.n2343 VSUBS 0.17fF $ **FLOATING
C2598 S.n2344 VSUBS 0.01fF $ **FLOATING
C2599 S.n2345 VSUBS 0.02fF $ **FLOATING
C2600 S.n2346 VSUBS 0.01fF $ **FLOATING
C2601 S.n2347 VSUBS 0.01fF $ **FLOATING
C2602 S.n2348 VSUBS 0.01fF $ **FLOATING
C2603 S.n2349 VSUBS 0.01fF $ **FLOATING
C2604 S.n2350 VSUBS 0.01fF $ **FLOATING
C2605 S.n2351 VSUBS 0.01fF $ **FLOATING
C2606 S.n2352 VSUBS 0.02fF $ **FLOATING
C2607 S.n2353 VSUBS 0.05fF $ **FLOATING
C2608 S.n2354 VSUBS 0.04fF $ **FLOATING
C2609 S.n2355 VSUBS 0.11fF $ **FLOATING
C2610 S.n2356 VSUBS 0.37fF $ **FLOATING
C2611 S.n2357 VSUBS 0.20fF $ **FLOATING
C2612 S.n2358 VSUBS 4.34fF $ **FLOATING
C2613 S.n2359 VSUBS 0.24fF $ **FLOATING
C2614 S.n2360 VSUBS 1.48fF $ **FLOATING
C2615 S.n2361 VSUBS 1.29fF $ **FLOATING
C2616 S.n2362 VSUBS 0.27fF $ **FLOATING
C2617 S.n2363 VSUBS 1.87fF $ **FLOATING
C2618 S.n2364 VSUBS 0.06fF $ **FLOATING
C2619 S.n2365 VSUBS 0.03fF $ **FLOATING
C2620 S.n2366 VSUBS 0.03fF $ **FLOATING
C2621 S.n2367 VSUBS 0.98fF $ **FLOATING
C2622 S.n2368 VSUBS 0.02fF $ **FLOATING
C2623 S.n2369 VSUBS 0.01fF $ **FLOATING
C2624 S.n2370 VSUBS 0.02fF $ **FLOATING
C2625 S.n2371 VSUBS 0.08fF $ **FLOATING
C2626 S.n2372 VSUBS 0.36fF $ **FLOATING
C2627 S.n2373 VSUBS 1.83fF $ **FLOATING
C2628 S.t122 VSUBS 0.02fF
C2629 S.n2374 VSUBS 0.24fF $ **FLOATING
C2630 S.n2375 VSUBS 0.35fF $ **FLOATING
C2631 S.n2376 VSUBS 0.60fF $ **FLOATING
C2632 S.n2377 VSUBS 0.12fF $ **FLOATING
C2633 S.t880 VSUBS 0.02fF
C2634 S.n2378 VSUBS 0.14fF $ **FLOATING
C2635 S.n2380 VSUBS 0.69fF $ **FLOATING
C2636 S.n2381 VSUBS 0.22fF $ **FLOATING
C2637 S.n2382 VSUBS 0.22fF $ **FLOATING
C2638 S.n2383 VSUBS 0.69fF $ **FLOATING
C2639 S.n2384 VSUBS 1.14fF $ **FLOATING
C2640 S.n2385 VSUBS 0.22fF $ **FLOATING
C2641 S.n2386 VSUBS 0.25fF $ **FLOATING
C2642 S.n2387 VSUBS 0.09fF $ **FLOATING
C2643 S.n2388 VSUBS 1.86fF $ **FLOATING
C2644 S.t244 VSUBS 0.02fF
C2645 S.n2389 VSUBS 0.24fF $ **FLOATING
C2646 S.n2390 VSUBS 0.90fF $ **FLOATING
C2647 S.n2391 VSUBS 0.05fF $ **FLOATING
C2648 S.t155 VSUBS 0.02fF
C2649 S.n2392 VSUBS 0.12fF $ **FLOATING
C2650 S.n2393 VSUBS 0.14fF $ **FLOATING
C2651 S.n2395 VSUBS 0.25fF $ **FLOATING
C2652 S.n2396 VSUBS 0.09fF $ **FLOATING
C2653 S.n2397 VSUBS 0.21fF $ **FLOATING
C2654 S.n2398 VSUBS 0.91fF $ **FLOATING
C2655 S.n2399 VSUBS 0.44fF $ **FLOATING
C2656 S.n2400 VSUBS 1.86fF $ **FLOATING
C2657 S.n2401 VSUBS 0.12fF $ **FLOATING
C2658 S.t699 VSUBS 0.02fF
C2659 S.n2402 VSUBS 0.14fF $ **FLOATING
C2660 S.t1054 VSUBS 0.02fF
C2661 S.n2404 VSUBS 0.24fF $ **FLOATING
C2662 S.n2405 VSUBS 0.35fF $ **FLOATING
C2663 S.n2406 VSUBS 0.60fF $ **FLOATING
C2664 S.n2407 VSUBS 0.02fF $ **FLOATING
C2665 S.n2408 VSUBS 0.01fF $ **FLOATING
C2666 S.n2409 VSUBS 0.02fF $ **FLOATING
C2667 S.n2410 VSUBS 0.08fF $ **FLOATING
C2668 S.n2411 VSUBS 0.06fF $ **FLOATING
C2669 S.n2412 VSUBS 0.03fF $ **FLOATING
C2670 S.n2413 VSUBS 0.03fF $ **FLOATING
C2671 S.n2414 VSUBS 0.99fF $ **FLOATING
C2672 S.n2415 VSUBS 0.35fF $ **FLOATING
C2673 S.n2416 VSUBS 1.85fF $ **FLOATING
C2674 S.n2417 VSUBS 1.97fF $ **FLOATING
C2675 S.t76 VSUBS 0.02fF
C2676 S.n2418 VSUBS 0.24fF $ **FLOATING
C2677 S.n2419 VSUBS 0.90fF $ **FLOATING
C2678 S.n2420 VSUBS 0.05fF $ **FLOATING
C2679 S.t1083 VSUBS 0.02fF
C2680 S.n2421 VSUBS 0.12fF $ **FLOATING
C2681 S.n2422 VSUBS 0.14fF $ **FLOATING
C2682 S.n2424 VSUBS 1.87fF $ **FLOATING
C2683 S.n2425 VSUBS 0.04fF $ **FLOATING
C2684 S.n2426 VSUBS 0.07fF $ **FLOATING
C2685 S.n2427 VSUBS 0.05fF $ **FLOATING
C2686 S.n2428 VSUBS 0.86fF $ **FLOATING
C2687 S.n2429 VSUBS 0.01fF $ **FLOATING
C2688 S.n2430 VSUBS 0.01fF $ **FLOATING
C2689 S.n2431 VSUBS 0.01fF $ **FLOATING
C2690 S.n2432 VSUBS 0.07fF $ **FLOATING
C2691 S.n2433 VSUBS 0.68fF $ **FLOATING
C2692 S.n2434 VSUBS 0.71fF $ **FLOATING
C2693 S.t295 VSUBS 0.02fF
C2694 S.n2435 VSUBS 0.24fF $ **FLOATING
C2695 S.n2436 VSUBS 0.35fF $ **FLOATING
C2696 S.n2437 VSUBS 0.60fF $ **FLOATING
C2697 S.n2438 VSUBS 0.12fF $ **FLOATING
C2698 S.t1040 VSUBS 0.02fF
C2699 S.n2439 VSUBS 0.14fF $ **FLOATING
C2700 S.n2441 VSUBS 0.69fF $ **FLOATING
C2701 S.n2442 VSUBS 0.22fF $ **FLOATING
C2702 S.n2443 VSUBS 0.22fF $ **FLOATING
C2703 S.n2444 VSUBS 0.69fF $ **FLOATING
C2704 S.n2445 VSUBS 1.14fF $ **FLOATING
C2705 S.n2446 VSUBS 0.22fF $ **FLOATING
C2706 S.n2447 VSUBS 0.25fF $ **FLOATING
C2707 S.n2448 VSUBS 0.09fF $ **FLOATING
C2708 S.n2449 VSUBS 2.29fF $ **FLOATING
C2709 S.t440 VSUBS 0.02fF
C2710 S.n2450 VSUBS 0.24fF $ **FLOATING
C2711 S.n2451 VSUBS 0.90fF $ **FLOATING
C2712 S.n2452 VSUBS 0.05fF $ **FLOATING
C2713 S.t315 VSUBS 0.02fF
C2714 S.n2453 VSUBS 0.12fF $ **FLOATING
C2715 S.n2454 VSUBS 0.14fF $ **FLOATING
C2716 S.n2456 VSUBS 1.86fF $ **FLOATING
C2717 S.n2457 VSUBS 0.45fF $ **FLOATING
C2718 S.n2458 VSUBS 0.22fF $ **FLOATING
C2719 S.n2459 VSUBS 0.38fF $ **FLOATING
C2720 S.n2460 VSUBS 0.16fF $ **FLOATING
C2721 S.n2461 VSUBS 0.28fF $ **FLOATING
C2722 S.n2462 VSUBS 0.21fF $ **FLOATING
C2723 S.n2463 VSUBS 0.30fF $ **FLOATING
C2724 S.n2464 VSUBS 0.41fF $ **FLOATING
C2725 S.n2465 VSUBS 0.20fF $ **FLOATING
C2726 S.t635 VSUBS 0.02fF
C2727 S.n2466 VSUBS 0.24fF $ **FLOATING
C2728 S.n2467 VSUBS 0.35fF $ **FLOATING
C2729 S.n2468 VSUBS 0.60fF $ **FLOATING
C2730 S.n2469 VSUBS 0.12fF $ **FLOATING
C2731 S.t282 VSUBS 0.02fF
C2732 S.n2470 VSUBS 0.14fF $ **FLOATING
C2733 S.n2472 VSUBS 0.04fF $ **FLOATING
C2734 S.n2473 VSUBS 0.03fF $ **FLOATING
C2735 S.n2474 VSUBS 0.03fF $ **FLOATING
C2736 S.n2475 VSUBS 0.10fF $ **FLOATING
C2737 S.n2476 VSUBS 0.36fF $ **FLOATING
C2738 S.n2477 VSUBS 0.37fF $ **FLOATING
C2739 S.n2478 VSUBS 0.10fF $ **FLOATING
C2740 S.n2479 VSUBS 0.12fF $ **FLOATING
C2741 S.n2480 VSUBS 0.07fF $ **FLOATING
C2742 S.n2481 VSUBS 0.12fF $ **FLOATING
C2743 S.n2482 VSUBS 0.18fF $ **FLOATING
C2744 S.n2483 VSUBS 3.95fF $ **FLOATING
C2745 S.t776 VSUBS 0.02fF
C2746 S.n2484 VSUBS 0.24fF $ **FLOATING
C2747 S.n2485 VSUBS 0.90fF $ **FLOATING
C2748 S.n2486 VSUBS 0.05fF $ **FLOATING
C2749 S.t660 VSUBS 0.02fF
C2750 S.n2487 VSUBS 0.12fF $ **FLOATING
C2751 S.n2488 VSUBS 0.14fF $ **FLOATING
C2752 S.n2490 VSUBS 0.25fF $ **FLOATING
C2753 S.n2491 VSUBS 0.09fF $ **FLOATING
C2754 S.n2492 VSUBS 0.21fF $ **FLOATING
C2755 S.n2493 VSUBS 1.27fF $ **FLOATING
C2756 S.n2494 VSUBS 0.52fF $ **FLOATING
C2757 S.n2495 VSUBS 1.86fF $ **FLOATING
C2758 S.n2496 VSUBS 0.12fF $ **FLOATING
C2759 S.t623 VSUBS 0.02fF
C2760 S.n2497 VSUBS 0.14fF $ **FLOATING
C2761 S.t986 VSUBS 0.02fF
C2762 S.n2499 VSUBS 0.24fF $ **FLOATING
C2763 S.n2500 VSUBS 0.35fF $ **FLOATING
C2764 S.n2501 VSUBS 0.60fF $ **FLOATING
C2765 S.n2502 VSUBS 1.56fF $ **FLOATING
C2766 S.n2503 VSUBS 2.42fF $ **FLOATING
C2767 S.t1123 VSUBS 0.02fF
C2768 S.n2504 VSUBS 0.24fF $ **FLOATING
C2769 S.n2505 VSUBS 0.90fF $ **FLOATING
C2770 S.n2506 VSUBS 0.05fF $ **FLOATING
C2771 S.t1010 VSUBS 0.02fF
C2772 S.n2507 VSUBS 0.12fF $ **FLOATING
C2773 S.n2508 VSUBS 0.14fF $ **FLOATING
C2774 S.n2510 VSUBS 1.87fF $ **FLOATING
C2775 S.n2511 VSUBS 0.06fF $ **FLOATING
C2776 S.n2512 VSUBS 0.03fF $ **FLOATING
C2777 S.n2513 VSUBS 0.03fF $ **FLOATING
C2778 S.n2514 VSUBS 0.98fF $ **FLOATING
C2779 S.n2515 VSUBS 0.02fF $ **FLOATING
C2780 S.n2516 VSUBS 0.01fF $ **FLOATING
C2781 S.n2517 VSUBS 0.02fF $ **FLOATING
C2782 S.n2518 VSUBS 0.08fF $ **FLOATING
C2783 S.n2519 VSUBS 0.36fF $ **FLOATING
C2784 S.n2520 VSUBS 1.83fF $ **FLOATING
C2785 S.t268 VSUBS 0.02fF
C2786 S.n2521 VSUBS 0.24fF $ **FLOATING
C2787 S.n2522 VSUBS 0.35fF $ **FLOATING
C2788 S.n2523 VSUBS 0.60fF $ **FLOATING
C2789 S.n2524 VSUBS 0.12fF $ **FLOATING
C2790 S.t371 VSUBS 0.02fF
C2791 S.n2525 VSUBS 0.14fF $ **FLOATING
C2792 S.n2527 VSUBS 0.69fF $ **FLOATING
C2793 S.n2528 VSUBS 0.22fF $ **FLOATING
C2794 S.n2529 VSUBS 0.22fF $ **FLOATING
C2795 S.n2530 VSUBS 0.69fF $ **FLOATING
C2796 S.n2531 VSUBS 1.14fF $ **FLOATING
C2797 S.n2532 VSUBS 0.22fF $ **FLOATING
C2798 S.n2533 VSUBS 0.25fF $ **FLOATING
C2799 S.n2534 VSUBS 0.09fF $ **FLOATING
C2800 S.n2535 VSUBS 1.86fF $ **FLOATING
C2801 S.t634 VSUBS 0.02fF
C2802 S.n2536 VSUBS 0.24fF $ **FLOATING
C2803 S.n2537 VSUBS 0.90fF $ **FLOATING
C2804 S.n2538 VSUBS 0.05fF $ **FLOATING
C2805 S.t303 VSUBS 0.02fF
C2806 S.n2539 VSUBS 0.12fF $ **FLOATING
C2807 S.n2540 VSUBS 0.14fF $ **FLOATING
C2808 S.n2542 VSUBS 14.09fF $ **FLOATING
C2809 S.n2543 VSUBS 0.06fF $ **FLOATING
C2810 S.n2544 VSUBS 0.20fF $ **FLOATING
C2811 S.n2545 VSUBS 0.09fF $ **FLOATING
C2812 S.n2546 VSUBS 0.20fF $ **FLOATING
C2813 S.n2547 VSUBS 0.09fF $ **FLOATING
C2814 S.n2548 VSUBS 0.30fF $ **FLOATING
C2815 S.n2549 VSUBS 0.69fF $ **FLOATING
C2816 S.n2550 VSUBS 0.44fF $ **FLOATING
C2817 S.n2551 VSUBS 2.30fF $ **FLOATING
C2818 S.n2552 VSUBS 0.12fF $ **FLOATING
C2819 S.t485 VSUBS 0.02fF
C2820 S.n2553 VSUBS 0.14fF $ **FLOATING
C2821 S.t844 VSUBS 0.02fF
C2822 S.n2555 VSUBS 0.24fF $ **FLOATING
C2823 S.n2556 VSUBS 0.35fF $ **FLOATING
C2824 S.n2557 VSUBS 0.60fF $ **FLOATING
C2825 S.n2558 VSUBS 1.88fF $ **FLOATING
C2826 S.n2559 VSUBS 0.17fF $ **FLOATING
C2827 S.n2560 VSUBS 0.76fF $ **FLOATING
C2828 S.n2561 VSUBS 0.31fF $ **FLOATING
C2829 S.n2562 VSUBS 0.25fF $ **FLOATING
C2830 S.n2563 VSUBS 0.29fF $ **FLOATING
C2831 S.n2564 VSUBS 0.46fF $ **FLOATING
C2832 S.n2565 VSUBS 0.16fF $ **FLOATING
C2833 S.n2566 VSUBS 1.90fF $ **FLOATING
C2834 S.t863 VSUBS 0.02fF
C2835 S.n2567 VSUBS 0.12fF $ **FLOATING
C2836 S.n2568 VSUBS 0.14fF $ **FLOATING
C2837 S.t958 VSUBS 0.02fF
C2838 S.n2570 VSUBS 0.24fF $ **FLOATING
C2839 S.n2571 VSUBS 0.90fF $ **FLOATING
C2840 S.n2572 VSUBS 0.05fF $ **FLOATING
C2841 S.n2573 VSUBS 1.86fF $ **FLOATING
C2842 S.n2574 VSUBS 0.12fF $ **FLOATING
C2843 S.t720 VSUBS 0.02fF
C2844 S.n2575 VSUBS 0.14fF $ **FLOATING
C2845 S.t1102 VSUBS 0.02fF
C2846 S.n2577 VSUBS 0.12fF $ **FLOATING
C2847 S.n2578 VSUBS 0.14fF $ **FLOATING
C2848 S.t995 VSUBS 0.02fF
C2849 S.n2580 VSUBS 0.24fF $ **FLOATING
C2850 S.n2581 VSUBS 0.90fF $ **FLOATING
C2851 S.n2582 VSUBS 0.05fF $ **FLOATING
C2852 S.t622 VSUBS 0.02fF
C2853 S.n2583 VSUBS 0.24fF $ **FLOATING
C2854 S.n2584 VSUBS 0.35fF $ **FLOATING
C2855 S.n2585 VSUBS 0.60fF $ **FLOATING
C2856 S.n2586 VSUBS 0.31fF $ **FLOATING
C2857 S.n2587 VSUBS 1.08fF $ **FLOATING
C2858 S.n2588 VSUBS 0.15fF $ **FLOATING
C2859 S.n2589 VSUBS 2.08fF $ **FLOATING
C2860 S.n2590 VSUBS 2.91fF $ **FLOATING
C2861 S.n2591 VSUBS 1.86fF $ **FLOATING
C2862 S.n2592 VSUBS 0.12fF $ **FLOATING
C2863 S.t705 VSUBS 0.02fF
C2864 S.n2593 VSUBS 0.14fF $ **FLOATING
C2865 S.t615 VSUBS 0.02fF
C2866 S.n2595 VSUBS 0.24fF $ **FLOATING
C2867 S.n2596 VSUBS 0.35fF $ **FLOATING
C2868 S.n2597 VSUBS 0.60fF $ **FLOATING
C2869 S.n2598 VSUBS 0.91fF $ **FLOATING
C2870 S.n2599 VSUBS 0.31fF $ **FLOATING
C2871 S.n2600 VSUBS 0.91fF $ **FLOATING
C2872 S.n2601 VSUBS 1.08fF $ **FLOATING
C2873 S.n2602 VSUBS 0.15fF $ **FLOATING
C2874 S.n2603 VSUBS 4.90fF $ **FLOATING
C2875 S.t1091 VSUBS 0.02fF
C2876 S.n2604 VSUBS 0.12fF $ **FLOATING
C2877 S.n2605 VSUBS 0.14fF $ **FLOATING
C2878 S.t985 VSUBS 0.02fF
C2879 S.n2607 VSUBS 0.24fF $ **FLOATING
C2880 S.n2608 VSUBS 0.90fF $ **FLOATING
C2881 S.n2609 VSUBS 0.05fF $ **FLOATING
C2882 S.n2610 VSUBS 1.86fF $ **FLOATING
C2883 S.n2611 VSUBS 2.64fF $ **FLOATING
C2884 S.t967 VSUBS 0.02fF
C2885 S.n2612 VSUBS 0.24fF $ **FLOATING
C2886 S.n2613 VSUBS 0.35fF $ **FLOATING
C2887 S.n2614 VSUBS 0.60fF $ **FLOATING
C2888 S.n2615 VSUBS 0.12fF $ **FLOATING
C2889 S.t1044 VSUBS 0.02fF
C2890 S.n2616 VSUBS 0.14fF $ **FLOATING
C2891 S.n2618 VSUBS 1.86fF $ **FLOATING
C2892 S.n2619 VSUBS 2.64fF $ **FLOATING
C2893 S.t974 VSUBS 0.02fF
C2894 S.n2620 VSUBS 0.24fF $ **FLOATING
C2895 S.n2621 VSUBS 0.35fF $ **FLOATING
C2896 S.n2622 VSUBS 0.60fF $ **FLOATING
C2897 S.t238 VSUBS 0.02fF
C2898 S.n2623 VSUBS 0.24fF $ **FLOATING
C2899 S.n2624 VSUBS 0.90fF $ **FLOATING
C2900 S.n2625 VSUBS 0.05fF $ **FLOATING
C2901 S.t334 VSUBS 0.02fF
C2902 S.n2626 VSUBS 0.12fF $ **FLOATING
C2903 S.n2627 VSUBS 0.14fF $ **FLOATING
C2904 S.n2629 VSUBS 0.12fF $ **FLOATING
C2905 S.t1055 VSUBS 0.02fF
C2906 S.n2630 VSUBS 0.14fF $ **FLOATING
C2907 S.n2632 VSUBS 2.27fF $ **FLOATING
C2908 S.n2633 VSUBS 2.91fF $ **FLOATING
C2909 S.n2634 VSUBS 5.10fF $ **FLOATING
C2910 S.t319 VSUBS 0.02fF
C2911 S.n2635 VSUBS 0.12fF $ **FLOATING
C2912 S.n2636 VSUBS 0.14fF $ **FLOATING
C2913 S.t225 VSUBS 0.02fF
C2914 S.n2638 VSUBS 0.24fF $ **FLOATING
C2915 S.n2639 VSUBS 0.90fF $ **FLOATING
C2916 S.n2640 VSUBS 0.05fF $ **FLOATING
C2917 S.n2641 VSUBS 1.86fF $ **FLOATING
C2918 S.n2642 VSUBS 2.64fF $ **FLOATING
C2919 S.t206 VSUBS 0.02fF
C2920 S.n2643 VSUBS 0.24fF $ **FLOATING
C2921 S.n2644 VSUBS 0.35fF $ **FLOATING
C2922 S.n2645 VSUBS 0.60fF $ **FLOATING
C2923 S.n2646 VSUBS 0.12fF $ **FLOATING
C2924 S.t284 VSUBS 0.02fF
C2925 S.n2647 VSUBS 0.14fF $ **FLOATING
C2926 S.n2649 VSUBS 4.84fF $ **FLOATING
C2927 S.t663 VSUBS 0.02fF
C2928 S.n2650 VSUBS 0.12fF $ **FLOATING
C2929 S.n2651 VSUBS 0.14fF $ **FLOATING
C2930 S.t574 VSUBS 0.02fF
C2931 S.n2653 VSUBS 0.24fF $ **FLOATING
C2932 S.n2654 VSUBS 0.90fF $ **FLOATING
C2933 S.n2655 VSUBS 0.05fF $ **FLOATING
C2934 S.n2656 VSUBS 1.86fF $ **FLOATING
C2935 S.n2657 VSUBS 2.64fF $ **FLOATING
C2936 S.t553 VSUBS 0.02fF
C2937 S.n2658 VSUBS 0.24fF $ **FLOATING
C2938 S.n2659 VSUBS 0.35fF $ **FLOATING
C2939 S.n2660 VSUBS 0.60fF $ **FLOATING
C2940 S.n2661 VSUBS 0.12fF $ **FLOATING
C2941 S.t627 VSUBS 0.02fF
C2942 S.n2662 VSUBS 0.14fF $ **FLOATING
C2943 S.n2664 VSUBS 1.86fF $ **FLOATING
C2944 S.n2665 VSUBS 2.65fF $ **FLOATING
C2945 S.t564 VSUBS 0.02fF
C2946 S.n2666 VSUBS 0.24fF $ **FLOATING
C2947 S.n2667 VSUBS 0.35fF $ **FLOATING
C2948 S.n2668 VSUBS 0.60fF $ **FLOATING
C2949 S.t1088 VSUBS 0.02fF
C2950 S.n2669 VSUBS 1.20fF $ **FLOATING
C2951 S.n2670 VSUBS 0.36fF $ **FLOATING
C2952 S.n2671 VSUBS 1.21fF $ **FLOATING
C2953 S.n2672 VSUBS 0.60fF $ **FLOATING
C2954 S.n2673 VSUBS 0.35fF $ **FLOATING
C2955 S.n2674 VSUBS 0.62fF $ **FLOATING
C2956 S.n2675 VSUBS 1.14fF $ **FLOATING
C2957 S.n2676 VSUBS 2.15fF $ **FLOATING
C2958 S.n2677 VSUBS 0.59fF $ **FLOATING
C2959 S.n2678 VSUBS 0.01fF $ **FLOATING
C2960 S.n2679 VSUBS 0.96fF $ **FLOATING
C2961 S.t140 VSUBS 14.53fF
C2962 S.n2680 VSUBS 14.40fF $ **FLOATING
C2963 S.n2682 VSUBS 0.37fF $ **FLOATING
C2964 S.n2683 VSUBS 0.23fF $ **FLOATING
C2965 S.n2684 VSUBS 2.76fF $ **FLOATING
C2966 S.n2685 VSUBS 2.43fF $ **FLOATING
C2967 S.n2686 VSUBS 3.96fF $ **FLOATING
C2968 S.n2687 VSUBS 0.25fF $ **FLOATING
C2969 S.n2688 VSUBS 0.01fF $ **FLOATING
C2970 S.t731 VSUBS 0.02fF
C2971 S.n2689 VSUBS 0.25fF $ **FLOATING
C2972 S.t108 VSUBS 0.02fF
C2973 S.n2690 VSUBS 0.94fF $ **FLOATING
C2974 S.n2691 VSUBS 0.70fF $ **FLOATING
C2975 S.n2692 VSUBS 1.87fF $ **FLOATING
C2976 S.n2693 VSUBS 1.86fF $ **FLOATING
C2977 S.t318 VSUBS 0.02fF
C2978 S.n2694 VSUBS 0.24fF $ **FLOATING
C2979 S.n2695 VSUBS 0.35fF $ **FLOATING
C2980 S.n2696 VSUBS 0.60fF $ **FLOATING
C2981 S.n2697 VSUBS 0.12fF $ **FLOATING
C2982 S.t1140 VSUBS 0.02fF
C2983 S.n2698 VSUBS 0.14fF $ **FLOATING
C2984 S.n2700 VSUBS 1.14fF $ **FLOATING
C2985 S.n2701 VSUBS 0.22fF $ **FLOATING
C2986 S.n2702 VSUBS 0.25fF $ **FLOATING
C2987 S.n2703 VSUBS 0.09fF $ **FLOATING
C2988 S.n2704 VSUBS 1.86fF $ **FLOATING
C2989 S.t463 VSUBS 0.02fF
C2990 S.n2705 VSUBS 0.24fF $ **FLOATING
C2991 S.n2706 VSUBS 0.90fF $ **FLOATING
C2992 S.n2707 VSUBS 0.05fF $ **FLOATING
C2993 S.t347 VSUBS 0.02fF
C2994 S.n2708 VSUBS 0.12fF $ **FLOATING
C2995 S.n2709 VSUBS 0.14fF $ **FLOATING
C2996 S.n2711 VSUBS 0.77fF $ **FLOATING
C2997 S.n2712 VSUBS 1.92fF $ **FLOATING
C2998 S.n2713 VSUBS 1.86fF $ **FLOATING
C2999 S.n2714 VSUBS 0.12fF $ **FLOATING
C3000 S.t961 VSUBS 0.02fF
C3001 S.n2715 VSUBS 0.14fF $ **FLOATING
C3002 S.t212 VSUBS 0.02fF
C3003 S.n2717 VSUBS 0.24fF $ **FLOATING
C3004 S.n2718 VSUBS 0.35fF $ **FLOATING
C3005 S.n2719 VSUBS 0.60fF $ **FLOATING
C3006 S.n2720 VSUBS 1.82fF $ **FLOATING
C3007 S.n2721 VSUBS 2.96fF $ **FLOATING
C3008 S.t329 VSUBS 0.02fF
C3009 S.n2722 VSUBS 0.24fF $ **FLOATING
C3010 S.n2723 VSUBS 0.90fF $ **FLOATING
C3011 S.n2724 VSUBS 0.05fF $ **FLOATING
C3012 S.t756 VSUBS 0.02fF
C3013 S.n2725 VSUBS 0.12fF $ **FLOATING
C3014 S.n2726 VSUBS 0.14fF $ **FLOATING
C3015 S.n2728 VSUBS 1.87fF $ **FLOATING
C3016 S.n2729 VSUBS 1.73fF $ **FLOATING
C3017 S.t562 VSUBS 0.02fF
C3018 S.n2730 VSUBS 0.24fF $ **FLOATING
C3019 S.n2731 VSUBS 0.35fF $ **FLOATING
C3020 S.n2732 VSUBS 0.60fF $ **FLOATING
C3021 S.n2733 VSUBS 0.12fF $ **FLOATING
C3022 S.t198 VSUBS 0.02fF
C3023 S.n2734 VSUBS 0.14fF $ **FLOATING
C3024 S.n2736 VSUBS 1.14fF $ **FLOATING
C3025 S.n2737 VSUBS 0.22fF $ **FLOATING
C3026 S.n2738 VSUBS 0.25fF $ **FLOATING
C3027 S.n2739 VSUBS 0.09fF $ **FLOATING
C3028 S.n2740 VSUBS 2.41fF $ **FLOATING
C3029 S.t675 VSUBS 0.02fF
C3030 S.n2741 VSUBS 0.24fF $ **FLOATING
C3031 S.n2742 VSUBS 0.90fF $ **FLOATING
C3032 S.n2743 VSUBS 0.05fF $ **FLOATING
C3033 S.t579 VSUBS 0.02fF
C3034 S.n2744 VSUBS 0.12fF $ **FLOATING
C3035 S.n2745 VSUBS 0.14fF $ **FLOATING
C3036 S.n2747 VSUBS 1.86fF $ **FLOATING
C3037 S.n2748 VSUBS 0.47fF $ **FLOATING
C3038 S.n2749 VSUBS 0.09fF $ **FLOATING
C3039 S.n2750 VSUBS 0.32fF $ **FLOATING
C3040 S.n2751 VSUBS 0.30fF $ **FLOATING
C3041 S.n2752 VSUBS 0.76fF $ **FLOATING
C3042 S.n2753 VSUBS 0.58fF $ **FLOATING
C3043 S.t907 VSUBS 0.02fF
C3044 S.n2754 VSUBS 0.24fF $ **FLOATING
C3045 S.n2755 VSUBS 0.35fF $ **FLOATING
C3046 S.n2756 VSUBS 0.60fF $ **FLOATING
C3047 S.n2757 VSUBS 0.12fF $ **FLOATING
C3048 S.t547 VSUBS 0.02fF
C3049 S.n2758 VSUBS 0.14fF $ **FLOATING
C3050 S.n2760 VSUBS 2.58fF $ **FLOATING
C3051 S.n2761 VSUBS 2.13fF $ **FLOATING
C3052 S.t1018 VSUBS 0.02fF
C3053 S.n2762 VSUBS 0.24fF $ **FLOATING
C3054 S.n2763 VSUBS 0.90fF $ **FLOATING
C3055 S.n2764 VSUBS 0.05fF $ **FLOATING
C3056 S.t925 VSUBS 0.02fF
C3057 S.n2765 VSUBS 0.12fF $ **FLOATING
C3058 S.n2766 VSUBS 0.14fF $ **FLOATING
C3059 S.n2768 VSUBS 0.77fF $ **FLOATING
C3060 S.n2769 VSUBS 2.27fF $ **FLOATING
C3061 S.n2770 VSUBS 1.86fF $ **FLOATING
C3062 S.n2771 VSUBS 0.12fF $ **FLOATING
C3063 S.t891 VSUBS 0.02fF
C3064 S.n2772 VSUBS 0.14fF $ **FLOATING
C3065 S.t141 VSUBS 0.02fF
C3066 S.n2774 VSUBS 0.24fF $ **FLOATING
C3067 S.n2775 VSUBS 0.35fF $ **FLOATING
C3068 S.n2776 VSUBS 0.60fF $ **FLOATING
C3069 S.n2777 VSUBS 1.37fF $ **FLOATING
C3070 S.n2778 VSUBS 0.70fF $ **FLOATING
C3071 S.n2779 VSUBS 1.13fF $ **FLOATING
C3072 S.n2780 VSUBS 0.35fF $ **FLOATING
C3073 S.n2781 VSUBS 2.00fF $ **FLOATING
C3074 S.t257 VSUBS 0.02fF
C3075 S.n2782 VSUBS 0.24fF $ **FLOATING
C3076 S.n2783 VSUBS 0.90fF $ **FLOATING
C3077 S.n2784 VSUBS 0.05fF $ **FLOATING
C3078 S.t169 VSUBS 0.02fF
C3079 S.n2785 VSUBS 0.12fF $ **FLOATING
C3080 S.n2786 VSUBS 0.14fF $ **FLOATING
C3081 S.n2788 VSUBS 1.87fF $ **FLOATING
C3082 S.n2789 VSUBS 1.86fF $ **FLOATING
C3083 S.t500 VSUBS 0.02fF
C3084 S.n2790 VSUBS 0.24fF $ **FLOATING
C3085 S.n2791 VSUBS 0.35fF $ **FLOATING
C3086 S.n2792 VSUBS 0.60fF $ **FLOATING
C3087 S.n2793 VSUBS 0.12fF $ **FLOATING
C3088 S.t185 VSUBS 0.02fF
C3089 S.n2794 VSUBS 0.14fF $ **FLOATING
C3090 S.n2796 VSUBS 1.14fF $ **FLOATING
C3091 S.n2797 VSUBS 0.22fF $ **FLOATING
C3092 S.n2798 VSUBS 0.25fF $ **FLOATING
C3093 S.n2799 VSUBS 0.09fF $ **FLOATING
C3094 S.n2800 VSUBS 1.86fF $ **FLOATING
C3095 S.t607 VSUBS 0.02fF
C3096 S.n2801 VSUBS 0.24fF $ **FLOATING
C3097 S.n2802 VSUBS 0.90fF $ **FLOATING
C3098 S.n2803 VSUBS 0.05fF $ **FLOATING
C3099 S.t516 VSUBS 0.02fF
C3100 S.n2804 VSUBS 0.12fF $ **FLOATING
C3101 S.n2805 VSUBS 0.14fF $ **FLOATING
C3102 S.n2807 VSUBS 14.09fF $ **FLOATING
C3103 S.n2808 VSUBS 1.86fF $ **FLOATING
C3104 S.n2809 VSUBS 2.64fF $ **FLOATING
C3105 S.t213 VSUBS 0.02fF
C3106 S.n2810 VSUBS 0.24fF $ **FLOATING
C3107 S.n2811 VSUBS 0.35fF $ **FLOATING
C3108 S.n2812 VSUBS 0.60fF $ **FLOATING
C3109 S.n2813 VSUBS 0.12fF $ **FLOATING
C3110 S.t297 VSUBS 0.02fF
C3111 S.n2814 VSUBS 0.14fF $ **FLOATING
C3112 S.n2816 VSUBS 2.77fF $ **FLOATING
C3113 S.n2817 VSUBS 2.27fF $ **FLOATING
C3114 S.t677 VSUBS 0.02fF
C3115 S.n2818 VSUBS 0.12fF $ **FLOATING
C3116 S.n2819 VSUBS 0.14fF $ **FLOATING
C3117 S.t586 VSUBS 0.02fF
C3118 S.n2821 VSUBS 0.24fF $ **FLOATING
C3119 S.n2822 VSUBS 0.90fF $ **FLOATING
C3120 S.n2823 VSUBS 0.05fF $ **FLOATING
C3121 S.n2824 VSUBS 2.70fF $ **FLOATING
C3122 S.n2825 VSUBS 1.58fF $ **FLOATING
C3123 S.n2826 VSUBS 0.12fF $ **FLOATING
C3124 S.t972 VSUBS 0.02fF
C3125 S.n2827 VSUBS 0.14fF $ **FLOATING
C3126 S.t337 VSUBS 0.02fF
C3127 S.n2829 VSUBS 0.24fF $ **FLOATING
C3128 S.n2830 VSUBS 0.35fF $ **FLOATING
C3129 S.n2831 VSUBS 0.60fF $ **FLOATING
C3130 S.n2832 VSUBS 0.07fF $ **FLOATING
C3131 S.n2833 VSUBS 0.01fF $ **FLOATING
C3132 S.n2834 VSUBS 0.23fF $ **FLOATING
C3133 S.n2835 VSUBS 1.15fF $ **FLOATING
C3134 S.n2836 VSUBS 1.33fF $ **FLOATING
C3135 S.n2837 VSUBS 2.27fF $ **FLOATING
C3136 S.t258 VSUBS 0.02fF
C3137 S.n2838 VSUBS 0.12fF $ **FLOATING
C3138 S.n2839 VSUBS 0.14fF $ **FLOATING
C3139 S.t952 VSUBS 0.02fF
C3140 S.n2841 VSUBS 0.24fF $ **FLOATING
C3141 S.n2842 VSUBS 0.90fF $ **FLOATING
C3142 S.n2843 VSUBS 0.05fF $ **FLOATING
C3143 S.t168 VSUBS 32.33fF
C3144 S.t932 VSUBS 0.02fF
C3145 S.n2844 VSUBS 0.24fF $ **FLOATING
C3146 S.n2845 VSUBS 0.90fF $ **FLOATING
C3147 S.n2846 VSUBS 0.05fF $ **FLOATING
C3148 S.t1022 VSUBS 0.02fF
C3149 S.n2847 VSUBS 0.12fF $ **FLOATING
C3150 S.n2848 VSUBS 0.14fF $ **FLOATING
C3151 S.n2850 VSUBS 0.12fF $ **FLOATING
C3152 S.t640 VSUBS 0.02fF
C3153 S.n2851 VSUBS 0.14fF $ **FLOATING
C3154 S.n2853 VSUBS 5.11fF $ **FLOATING
C3155 S.n2854 VSUBS 5.38fF $ **FLOATING
C3156 S.t1013 VSUBS 0.02fF
C3157 S.n2855 VSUBS 0.12fF $ **FLOATING
C3158 S.n2856 VSUBS 0.14fF $ **FLOATING
C3159 S.t920 VSUBS 0.02fF
C3160 S.n2858 VSUBS 0.24fF $ **FLOATING
C3161 S.n2859 VSUBS 0.90fF $ **FLOATING
C3162 S.n2860 VSUBS 0.05fF $ **FLOATING
C3163 S.t154 VSUBS 31.95fF
C3164 S.t480 VSUBS 0.02fF
C3165 S.n2861 VSUBS 0.01fF $ **FLOATING
C3166 S.n2862 VSUBS 0.25fF $ **FLOATING
C3167 S.t851 VSUBS 0.02fF
C3168 S.n2864 VSUBS 1.18fF $ **FLOATING
C3169 S.n2865 VSUBS 0.05fF $ **FLOATING
C3170 S.t715 VSUBS 0.02fF
C3171 S.n2866 VSUBS 0.63fF $ **FLOATING
C3172 S.n2867 VSUBS 0.60fF $ **FLOATING
C3173 S.n2868 VSUBS 8.88fF $ **FLOATING
C3174 S.n2869 VSUBS 8.88fF $ **FLOATING
C3175 S.n2870 VSUBS 0.59fF $ **FLOATING
C3176 S.n2871 VSUBS 0.21fF $ **FLOATING
C3177 S.n2872 VSUBS 0.59fF $ **FLOATING
C3178 S.n2873 VSUBS 2.55fF $ **FLOATING
C3179 S.n2874 VSUBS 0.28fF $ **FLOATING
C3180 S.t107 VSUBS 14.53fF
C3181 S.n2875 VSUBS 15.80fF $ **FLOATING
C3182 S.n2876 VSUBS 0.76fF $ **FLOATING
C3183 S.n2877 VSUBS 0.27fF $ **FLOATING
C3184 S.n2878 VSUBS 3.96fF $ **FLOATING
C3185 S.n2879 VSUBS 1.34fF $ **FLOATING
C3186 S.n2880 VSUBS 0.01fF $ **FLOATING
C3187 S.n2881 VSUBS 0.02fF $ **FLOATING
C3188 S.n2882 VSUBS 0.03fF $ **FLOATING
C3189 S.n2883 VSUBS 0.04fF $ **FLOATING
C3190 S.n2884 VSUBS 0.17fF $ **FLOATING
C3191 S.n2885 VSUBS 0.01fF $ **FLOATING
C3192 S.n2886 VSUBS 0.02fF $ **FLOATING
C3193 S.n2887 VSUBS 0.01fF $ **FLOATING
C3194 S.n2888 VSUBS 0.01fF $ **FLOATING
C3195 S.n2889 VSUBS 0.01fF $ **FLOATING
C3196 S.n2890 VSUBS 0.01fF $ **FLOATING
C3197 S.n2891 VSUBS 0.01fF $ **FLOATING
C3198 S.n2892 VSUBS 0.01fF $ **FLOATING
C3199 S.n2893 VSUBS 0.02fF $ **FLOATING
C3200 S.n2894 VSUBS 0.05fF $ **FLOATING
C3201 S.n2895 VSUBS 0.04fF $ **FLOATING
C3202 S.n2896 VSUBS 0.11fF $ **FLOATING
C3203 S.n2897 VSUBS 0.37fF $ **FLOATING
C3204 S.n2898 VSUBS 0.20fF $ **FLOATING
C3205 S.n2899 VSUBS 4.34fF $ **FLOATING
C3206 S.n2900 VSUBS 0.24fF $ **FLOATING
C3207 S.n2901 VSUBS 1.48fF $ **FLOATING
C3208 S.n2902 VSUBS 1.29fF $ **FLOATING
C3209 S.n2903 VSUBS 0.27fF $ **FLOATING
C3210 S.n2904 VSUBS 0.25fF $ **FLOATING
C3211 S.n2905 VSUBS 0.09fF $ **FLOATING
C3212 S.n2906 VSUBS 0.21fF $ **FLOATING
C3213 S.n2907 VSUBS 0.91fF $ **FLOATING
C3214 S.n2908 VSUBS 0.44fF $ **FLOATING
C3215 S.n2909 VSUBS 1.86fF $ **FLOATING
C3216 S.n2910 VSUBS 0.12fF $ **FLOATING
C3217 S.t618 VSUBS 0.02fF
C3218 S.n2911 VSUBS 0.14fF $ **FLOATING
C3219 S.t979 VSUBS 0.02fF
C3220 S.n2913 VSUBS 0.24fF $ **FLOATING
C3221 S.n2914 VSUBS 0.35fF $ **FLOATING
C3222 S.n2915 VSUBS 0.60fF $ **FLOATING
C3223 S.n2916 VSUBS 0.02fF $ **FLOATING
C3224 S.n2917 VSUBS 0.01fF $ **FLOATING
C3225 S.n2918 VSUBS 0.02fF $ **FLOATING
C3226 S.n2919 VSUBS 0.08fF $ **FLOATING
C3227 S.n2920 VSUBS 0.06fF $ **FLOATING
C3228 S.n2921 VSUBS 0.03fF $ **FLOATING
C3229 S.n2922 VSUBS 0.03fF $ **FLOATING
C3230 S.n2923 VSUBS 0.99fF $ **FLOATING
C3231 S.n2924 VSUBS 0.35fF $ **FLOATING
C3232 S.n2925 VSUBS 1.85fF $ **FLOATING
C3233 S.n2926 VSUBS 1.97fF $ **FLOATING
C3234 S.t1112 VSUBS 0.02fF
C3235 S.n2927 VSUBS 0.24fF $ **FLOATING
C3236 S.n2928 VSUBS 0.90fF $ **FLOATING
C3237 S.n2929 VSUBS 0.05fF $ **FLOATING
C3238 S.t999 VSUBS 0.02fF
C3239 S.n2930 VSUBS 0.12fF $ **FLOATING
C3240 S.n2931 VSUBS 0.14fF $ **FLOATING
C3241 S.n2933 VSUBS 1.87fF $ **FLOATING
C3242 S.n2934 VSUBS 0.07fF $ **FLOATING
C3243 S.n2935 VSUBS 0.04fF $ **FLOATING
C3244 S.n2936 VSUBS 0.05fF $ **FLOATING
C3245 S.n2937 VSUBS 0.86fF $ **FLOATING
C3246 S.n2938 VSUBS 0.01fF $ **FLOATING
C3247 S.n2939 VSUBS 0.01fF $ **FLOATING
C3248 S.n2940 VSUBS 0.01fF $ **FLOATING
C3249 S.n2941 VSUBS 0.07fF $ **FLOATING
C3250 S.n2942 VSUBS 0.68fF $ **FLOATING
C3251 S.n2943 VSUBS 0.71fF $ **FLOATING
C3252 S.t823 VSUBS 0.02fF
C3253 S.n2944 VSUBS 0.24fF $ **FLOATING
C3254 S.n2945 VSUBS 0.35fF $ **FLOATING
C3255 S.n2946 VSUBS 0.60fF $ **FLOATING
C3256 S.n2947 VSUBS 0.12fF $ **FLOATING
C3257 S.t466 VSUBS 0.02fF
C3258 S.n2948 VSUBS 0.14fF $ **FLOATING
C3259 S.n2950 VSUBS 0.69fF $ **FLOATING
C3260 S.n2951 VSUBS 0.22fF $ **FLOATING
C3261 S.n2952 VSUBS 0.22fF $ **FLOATING
C3262 S.n2953 VSUBS 0.69fF $ **FLOATING
C3263 S.n2954 VSUBS 1.14fF $ **FLOATING
C3264 S.n2955 VSUBS 0.22fF $ **FLOATING
C3265 S.n2956 VSUBS 0.25fF $ **FLOATING
C3266 S.n2957 VSUBS 0.09fF $ **FLOATING
C3267 S.n2958 VSUBS 2.29fF $ **FLOATING
C3268 S.t940 VSUBS 0.02fF
C3269 S.n2959 VSUBS 0.24fF $ **FLOATING
C3270 S.n2960 VSUBS 0.90fF $ **FLOATING
C3271 S.n2961 VSUBS 0.05fF $ **FLOATING
C3272 S.t847 VSUBS 0.02fF
C3273 S.n2962 VSUBS 0.12fF $ **FLOATING
C3274 S.n2963 VSUBS 0.14fF $ **FLOATING
C3275 S.n2965 VSUBS 1.86fF $ **FLOATING
C3276 S.n2966 VSUBS 0.45fF $ **FLOATING
C3277 S.n2967 VSUBS 0.22fF $ **FLOATING
C3278 S.n2968 VSUBS 0.38fF $ **FLOATING
C3279 S.n2969 VSUBS 0.16fF $ **FLOATING
C3280 S.n2970 VSUBS 0.28fF $ **FLOATING
C3281 S.n2971 VSUBS 0.21fF $ **FLOATING
C3282 S.n2972 VSUBS 0.30fF $ **FLOATING
C3283 S.n2973 VSUBS 0.41fF $ **FLOATING
C3284 S.n2974 VSUBS 0.20fF $ **FLOATING
C3285 S.t34 VSUBS 0.02fF
C3286 S.n2975 VSUBS 0.24fF $ **FLOATING
C3287 S.n2976 VSUBS 0.35fF $ **FLOATING
C3288 S.n2977 VSUBS 0.60fF $ **FLOATING
C3289 S.n2978 VSUBS 0.12fF $ **FLOATING
C3290 S.t806 VSUBS 0.02fF
C3291 S.n2979 VSUBS 0.14fF $ **FLOATING
C3292 S.n2981 VSUBS 0.04fF $ **FLOATING
C3293 S.n2982 VSUBS 0.03fF $ **FLOATING
C3294 S.n2983 VSUBS 0.03fF $ **FLOATING
C3295 S.n2984 VSUBS 0.10fF $ **FLOATING
C3296 S.n2985 VSUBS 0.36fF $ **FLOATING
C3297 S.n2986 VSUBS 0.37fF $ **FLOATING
C3298 S.n2987 VSUBS 0.10fF $ **FLOATING
C3299 S.n2988 VSUBS 0.12fF $ **FLOATING
C3300 S.n2989 VSUBS 0.07fF $ **FLOATING
C3301 S.n2990 VSUBS 0.12fF $ **FLOATING
C3302 S.n2991 VSUBS 0.18fF $ **FLOATING
C3303 S.n2992 VSUBS 3.95fF $ **FLOATING
C3304 S.t180 VSUBS 0.02fF
C3305 S.n2993 VSUBS 0.24fF $ **FLOATING
C3306 S.n2994 VSUBS 0.90fF $ **FLOATING
C3307 S.n2995 VSUBS 0.05fF $ **FLOATING
C3308 S.t70 VSUBS 0.02fF
C3309 S.n2996 VSUBS 0.12fF $ **FLOATING
C3310 S.n2997 VSUBS 0.14fF $ **FLOATING
C3311 S.n2999 VSUBS 0.25fF $ **FLOATING
C3312 S.n3000 VSUBS 0.09fF $ **FLOATING
C3313 S.n3001 VSUBS 0.21fF $ **FLOATING
C3314 S.n3002 VSUBS 1.27fF $ **FLOATING
C3315 S.n3003 VSUBS 0.52fF $ **FLOATING
C3316 S.n3004 VSUBS 1.86fF $ **FLOATING
C3317 S.n3005 VSUBS 0.12fF $ **FLOATING
C3318 S.t15 VSUBS 0.02fF
C3319 S.n3006 VSUBS 0.14fF $ **FLOATING
C3320 S.t405 VSUBS 0.02fF
C3321 S.n3008 VSUBS 0.24fF $ **FLOATING
C3322 S.n3009 VSUBS 0.35fF $ **FLOATING
C3323 S.n3010 VSUBS 0.60fF $ **FLOATING
C3324 S.n3011 VSUBS 1.56fF $ **FLOATING
C3325 S.n3012 VSUBS 2.42fF $ **FLOATING
C3326 S.t530 VSUBS 0.02fF
C3327 S.n3013 VSUBS 0.24fF $ **FLOATING
C3328 S.n3014 VSUBS 0.90fF $ **FLOATING
C3329 S.n3015 VSUBS 0.05fF $ **FLOATING
C3330 S.t429 VSUBS 0.02fF
C3331 S.n3016 VSUBS 0.12fF $ **FLOATING
C3332 S.n3017 VSUBS 0.14fF $ **FLOATING
C3333 S.n3019 VSUBS 1.87fF $ **FLOATING
C3334 S.n3020 VSUBS 0.06fF $ **FLOATING
C3335 S.n3021 VSUBS 0.03fF $ **FLOATING
C3336 S.n3022 VSUBS 0.03fF $ **FLOATING
C3337 S.n3023 VSUBS 0.98fF $ **FLOATING
C3338 S.n3024 VSUBS 0.02fF $ **FLOATING
C3339 S.n3025 VSUBS 0.01fF $ **FLOATING
C3340 S.n3026 VSUBS 0.02fF $ **FLOATING
C3341 S.n3027 VSUBS 0.08fF $ **FLOATING
C3342 S.n3028 VSUBS 0.36fF $ **FLOATING
C3343 S.n3029 VSUBS 1.83fF $ **FLOATING
C3344 S.t747 VSUBS 0.02fF
C3345 S.n3030 VSUBS 0.24fF $ **FLOATING
C3346 S.n3031 VSUBS 0.35fF $ **FLOATING
C3347 S.n3032 VSUBS 0.60fF $ **FLOATING
C3348 S.n3033 VSUBS 0.12fF $ **FLOATING
C3349 S.t389 VSUBS 0.02fF
C3350 S.n3034 VSUBS 0.14fF $ **FLOATING
C3351 S.n3036 VSUBS 0.69fF $ **FLOATING
C3352 S.n3037 VSUBS 0.22fF $ **FLOATING
C3353 S.n3038 VSUBS 0.22fF $ **FLOATING
C3354 S.n3039 VSUBS 0.69fF $ **FLOATING
C3355 S.n3040 VSUBS 1.14fF $ **FLOATING
C3356 S.n3041 VSUBS 0.22fF $ **FLOATING
C3357 S.n3042 VSUBS 0.25fF $ **FLOATING
C3358 S.n3043 VSUBS 0.09fF $ **FLOATING
C3359 S.n3044 VSUBS 1.86fF $ **FLOATING
C3360 S.t873 VSUBS 0.02fF
C3361 S.n3045 VSUBS 0.24fF $ **FLOATING
C3362 S.n3046 VSUBS 0.90fF $ **FLOATING
C3363 S.n3047 VSUBS 0.05fF $ **FLOATING
C3364 S.t770 VSUBS 0.02fF
C3365 S.n3048 VSUBS 0.12fF $ **FLOATING
C3366 S.n3049 VSUBS 0.14fF $ **FLOATING
C3367 S.n3051 VSUBS 14.09fF $ **FLOATING
C3368 S.n3052 VSUBS 1.70fF $ **FLOATING
C3369 S.n3053 VSUBS 3.01fF $ **FLOATING
C3370 S.t585 VSUBS 0.02fF
C3371 S.n3054 VSUBS 0.24fF $ **FLOATING
C3372 S.n3055 VSUBS 0.35fF $ **FLOATING
C3373 S.n3056 VSUBS 0.60fF $ **FLOATING
C3374 S.n3057 VSUBS 0.12fF $ **FLOATING
C3375 S.t220 VSUBS 0.02fF
C3376 S.n3058 VSUBS 0.14fF $ **FLOATING
C3377 S.n3060 VSUBS 0.31fF $ **FLOATING
C3378 S.n3061 VSUBS 0.22fF $ **FLOATING
C3379 S.n3062 VSUBS 0.65fF $ **FLOATING
C3380 S.n3063 VSUBS 0.94fF $ **FLOATING
C3381 S.n3064 VSUBS 0.22fF $ **FLOATING
C3382 S.n3065 VSUBS 0.20fF $ **FLOATING
C3383 S.n3066 VSUBS 0.20fF $ **FLOATING
C3384 S.n3067 VSUBS 0.06fF $ **FLOATING
C3385 S.n3068 VSUBS 0.09fF $ **FLOATING
C3386 S.n3069 VSUBS 0.09fF $ **FLOATING
C3387 S.n3070 VSUBS 1.97fF $ **FLOATING
C3388 S.t600 VSUBS 0.02fF
C3389 S.n3071 VSUBS 0.12fF $ **FLOATING
C3390 S.n3072 VSUBS 0.14fF $ **FLOATING
C3391 S.t704 VSUBS 0.02fF
C3392 S.n3074 VSUBS 0.24fF $ **FLOATING
C3393 S.n3075 VSUBS 0.90fF $ **FLOATING
C3394 S.n3076 VSUBS 0.05fF $ **FLOATING
C3395 S.n3077 VSUBS 1.86fF $ **FLOATING
C3396 S.n3078 VSUBS 0.12fF $ **FLOATING
C3397 S.t1031 VSUBS 0.02fF
C3398 S.n3079 VSUBS 0.14fF $ **FLOATING
C3399 S.t249 VSUBS 0.02fF
C3400 S.n3081 VSUBS 0.12fF $ **FLOATING
C3401 S.n3082 VSUBS 0.14fF $ **FLOATING
C3402 S.t362 VSUBS 0.02fF
C3403 S.n3084 VSUBS 0.24fF $ **FLOATING
C3404 S.n3085 VSUBS 0.90fF $ **FLOATING
C3405 S.n3086 VSUBS 0.05fF $ **FLOATING
C3406 S.t229 VSUBS 0.02fF
C3407 S.n3087 VSUBS 0.24fF $ **FLOATING
C3408 S.n3088 VSUBS 0.35fF $ **FLOATING
C3409 S.n3089 VSUBS 0.60fF $ **FLOATING
C3410 S.n3090 VSUBS 0.31fF $ **FLOATING
C3411 S.n3091 VSUBS 1.08fF $ **FLOATING
C3412 S.n3092 VSUBS 0.15fF $ **FLOATING
C3413 S.n3093 VSUBS 2.08fF $ **FLOATING
C3414 S.n3094 VSUBS 2.91fF $ **FLOATING
C3415 S.n3095 VSUBS 1.86fF $ **FLOATING
C3416 S.n3096 VSUBS 0.12fF $ **FLOATING
C3417 S.t733 VSUBS 0.02fF
C3418 S.n3097 VSUBS 0.14fF $ **FLOATING
C3419 S.t633 VSUBS 0.02fF
C3420 S.n3099 VSUBS 0.24fF $ **FLOATING
C3421 S.n3100 VSUBS 0.35fF $ **FLOATING
C3422 S.n3101 VSUBS 0.60fF $ **FLOATING
C3423 S.n3102 VSUBS 0.91fF $ **FLOATING
C3424 S.n3103 VSUBS 0.31fF $ **FLOATING
C3425 S.n3104 VSUBS 0.91fF $ **FLOATING
C3426 S.n3105 VSUBS 1.08fF $ **FLOATING
C3427 S.n3106 VSUBS 0.15fF $ **FLOATING
C3428 S.n3107 VSUBS 4.90fF $ **FLOATING
C3429 S.t47 VSUBS 0.02fF
C3430 S.n3108 VSUBS 0.12fF $ **FLOATING
C3431 S.n3109 VSUBS 0.14fF $ **FLOATING
C3432 S.t1008 VSUBS 0.02fF
C3433 S.n3111 VSUBS 0.24fF $ **FLOATING
C3434 S.n3112 VSUBS 0.90fF $ **FLOATING
C3435 S.n3113 VSUBS 0.05fF $ **FLOATING
C3436 S.n3114 VSUBS 1.86fF $ **FLOATING
C3437 S.n3115 VSUBS 2.64fF $ **FLOATING
C3438 S.t983 VSUBS 0.02fF
C3439 S.n3116 VSUBS 0.24fF $ **FLOATING
C3440 S.n3117 VSUBS 0.35fF $ **FLOATING
C3441 S.n3118 VSUBS 0.60fF $ **FLOATING
C3442 S.n3119 VSUBS 0.12fF $ **FLOATING
C3443 S.t1067 VSUBS 0.02fF
C3444 S.n3120 VSUBS 0.14fF $ **FLOATING
C3445 S.n3122 VSUBS 1.86fF $ **FLOATING
C3446 S.n3123 VSUBS 2.64fF $ **FLOATING
C3447 S.t993 VSUBS 0.02fF
C3448 S.n3124 VSUBS 0.24fF $ **FLOATING
C3449 S.n3125 VSUBS 0.35fF $ **FLOATING
C3450 S.n3126 VSUBS 0.60fF $ **FLOATING
C3451 S.t252 VSUBS 0.02fF
C3452 S.n3127 VSUBS 0.24fF $ **FLOATING
C3453 S.n3128 VSUBS 0.90fF $ **FLOATING
C3454 S.n3129 VSUBS 0.05fF $ **FLOATING
C3455 S.t367 VSUBS 0.02fF
C3456 S.n3130 VSUBS 0.12fF $ **FLOATING
C3457 S.n3131 VSUBS 0.14fF $ **FLOATING
C3458 S.n3133 VSUBS 0.12fF $ **FLOATING
C3459 S.t1085 VSUBS 0.02fF
C3460 S.n3134 VSUBS 0.14fF $ **FLOATING
C3461 S.n3136 VSUBS 2.27fF $ **FLOATING
C3462 S.n3137 VSUBS 2.91fF $ **FLOATING
C3463 S.n3138 VSUBS 5.10fF $ **FLOATING
C3464 S.t349 VSUBS 0.02fF
C3465 S.n3139 VSUBS 0.12fF $ **FLOATING
C3466 S.n3140 VSUBS 0.14fF $ **FLOATING
C3467 S.t242 VSUBS 0.02fF
C3468 S.n3142 VSUBS 0.24fF $ **FLOATING
C3469 S.n3143 VSUBS 0.90fF $ **FLOATING
C3470 S.n3144 VSUBS 0.05fF $ **FLOATING
C3471 S.n3145 VSUBS 1.86fF $ **FLOATING
C3472 S.n3146 VSUBS 2.64fF $ **FLOATING
C3473 S.t222 VSUBS 0.02fF
C3474 S.n3147 VSUBS 0.24fF $ **FLOATING
C3475 S.n3148 VSUBS 0.35fF $ **FLOATING
C3476 S.n3149 VSUBS 0.60fF $ **FLOATING
C3477 S.n3150 VSUBS 0.12fF $ **FLOATING
C3478 S.t306 VSUBS 0.02fF
C3479 S.n3151 VSUBS 0.14fF $ **FLOATING
C3480 S.n3153 VSUBS 5.11fF $ **FLOATING
C3481 S.t687 VSUBS 0.02fF
C3482 S.n3154 VSUBS 0.12fF $ **FLOATING
C3483 S.n3155 VSUBS 0.14fF $ **FLOATING
C3484 S.t595 VSUBS 0.02fF
C3485 S.n3157 VSUBS 0.24fF $ **FLOATING
C3486 S.n3158 VSUBS 0.90fF $ **FLOATING
C3487 S.n3159 VSUBS 0.05fF $ **FLOATING
C3488 S.n3160 VSUBS 1.86fF $ **FLOATING
C3489 S.n3161 VSUBS 2.64fF $ **FLOATING
C3490 S.t572 VSUBS 0.02fF
C3491 S.n3162 VSUBS 0.24fF $ **FLOATING
C3492 S.n3163 VSUBS 0.35fF $ **FLOATING
C3493 S.n3164 VSUBS 0.60fF $ **FLOATING
C3494 S.n3165 VSUBS 0.12fF $ **FLOATING
C3495 S.t653 VSUBS 0.02fF
C3496 S.n3166 VSUBS 0.14fF $ **FLOATING
C3497 S.n3168 VSUBS 4.84fF $ **FLOATING
C3498 S.t1032 VSUBS 0.02fF
C3499 S.n3169 VSUBS 0.12fF $ **FLOATING
C3500 S.n3170 VSUBS 0.14fF $ **FLOATING
C3501 S.t941 VSUBS 0.02fF
C3502 S.n3172 VSUBS 0.24fF $ **FLOATING
C3503 S.n3173 VSUBS 0.90fF $ **FLOATING
C3504 S.n3174 VSUBS 0.05fF $ **FLOATING
C3505 S.n3175 VSUBS 1.86fF $ **FLOATING
C3506 S.n3176 VSUBS 2.64fF $ **FLOATING
C3507 S.t919 VSUBS 0.02fF
C3508 S.n3177 VSUBS 0.24fF $ **FLOATING
C3509 S.n3178 VSUBS 0.35fF $ **FLOATING
C3510 S.n3179 VSUBS 0.60fF $ **FLOATING
C3511 S.n3180 VSUBS 0.12fF $ **FLOATING
C3512 S.t997 VSUBS 0.02fF
C3513 S.n3181 VSUBS 0.14fF $ **FLOATING
C3514 S.n3183 VSUBS 1.86fF $ **FLOATING
C3515 S.n3184 VSUBS 2.65fF $ **FLOATING
C3516 S.t929 VSUBS 0.02fF
C3517 S.n3185 VSUBS 0.24fF $ **FLOATING
C3518 S.n3186 VSUBS 0.35fF $ **FLOATING
C3519 S.n3187 VSUBS 0.60fF $ **FLOATING
C3520 S.t850 VSUBS 0.02fF
C3521 S.n3188 VSUBS 1.20fF $ **FLOATING
C3522 S.n3189 VSUBS 0.60fF $ **FLOATING
C3523 S.n3190 VSUBS 0.35fF $ **FLOATING
C3524 S.n3191 VSUBS 0.62fF $ **FLOATING
C3525 S.n3192 VSUBS 1.14fF $ **FLOATING
C3526 S.n3193 VSUBS 2.15fF $ **FLOATING
C3527 S.n3194 VSUBS 0.59fF $ **FLOATING
C3528 S.n3195 VSUBS 0.01fF $ **FLOATING
C3529 S.n3196 VSUBS 0.96fF $ **FLOATING
C3530 S.t72 VSUBS 14.53fF
C3531 S.n3197 VSUBS 14.40fF $ **FLOATING
C3532 S.n3199 VSUBS 0.37fF $ **FLOATING
C3533 S.n3200 VSUBS 0.23fF $ **FLOATING
C3534 S.n3201 VSUBS 2.87fF $ **FLOATING
C3535 S.n3202 VSUBS 2.43fF $ **FLOATING
C3536 S.n3203 VSUBS 1.94fF $ **FLOATING
C3537 S.n3204 VSUBS 3.89fF $ **FLOATING
C3538 S.n3205 VSUBS 0.25fF $ **FLOATING
C3539 S.n3206 VSUBS 0.01fF $ **FLOATING
C3540 S.t492 VSUBS 0.02fF
C3541 S.n3207 VSUBS 0.25fF $ **FLOATING
C3542 S.t964 VSUBS 0.02fF
C3543 S.n3208 VSUBS 0.94fF $ **FLOATING
C3544 S.n3209 VSUBS 0.70fF $ **FLOATING
C3545 S.n3210 VSUBS 0.77fF $ **FLOATING
C3546 S.n3211 VSUBS 1.91fF $ **FLOATING
C3547 S.n3212 VSUBS 1.86fF $ **FLOATING
C3548 S.n3213 VSUBS 0.12fF $ **FLOATING
C3549 S.t884 VSUBS 0.02fF
C3550 S.n3214 VSUBS 0.14fF $ **FLOATING
C3551 S.t73 VSUBS 0.02fF
C3552 S.n3216 VSUBS 0.24fF $ **FLOATING
C3553 S.n3217 VSUBS 0.35fF $ **FLOATING
C3554 S.n3218 VSUBS 0.60fF $ **FLOATING
C3555 S.n3219 VSUBS 1.50fF $ **FLOATING
C3556 S.n3220 VSUBS 2.96fF $ **FLOATING
C3557 S.t201 VSUBS 0.02fF
C3558 S.n3221 VSUBS 0.24fF $ **FLOATING
C3559 S.n3222 VSUBS 0.90fF $ **FLOATING
C3560 S.n3223 VSUBS 0.05fF $ **FLOATING
C3561 S.t96 VSUBS 0.02fF
C3562 S.n3224 VSUBS 0.12fF $ **FLOATING
C3563 S.n3225 VSUBS 0.14fF $ **FLOATING
C3564 S.n3227 VSUBS 1.87fF $ **FLOATING
C3565 S.n3228 VSUBS 1.73fF $ **FLOATING
C3566 S.t1060 VSUBS 0.02fF
C3567 S.n3229 VSUBS 0.24fF $ **FLOATING
C3568 S.n3230 VSUBS 0.35fF $ **FLOATING
C3569 S.n3231 VSUBS 0.60fF $ **FLOATING
C3570 S.n3232 VSUBS 0.12fF $ **FLOATING
C3571 S.t709 VSUBS 0.02fF
C3572 S.n3233 VSUBS 0.14fF $ **FLOATING
C3573 S.n3235 VSUBS 1.14fF $ **FLOATING
C3574 S.n3236 VSUBS 0.22fF $ **FLOATING
C3575 S.n3237 VSUBS 0.25fF $ **FLOATING
C3576 S.n3238 VSUBS 0.09fF $ **FLOATING
C3577 S.n3239 VSUBS 2.41fF $ **FLOATING
C3578 S.t83 VSUBS 0.02fF
C3579 S.n3240 VSUBS 0.24fF $ **FLOATING
C3580 S.n3241 VSUBS 0.90fF $ **FLOATING
C3581 S.n3242 VSUBS 0.05fF $ **FLOATING
C3582 S.t510 VSUBS 0.02fF
C3583 S.n3243 VSUBS 0.12fF $ **FLOATING
C3584 S.n3244 VSUBS 0.14fF $ **FLOATING
C3585 S.n3246 VSUBS 1.86fF $ **FLOATING
C3586 S.n3247 VSUBS 0.47fF $ **FLOATING
C3587 S.n3248 VSUBS 0.09fF $ **FLOATING
C3588 S.n3249 VSUBS 0.32fF $ **FLOATING
C3589 S.n3250 VSUBS 0.30fF $ **FLOATING
C3590 S.n3251 VSUBS 0.76fF $ **FLOATING
C3591 S.n3252 VSUBS 0.58fF $ **FLOATING
C3592 S.t301 VSUBS 0.02fF
C3593 S.n3253 VSUBS 0.24fF $ **FLOATING
C3594 S.n3254 VSUBS 0.35fF $ **FLOATING
C3595 S.n3255 VSUBS 0.60fF $ **FLOATING
C3596 S.n3256 VSUBS 0.12fF $ **FLOATING
C3597 S.t1047 VSUBS 0.02fF
C3598 S.n3257 VSUBS 0.14fF $ **FLOATING
C3599 S.n3259 VSUBS 2.58fF $ **FLOATING
C3600 S.n3260 VSUBS 2.13fF $ **FLOATING
C3601 S.t445 VSUBS 0.02fF
C3602 S.n3261 VSUBS 0.24fF $ **FLOATING
C3603 S.n3262 VSUBS 0.90fF $ **FLOATING
C3604 S.n3263 VSUBS 0.05fF $ **FLOATING
C3605 S.t323 VSUBS 0.02fF
C3606 S.n3264 VSUBS 0.12fF $ **FLOATING
C3607 S.n3265 VSUBS 0.14fF $ **FLOATING
C3608 S.n3267 VSUBS 0.77fF $ **FLOATING
C3609 S.n3268 VSUBS 2.27fF $ **FLOATING
C3610 S.n3269 VSUBS 1.86fF $ **FLOATING
C3611 S.n3270 VSUBS 0.12fF $ **FLOATING
C3612 S.t285 VSUBS 0.02fF
C3613 S.n3271 VSUBS 0.14fF $ **FLOATING
C3614 S.t641 VSUBS 0.02fF
C3615 S.n3273 VSUBS 0.24fF $ **FLOATING
C3616 S.n3274 VSUBS 0.35fF $ **FLOATING
C3617 S.n3275 VSUBS 0.60fF $ **FLOATING
C3618 S.n3276 VSUBS 1.37fF $ **FLOATING
C3619 S.n3277 VSUBS 0.70fF $ **FLOATING
C3620 S.n3278 VSUBS 1.13fF $ **FLOATING
C3621 S.n3279 VSUBS 0.35fF $ **FLOATING
C3622 S.n3280 VSUBS 2.00fF $ **FLOATING
C3623 S.t782 VSUBS 0.02fF
C3624 S.n3281 VSUBS 0.24fF $ **FLOATING
C3625 S.n3282 VSUBS 0.90fF $ **FLOATING
C3626 S.n3283 VSUBS 0.05fF $ **FLOATING
C3627 S.t666 VSUBS 0.02fF
C3628 S.n3284 VSUBS 0.12fF $ **FLOATING
C3629 S.n3285 VSUBS 0.14fF $ **FLOATING
C3630 S.n3287 VSUBS 1.87fF $ **FLOATING
C3631 S.n3288 VSUBS 1.86fF $ **FLOATING
C3632 S.t991 VSUBS 0.02fF
C3633 S.n3289 VSUBS 0.24fF $ **FLOATING
C3634 S.n3290 VSUBS 0.35fF $ **FLOATING
C3635 S.n3291 VSUBS 0.60fF $ **FLOATING
C3636 S.n3292 VSUBS 0.12fF $ **FLOATING
C3637 S.t629 VSUBS 0.02fF
C3638 S.n3293 VSUBS 0.14fF $ **FLOATING
C3639 S.n3295 VSUBS 1.14fF $ **FLOATING
C3640 S.n3296 VSUBS 0.22fF $ **FLOATING
C3641 S.n3297 VSUBS 0.25fF $ **FLOATING
C3642 S.n3298 VSUBS 0.09fF $ **FLOATING
C3643 S.n3299 VSUBS 1.86fF $ **FLOATING
C3644 S.t1126 VSUBS 0.02fF
C3645 S.n3300 VSUBS 0.24fF $ **FLOATING
C3646 S.n3301 VSUBS 0.90fF $ **FLOATING
C3647 S.n3302 VSUBS 0.05fF $ **FLOATING
C3648 S.t1014 VSUBS 0.02fF
C3649 S.n3303 VSUBS 0.12fF $ **FLOATING
C3650 S.n3304 VSUBS 0.14fF $ **FLOATING
C3651 S.n3306 VSUBS 14.09fF $ **FLOATING
C3652 S.n3307 VSUBS 1.86fF $ **FLOATING
C3653 S.n3308 VSUBS 2.64fF $ **FLOATING
C3654 S.t236 VSUBS 0.02fF
C3655 S.n3309 VSUBS 0.24fF $ **FLOATING
C3656 S.n3310 VSUBS 0.35fF $ **FLOATING
C3657 S.n3311 VSUBS 0.60fF $ **FLOATING
C3658 S.n3312 VSUBS 0.12fF $ **FLOATING
C3659 S.t316 VSUBS 0.02fF
C3660 S.n3313 VSUBS 0.14fF $ **FLOATING
C3661 S.n3315 VSUBS 2.77fF $ **FLOATING
C3662 S.n3316 VSUBS 2.27fF $ **FLOATING
C3663 S.t700 VSUBS 0.02fF
C3664 S.n3317 VSUBS 0.12fF $ **FLOATING
C3665 S.n3318 VSUBS 0.14fF $ **FLOATING
C3666 S.t603 VSUBS 0.02fF
C3667 S.n3320 VSUBS 0.24fF $ **FLOATING
C3668 S.n3321 VSUBS 0.90fF $ **FLOATING
C3669 S.n3322 VSUBS 0.05fF $ **FLOATING
C3670 S.n3323 VSUBS 1.86fF $ **FLOATING
C3671 S.n3324 VSUBS 2.64fF $ **FLOATING
C3672 S.t583 VSUBS 0.02fF
C3673 S.n3325 VSUBS 0.24fF $ **FLOATING
C3674 S.n3326 VSUBS 0.35fF $ **FLOATING
C3675 S.n3327 VSUBS 0.60fF $ **FLOATING
C3676 S.n3328 VSUBS 0.12fF $ **FLOATING
C3677 S.t662 VSUBS 0.02fF
C3678 S.n3329 VSUBS 0.14fF $ **FLOATING
C3679 S.n3331 VSUBS 2.77fF $ **FLOATING
C3680 S.n3332 VSUBS 2.27fF $ **FLOATING
C3681 S.t1041 VSUBS 0.02fF
C3682 S.n3333 VSUBS 0.12fF $ **FLOATING
C3683 S.n3334 VSUBS 0.14fF $ **FLOATING
C3684 S.t948 VSUBS 0.02fF
C3685 S.n3336 VSUBS 0.24fF $ **FLOATING
C3686 S.n3337 VSUBS 0.90fF $ **FLOATING
C3687 S.n3338 VSUBS 0.05fF $ **FLOATING
C3688 S.n3339 VSUBS 2.70fF $ **FLOATING
C3689 S.n3340 VSUBS 1.58fF $ **FLOATING
C3690 S.n3341 VSUBS 0.12fF $ **FLOATING
C3691 S.t888 VSUBS 0.02fF
C3692 S.n3342 VSUBS 0.14fF $ **FLOATING
C3693 S.t843 VSUBS 0.02fF
C3694 S.n3344 VSUBS 0.24fF $ **FLOATING
C3695 S.n3345 VSUBS 0.90fF $ **FLOATING
C3696 S.n3346 VSUBS 0.05fF $ **FLOATING
C3697 S.t218 VSUBS 0.02fF
C3698 S.n3347 VSUBS 0.24fF $ **FLOATING
C3699 S.n3348 VSUBS 0.35fF $ **FLOATING
C3700 S.n3349 VSUBS 0.60fF $ **FLOATING
C3701 S.n3350 VSUBS 0.07fF $ **FLOATING
C3702 S.n3351 VSUBS 0.01fF $ **FLOATING
C3703 S.n3352 VSUBS 0.23fF $ **FLOATING
C3704 S.n3353 VSUBS 1.15fF $ **FLOATING
C3705 S.n3354 VSUBS 1.33fF $ **FLOATING
C3706 S.n3355 VSUBS 2.27fF $ **FLOATING
C3707 S.t624 VSUBS 0.02fF
C3708 S.n3356 VSUBS 0.12fF $ **FLOATING
C3709 S.n3357 VSUBS 0.14fF $ **FLOATING
C3710 S.t95 VSUBS 32.33fF
C3711 S.t191 VSUBS 0.02fF
C3712 S.n3359 VSUBS 0.24fF $ **FLOATING
C3713 S.n3360 VSUBS 0.90fF $ **FLOATING
C3714 S.n3361 VSUBS 0.05fF $ **FLOATING
C3715 S.t283 VSUBS 0.02fF
C3716 S.n3362 VSUBS 0.12fF $ **FLOATING
C3717 S.n3363 VSUBS 0.14fF $ **FLOATING
C3718 S.n3365 VSUBS 0.12fF $ **FLOATING
C3719 S.t1011 VSUBS 0.02fF
C3720 S.n3366 VSUBS 0.14fF $ **FLOATING
C3721 S.n3368 VSUBS 5.11fF $ **FLOATING
C3722 S.n3369 VSUBS 5.38fF $ **FLOATING
C3723 S.t272 VSUBS 0.02fF
C3724 S.n3370 VSUBS 0.12fF $ **FLOATING
C3725 S.n3371 VSUBS 0.14fF $ **FLOATING
C3726 S.t182 VSUBS 0.02fF
C3727 S.n3373 VSUBS 0.24fF $ **FLOATING
C3728 S.n3374 VSUBS 0.90fF $ **FLOATING
C3729 S.n3375 VSUBS 0.05fF $ **FLOATING
C3730 S.t14 VSUBS 31.95fF
C3731 S.t383 VSUBS 0.02fF
C3732 S.n3376 VSUBS 0.01fF $ **FLOATING
C3733 S.n3377 VSUBS 0.25fF $ **FLOATING
C3734 S.t592 VSUBS 0.02fF
C3735 S.n3379 VSUBS 1.18fF $ **FLOATING
C3736 S.n3380 VSUBS 0.05fF $ **FLOATING
C3737 S.t475 VSUBS 0.02fF
C3738 S.n3381 VSUBS 0.63fF $ **FLOATING
C3739 S.n3382 VSUBS 0.60fF $ **FLOATING
C3740 S.n3383 VSUBS 8.88fF $ **FLOATING
C3741 S.n3384 VSUBS 8.88fF $ **FLOATING
C3742 S.n3385 VSUBS 0.59fF $ **FLOATING
C3743 S.n3386 VSUBS 0.21fF $ **FLOATING
C3744 S.n3387 VSUBS 0.59fF $ **FLOATING
C3745 S.n3388 VSUBS 2.55fF $ **FLOATING
C3746 S.n3389 VSUBS 0.28fF $ **FLOATING
C3747 S.t33 VSUBS 14.53fF
C3748 S.n3390 VSUBS 15.80fF $ **FLOATING
C3749 S.n3391 VSUBS 0.76fF $ **FLOATING
C3750 S.n3392 VSUBS 0.27fF $ **FLOATING
C3751 S.n3393 VSUBS 3.96fF $ **FLOATING
C3752 S.n3394 VSUBS 1.34fF $ **FLOATING
C3753 S.n3395 VSUBS 0.01fF $ **FLOATING
C3754 S.n3396 VSUBS 0.02fF $ **FLOATING
C3755 S.n3397 VSUBS 0.03fF $ **FLOATING
C3756 S.n3398 VSUBS 0.04fF $ **FLOATING
C3757 S.n3399 VSUBS 0.17fF $ **FLOATING
C3758 S.n3400 VSUBS 0.01fF $ **FLOATING
C3759 S.n3401 VSUBS 0.02fF $ **FLOATING
C3760 S.n3402 VSUBS 0.01fF $ **FLOATING
C3761 S.n3403 VSUBS 0.01fF $ **FLOATING
C3762 S.n3404 VSUBS 0.01fF $ **FLOATING
C3763 S.n3405 VSUBS 0.01fF $ **FLOATING
C3764 S.n3406 VSUBS 0.01fF $ **FLOATING
C3765 S.n3407 VSUBS 0.01fF $ **FLOATING
C3766 S.n3408 VSUBS 0.02fF $ **FLOATING
C3767 S.n3409 VSUBS 0.05fF $ **FLOATING
C3768 S.n3410 VSUBS 0.04fF $ **FLOATING
C3769 S.n3411 VSUBS 0.11fF $ **FLOATING
C3770 S.n3412 VSUBS 0.37fF $ **FLOATING
C3771 S.n3413 VSUBS 0.20fF $ **FLOATING
C3772 S.n3414 VSUBS 4.34fF $ **FLOATING
C3773 S.n3415 VSUBS 0.24fF $ **FLOATING
C3774 S.n3416 VSUBS 1.48fF $ **FLOATING
C3775 S.n3417 VSUBS 1.29fF $ **FLOATING
C3776 S.n3418 VSUBS 0.27fF $ **FLOATING
C3777 S.n3419 VSUBS 1.87fF $ **FLOATING
C3778 S.n3420 VSUBS 0.04fF $ **FLOATING
C3779 S.n3421 VSUBS 0.07fF $ **FLOATING
C3780 S.n3422 VSUBS 0.05fF $ **FLOATING
C3781 S.n3423 VSUBS 0.86fF $ **FLOATING
C3782 S.n3424 VSUBS 0.01fF $ **FLOATING
C3783 S.n3425 VSUBS 0.01fF $ **FLOATING
C3784 S.n3426 VSUBS 0.01fF $ **FLOATING
C3785 S.n3427 VSUBS 0.07fF $ **FLOATING
C3786 S.n3428 VSUBS 0.68fF $ **FLOATING
C3787 S.n3429 VSUBS 0.71fF $ **FLOATING
C3788 S.t832 VSUBS 0.02fF
C3789 S.n3430 VSUBS 0.24fF $ **FLOATING
C3790 S.n3431 VSUBS 0.35fF $ **FLOATING
C3791 S.n3432 VSUBS 0.60fF $ **FLOATING
C3792 S.n3433 VSUBS 0.12fF $ **FLOATING
C3793 S.t378 VSUBS 0.02fF
C3794 S.n3434 VSUBS 0.14fF $ **FLOATING
C3795 S.n3436 VSUBS 0.69fF $ **FLOATING
C3796 S.n3437 VSUBS 0.22fF $ **FLOATING
C3797 S.n3438 VSUBS 0.22fF $ **FLOATING
C3798 S.n3439 VSUBS 0.69fF $ **FLOATING
C3799 S.n3440 VSUBS 1.14fF $ **FLOATING
C3800 S.n3441 VSUBS 0.22fF $ **FLOATING
C3801 S.n3442 VSUBS 0.25fF $ **FLOATING
C3802 S.n3443 VSUBS 0.09fF $ **FLOATING
C3803 S.n3444 VSUBS 2.29fF $ **FLOATING
C3804 S.t867 VSUBS 0.02fF
C3805 S.n3445 VSUBS 0.24fF $ **FLOATING
C3806 S.n3446 VSUBS 0.90fF $ **FLOATING
C3807 S.n3447 VSUBS 0.05fF $ **FLOATING
C3808 S.t761 VSUBS 0.02fF
C3809 S.n3448 VSUBS 0.12fF $ **FLOATING
C3810 S.n3449 VSUBS 0.14fF $ **FLOATING
C3811 S.n3451 VSUBS 1.86fF $ **FLOATING
C3812 S.n3452 VSUBS 0.45fF $ **FLOATING
C3813 S.n3453 VSUBS 0.22fF $ **FLOATING
C3814 S.n3454 VSUBS 0.38fF $ **FLOATING
C3815 S.n3455 VSUBS 0.16fF $ **FLOATING
C3816 S.n3456 VSUBS 0.28fF $ **FLOATING
C3817 S.n3457 VSUBS 0.21fF $ **FLOATING
C3818 S.n3458 VSUBS 0.30fF $ **FLOATING
C3819 S.n3459 VSUBS 0.41fF $ **FLOATING
C3820 S.n3460 VSUBS 0.20fF $ **FLOATING
C3821 S.t645 VSUBS 0.02fF
C3822 S.n3461 VSUBS 0.24fF $ **FLOATING
C3823 S.n3462 VSUBS 0.35fF $ **FLOATING
C3824 S.n3463 VSUBS 0.60fF $ **FLOATING
C3825 S.n3464 VSUBS 0.12fF $ **FLOATING
C3826 S.t205 VSUBS 0.02fF
C3827 S.n3465 VSUBS 0.14fF $ **FLOATING
C3828 S.n3467 VSUBS 0.04fF $ **FLOATING
C3829 S.n3468 VSUBS 0.03fF $ **FLOATING
C3830 S.n3469 VSUBS 0.03fF $ **FLOATING
C3831 S.n3470 VSUBS 0.10fF $ **FLOATING
C3832 S.n3471 VSUBS 0.36fF $ **FLOATING
C3833 S.n3472 VSUBS 0.37fF $ **FLOATING
C3834 S.n3473 VSUBS 0.10fF $ **FLOATING
C3835 S.n3474 VSUBS 0.12fF $ **FLOATING
C3836 S.n3475 VSUBS 0.07fF $ **FLOATING
C3837 S.n3476 VSUBS 0.12fF $ **FLOATING
C3838 S.n3477 VSUBS 0.18fF $ **FLOATING
C3839 S.n3478 VSUBS 3.95fF $ **FLOATING
C3840 S.t682 VSUBS 0.02fF
C3841 S.n3479 VSUBS 0.24fF $ **FLOATING
C3842 S.n3480 VSUBS 0.90fF $ **FLOATING
C3843 S.n3481 VSUBS 0.05fF $ **FLOATING
C3844 S.t589 VSUBS 0.02fF
C3845 S.n3482 VSUBS 0.12fF $ **FLOATING
C3846 S.n3483 VSUBS 0.14fF $ **FLOATING
C3847 S.n3485 VSUBS 0.25fF $ **FLOATING
C3848 S.n3486 VSUBS 0.09fF $ **FLOATING
C3849 S.n3487 VSUBS 0.21fF $ **FLOATING
C3850 S.n3488 VSUBS 1.27fF $ **FLOATING
C3851 S.n3489 VSUBS 0.52fF $ **FLOATING
C3852 S.n3490 VSUBS 1.86fF $ **FLOATING
C3853 S.n3491 VSUBS 0.12fF $ **FLOATING
C3854 S.t551 VSUBS 0.02fF
C3855 S.n3492 VSUBS 0.14fF $ **FLOATING
C3856 S.t992 VSUBS 0.02fF
C3857 S.n3494 VSUBS 0.24fF $ **FLOATING
C3858 S.n3495 VSUBS 0.35fF $ **FLOATING
C3859 S.n3496 VSUBS 0.60fF $ **FLOATING
C3860 S.n3497 VSUBS 1.56fF $ **FLOATING
C3861 S.n3498 VSUBS 2.42fF $ **FLOATING
C3862 S.t1023 VSUBS 0.02fF
C3863 S.n3499 VSUBS 0.24fF $ **FLOATING
C3864 S.n3500 VSUBS 0.90fF $ **FLOATING
C3865 S.n3501 VSUBS 0.05fF $ **FLOATING
C3866 S.t931 VSUBS 0.02fF
C3867 S.n3502 VSUBS 0.12fF $ **FLOATING
C3868 S.n3503 VSUBS 0.14fF $ **FLOATING
C3869 S.n3505 VSUBS 1.87fF $ **FLOATING
C3870 S.n3506 VSUBS 0.06fF $ **FLOATING
C3871 S.n3507 VSUBS 0.03fF $ **FLOATING
C3872 S.n3508 VSUBS 0.03fF $ **FLOATING
C3873 S.n3509 VSUBS 0.98fF $ **FLOATING
C3874 S.n3510 VSUBS 0.02fF $ **FLOATING
C3875 S.n3511 VSUBS 0.01fF $ **FLOATING
C3876 S.n3512 VSUBS 0.02fF $ **FLOATING
C3877 S.n3513 VSUBS 0.08fF $ **FLOATING
C3878 S.n3514 VSUBS 0.36fF $ **FLOATING
C3879 S.n3515 VSUBS 1.83fF $ **FLOATING
C3880 S.t235 VSUBS 0.02fF
C3881 S.n3516 VSUBS 0.24fF $ **FLOATING
C3882 S.n3517 VSUBS 0.35fF $ **FLOATING
C3883 S.n3518 VSUBS 0.60fF $ **FLOATING
C3884 S.n3519 VSUBS 0.12fF $ **FLOATING
C3885 S.t897 VSUBS 0.02fF
C3886 S.n3520 VSUBS 0.14fF $ **FLOATING
C3887 S.n3522 VSUBS 0.69fF $ **FLOATING
C3888 S.n3523 VSUBS 0.22fF $ **FLOATING
C3889 S.n3524 VSUBS 0.22fF $ **FLOATING
C3890 S.n3525 VSUBS 0.69fF $ **FLOATING
C3891 S.n3526 VSUBS 1.14fF $ **FLOATING
C3892 S.n3527 VSUBS 0.22fF $ **FLOATING
C3893 S.n3528 VSUBS 0.25fF $ **FLOATING
C3894 S.n3529 VSUBS 0.09fF $ **FLOATING
C3895 S.n3530 VSUBS 1.86fF $ **FLOATING
C3896 S.t262 VSUBS 0.02fF
C3897 S.n3531 VSUBS 0.24fF $ **FLOATING
C3898 S.n3532 VSUBS 0.90fF $ **FLOATING
C3899 S.n3533 VSUBS 0.05fF $ **FLOATING
C3900 S.t172 VSUBS 0.02fF
C3901 S.n3534 VSUBS 0.12fF $ **FLOATING
C3902 S.n3535 VSUBS 0.14fF $ **FLOATING
C3903 S.n3537 VSUBS 14.09fF $ **FLOATING
C3904 S.n3538 VSUBS 0.06fF $ **FLOATING
C3905 S.n3539 VSUBS 0.20fF $ **FLOATING
C3906 S.n3540 VSUBS 0.09fF $ **FLOATING
C3907 S.n3541 VSUBS 0.20fF $ **FLOATING
C3908 S.n3542 VSUBS 0.09fF $ **FLOATING
C3909 S.n3543 VSUBS 0.30fF $ **FLOATING
C3910 S.n3544 VSUBS 0.69fF $ **FLOATING
C3911 S.n3545 VSUBS 0.44fF $ **FLOATING
C3912 S.n3546 VSUBS 2.30fF $ **FLOATING
C3913 S.n3547 VSUBS 0.12fF $ **FLOATING
C3914 S.t1075 VSUBS 0.02fF
C3915 S.n3548 VSUBS 0.14fF $ **FLOATING
C3916 S.t433 VSUBS 0.02fF
C3917 S.n3550 VSUBS 0.24fF $ **FLOATING
C3918 S.n3551 VSUBS 0.35fF $ **FLOATING
C3919 S.n3552 VSUBS 0.60fF $ **FLOATING
C3920 S.n3553 VSUBS 1.88fF $ **FLOATING
C3921 S.n3554 VSUBS 0.17fF $ **FLOATING
C3922 S.n3555 VSUBS 0.76fF $ **FLOATING
C3923 S.n3556 VSUBS 0.25fF $ **FLOATING
C3924 S.n3557 VSUBS 0.29fF $ **FLOATING
C3925 S.n3558 VSUBS 0.31fF $ **FLOATING
C3926 S.n3559 VSUBS 0.46fF $ **FLOATING
C3927 S.n3560 VSUBS 0.16fF $ **FLOATING
C3928 S.n3561 VSUBS 1.90fF $ **FLOATING
C3929 S.t355 VSUBS 0.02fF
C3930 S.n3562 VSUBS 0.12fF $ **FLOATING
C3931 S.n3563 VSUBS 0.14fF $ **FLOATING
C3932 S.t470 VSUBS 0.02fF
C3933 S.n3565 VSUBS 0.24fF $ **FLOATING
C3934 S.n3566 VSUBS 0.90fF $ **FLOATING
C3935 S.n3567 VSUBS 0.05fF $ **FLOATING
C3936 S.n3568 VSUBS 1.86fF $ **FLOATING
C3937 S.n3569 VSUBS 0.12fF $ **FLOATING
C3938 S.t491 VSUBS 0.02fF
C3939 S.n3570 VSUBS 0.14fF $ **FLOATING
C3940 S.t671 VSUBS 0.02fF
C3941 S.n3572 VSUBS 1.20fF $ **FLOATING
C3942 S.n3573 VSUBS 0.36fF $ **FLOATING
C3943 S.n3574 VSUBS 1.21fF $ **FLOATING
C3944 S.n3575 VSUBS 0.60fF $ **FLOATING
C3945 S.n3576 VSUBS 0.35fF $ **FLOATING
C3946 S.n3577 VSUBS 0.62fF $ **FLOATING
C3947 S.n3578 VSUBS 1.14fF $ **FLOATING
C3948 S.n3579 VSUBS 2.15fF $ **FLOATING
C3949 S.n3580 VSUBS 0.59fF $ **FLOATING
C3950 S.n3581 VSUBS 0.01fF $ **FLOATING
C3951 S.n3582 VSUBS 0.96fF $ **FLOATING
C3952 S.t27 VSUBS 14.53fF
C3953 S.n3583 VSUBS 14.40fF $ **FLOATING
C3954 S.n3585 VSUBS 0.37fF $ **FLOATING
C3955 S.n3586 VSUBS 0.23fF $ **FLOATING
C3956 S.n3587 VSUBS 2.76fF $ **FLOATING
C3957 S.n3588 VSUBS 2.43fF $ **FLOATING
C3958 S.n3589 VSUBS 3.96fF $ **FLOATING
C3959 S.n3590 VSUBS 0.25fF $ **FLOATING
C3960 S.n3591 VSUBS 0.01fF $ **FLOATING
C3961 S.t314 VSUBS 0.02fF
C3962 S.n3592 VSUBS 0.25fF $ **FLOATING
C3963 S.t811 VSUBS 0.02fF
C3964 S.n3593 VSUBS 0.94fF $ **FLOATING
C3965 S.n3594 VSUBS 0.70fF $ **FLOATING
C3966 S.n3595 VSUBS 1.87fF $ **FLOATING
C3967 S.n3596 VSUBS 1.71fF $ **FLOATING
C3968 S.t1017 VSUBS 0.02fF
C3969 S.n3597 VSUBS 0.24fF $ **FLOATING
C3970 S.n3598 VSUBS 0.35fF $ **FLOATING
C3971 S.n3599 VSUBS 0.60fF $ **FLOATING
C3972 S.n3600 VSUBS 0.12fF $ **FLOATING
C3973 S.t721 VSUBS 0.02fF
C3974 S.n3601 VSUBS 0.14fF $ **FLOATING
C3975 S.n3603 VSUBS 1.14fF $ **FLOATING
C3976 S.n3604 VSUBS 0.22fF $ **FLOATING
C3977 S.n3605 VSUBS 0.25fF $ **FLOATING
C3978 S.n3606 VSUBS 0.09fF $ **FLOATING
C3979 S.n3607 VSUBS 2.41fF $ **FLOATING
C3980 S.t19 VSUBS 0.02fF
C3981 S.n3608 VSUBS 0.24fF $ **FLOATING
C3982 S.n3609 VSUBS 0.90fF $ **FLOATING
C3983 S.n3610 VSUBS 0.05fF $ **FLOATING
C3984 S.t1038 VSUBS 0.02fF
C3985 S.n3611 VSUBS 0.12fF $ **FLOATING
C3986 S.n3612 VSUBS 0.14fF $ **FLOATING
C3987 S.n3614 VSUBS 1.86fF $ **FLOATING
C3988 S.n3615 VSUBS 0.47fF $ **FLOATING
C3989 S.n3616 VSUBS 0.09fF $ **FLOATING
C3990 S.n3617 VSUBS 0.32fF $ **FLOATING
C3991 S.n3618 VSUBS 0.30fF $ **FLOATING
C3992 S.n3619 VSUBS 0.76fF $ **FLOATING
C3993 S.n3620 VSUBS 0.58fF $ **FLOATING
C3994 S.t911 VSUBS 0.02fF
C3995 S.n3621 VSUBS 0.24fF $ **FLOATING
C3996 S.n3622 VSUBS 0.35fF $ **FLOATING
C3997 S.n3623 VSUBS 0.60fF $ **FLOATING
C3998 S.n3624 VSUBS 0.12fF $ **FLOATING
C3999 S.t554 VSUBS 0.02fF
C4000 S.n3625 VSUBS 0.14fF $ **FLOATING
C4001 S.n3627 VSUBS 2.58fF $ **FLOATING
C4002 S.n3628 VSUBS 2.13fF $ **FLOATING
C4003 S.t1028 VSUBS 0.02fF
C4004 S.n3629 VSUBS 0.24fF $ **FLOATING
C4005 S.n3630 VSUBS 0.90fF $ **FLOATING
C4006 S.n3631 VSUBS 0.05fF $ **FLOATING
C4007 S.t338 VSUBS 0.02fF
C4008 S.n3632 VSUBS 0.12fF $ **FLOATING
C4009 S.n3633 VSUBS 0.14fF $ **FLOATING
C4010 S.n3635 VSUBS 0.77fF $ **FLOATING
C4011 S.n3636 VSUBS 2.27fF $ **FLOATING
C4012 S.n3637 VSUBS 1.86fF $ **FLOATING
C4013 S.n3638 VSUBS 0.12fF $ **FLOATING
C4014 S.t902 VSUBS 0.02fF
C4015 S.n3639 VSUBS 0.14fF $ **FLOATING
C4016 S.t148 VSUBS 0.02fF
C4017 S.n3641 VSUBS 0.24fF $ **FLOATING
C4018 S.n3642 VSUBS 0.35fF $ **FLOATING
C4019 S.n3643 VSUBS 0.60fF $ **FLOATING
C4020 S.n3644 VSUBS 1.37fF $ **FLOATING
C4021 S.n3645 VSUBS 0.70fF $ **FLOATING
C4022 S.n3646 VSUBS 1.13fF $ **FLOATING
C4023 S.n3647 VSUBS 0.35fF $ **FLOATING
C4024 S.n3648 VSUBS 2.00fF $ **FLOATING
C4025 S.t265 VSUBS 0.02fF
C4026 S.n3649 VSUBS 0.24fF $ **FLOATING
C4027 S.n3650 VSUBS 0.90fF $ **FLOATING
C4028 S.n3651 VSUBS 0.05fF $ **FLOATING
C4029 S.t174 VSUBS 0.02fF
C4030 S.n3652 VSUBS 0.12fF $ **FLOATING
C4031 S.n3653 VSUBS 0.14fF $ **FLOATING
C4032 S.n3655 VSUBS 1.87fF $ **FLOATING
C4033 S.n3656 VSUBS 1.86fF $ **FLOATING
C4034 S.t507 VSUBS 0.02fF
C4035 S.n3657 VSUBS 0.24fF $ **FLOATING
C4036 S.n3658 VSUBS 0.35fF $ **FLOATING
C4037 S.n3659 VSUBS 0.60fF $ **FLOATING
C4038 S.n3660 VSUBS 0.12fF $ **FLOATING
C4039 S.t134 VSUBS 0.02fF
C4040 S.n3661 VSUBS 0.14fF $ **FLOATING
C4041 S.n3663 VSUBS 1.14fF $ **FLOATING
C4042 S.n3664 VSUBS 0.22fF $ **FLOATING
C4043 S.n3665 VSUBS 0.25fF $ **FLOATING
C4044 S.n3666 VSUBS 0.09fF $ **FLOATING
C4045 S.n3667 VSUBS 1.86fF $ **FLOATING
C4046 S.t612 VSUBS 0.02fF
C4047 S.n3668 VSUBS 0.24fF $ **FLOATING
C4048 S.n3669 VSUBS 0.90fF $ **FLOATING
C4049 S.n3670 VSUBS 0.05fF $ **FLOATING
C4050 S.t523 VSUBS 0.02fF
C4051 S.n3671 VSUBS 0.12fF $ **FLOATING
C4052 S.n3672 VSUBS 0.14fF $ **FLOATING
C4053 S.n3674 VSUBS 14.09fF $ **FLOATING
C4054 S.n3675 VSUBS 1.86fF $ **FLOATING
C4055 S.n3676 VSUBS 2.64fF $ **FLOATING
C4056 S.t439 VSUBS 0.02fF
C4057 S.n3677 VSUBS 0.24fF $ **FLOATING
C4058 S.n3678 VSUBS 0.35fF $ **FLOATING
C4059 S.n3679 VSUBS 0.60fF $ **FLOATING
C4060 S.n3680 VSUBS 0.12fF $ **FLOATING
C4061 S.t525 VSUBS 0.02fF
C4062 S.n3681 VSUBS 0.14fF $ **FLOATING
C4063 S.n3683 VSUBS 2.77fF $ **FLOATING
C4064 S.n3684 VSUBS 2.27fF $ **FLOATING
C4065 S.t900 VSUBS 0.02fF
C4066 S.n3685 VSUBS 0.12fF $ **FLOATING
C4067 S.n3686 VSUBS 0.14fF $ **FLOATING
C4068 S.t804 VSUBS 0.02fF
C4069 S.n3688 VSUBS 0.24fF $ **FLOATING
C4070 S.n3689 VSUBS 0.90fF $ **FLOATING
C4071 S.n3690 VSUBS 0.05fF $ **FLOATING
C4072 S.n3691 VSUBS 1.86fF $ **FLOATING
C4073 S.n3692 VSUBS 2.64fF $ **FLOATING
C4074 S.t778 VSUBS 0.02fF
C4075 S.n3693 VSUBS 0.24fF $ **FLOATING
C4076 S.n3694 VSUBS 0.35fF $ **FLOATING
C4077 S.n3695 VSUBS 0.60fF $ **FLOATING
C4078 S.n3696 VSUBS 0.12fF $ **FLOATING
C4079 S.t868 VSUBS 0.02fF
C4080 S.n3697 VSUBS 0.14fF $ **FLOATING
C4081 S.n3699 VSUBS 2.77fF $ **FLOATING
C4082 S.n3700 VSUBS 2.27fF $ **FLOATING
C4083 S.t133 VSUBS 0.02fF
C4084 S.n3701 VSUBS 0.12fF $ **FLOATING
C4085 S.n3702 VSUBS 0.14fF $ **FLOATING
C4086 S.t11 VSUBS 0.02fF
C4087 S.n3704 VSUBS 0.24fF $ **FLOATING
C4088 S.n3705 VSUBS 0.90fF $ **FLOATING
C4089 S.n3706 VSUBS 0.05fF $ **FLOATING
C4090 S.n3707 VSUBS 1.86fF $ **FLOATING
C4091 S.n3708 VSUBS 2.64fF $ **FLOATING
C4092 S.t1122 VSUBS 0.02fF
C4093 S.n3709 VSUBS 0.24fF $ **FLOATING
C4094 S.n3710 VSUBS 0.35fF $ **FLOATING
C4095 S.n3711 VSUBS 0.60fF $ **FLOATING
C4096 S.n3712 VSUBS 0.12fF $ **FLOATING
C4097 S.t93 VSUBS 0.02fF
C4098 S.n3713 VSUBS 0.14fF $ **FLOATING
C4099 S.n3715 VSUBS 2.77fF $ **FLOATING
C4100 S.n3716 VSUBS 2.27fF $ **FLOATING
C4101 S.t489 VSUBS 0.02fF
C4102 S.n3717 VSUBS 0.12fF $ **FLOATING
C4103 S.n3718 VSUBS 0.14fF $ **FLOATING
C4104 S.t387 VSUBS 0.02fF
C4105 S.n3720 VSUBS 0.24fF $ **FLOATING
C4106 S.n3721 VSUBS 0.90fF $ **FLOATING
C4107 S.n3722 VSUBS 0.05fF $ **FLOATING
C4108 S.n3723 VSUBS 1.86fF $ **FLOATING
C4109 S.n3724 VSUBS 2.65fF $ **FLOATING
C4110 S.t356 VSUBS 0.02fF
C4111 S.n3725 VSUBS 0.24fF $ **FLOATING
C4112 S.n3726 VSUBS 0.35fF $ **FLOATING
C4113 S.n3727 VSUBS 0.60fF $ **FLOATING
C4114 S.n3728 VSUBS 0.12fF $ **FLOATING
C4115 S.t456 VSUBS 0.02fF
C4116 S.n3729 VSUBS 0.14fF $ **FLOATING
C4117 S.n3731 VSUBS 5.11fF $ **FLOATING
C4118 S.t833 VSUBS 0.02fF
C4119 S.n3732 VSUBS 0.12fF $ **FLOATING
C4120 S.n3733 VSUBS 0.14fF $ **FLOATING
C4121 S.t726 VSUBS 0.02fF
C4122 S.n3735 VSUBS 0.24fF $ **FLOATING
C4123 S.n3736 VSUBS 0.90fF $ **FLOATING
C4124 S.n3737 VSUBS 0.05fF $ **FLOATING
C4125 S.n3738 VSUBS 2.70fF $ **FLOATING
C4126 S.n3739 VSUBS 1.58fF $ **FLOATING
C4127 S.n3740 VSUBS 0.12fF $ **FLOATING
C4128 S.t493 VSUBS 0.02fF
C4129 S.n3741 VSUBS 0.14fF $ **FLOATING
C4130 S.t490 VSUBS 0.02fF
C4131 S.n3743 VSUBS 0.24fF $ **FLOATING
C4132 S.n3744 VSUBS 0.35fF $ **FLOATING
C4133 S.n3745 VSUBS 0.60fF $ **FLOATING
C4134 S.n3746 VSUBS 0.07fF $ **FLOATING
C4135 S.n3747 VSUBS 0.01fF $ **FLOATING
C4136 S.n3748 VSUBS 0.23fF $ **FLOATING
C4137 S.n3749 VSUBS 1.15fF $ **FLOATING
C4138 S.n3750 VSUBS 1.33fF $ **FLOATING
C4139 S.n3751 VSUBS 2.27fF $ **FLOATING
C4140 S.t54 VSUBS 0.02fF
C4141 S.n3752 VSUBS 0.12fF $ **FLOATING
C4142 S.n3753 VSUBS 0.14fF $ **FLOATING
C4143 S.t1096 VSUBS 0.02fF
C4144 S.n3755 VSUBS 0.24fF $ **FLOATING
C4145 S.n3756 VSUBS 0.90fF $ **FLOATING
C4146 S.n3757 VSUBS 0.05fF $ **FLOATING
C4147 S.t53 VSUBS 32.33fF
C4148 S.t869 VSUBS 0.02fF
C4149 S.n3758 VSUBS 0.12fF $ **FLOATING
C4150 S.n3759 VSUBS 0.14fF $ **FLOATING
C4151 S.t959 VSUBS 0.02fF
C4152 S.n3761 VSUBS 0.24fF $ **FLOATING
C4153 S.n3762 VSUBS 0.90fF $ **FLOATING
C4154 S.n3763 VSUBS 0.05fF $ **FLOATING
C4155 S.t846 VSUBS 0.02fF
C4156 S.n3764 VSUBS 0.24fF $ **FLOATING
C4157 S.n3765 VSUBS 0.35fF $ **FLOATING
C4158 S.n3766 VSUBS 0.60fF $ **FLOATING
C4159 S.n3767 VSUBS 0.31fF $ **FLOATING
C4160 S.n3768 VSUBS 1.08fF $ **FLOATING
C4161 S.n3769 VSUBS 0.15fF $ **FLOATING
C4162 S.n3770 VSUBS 2.08fF $ **FLOATING
C4163 S.n3771 VSUBS 2.91fF $ **FLOATING
C4164 S.n3772 VSUBS 1.86fF $ **FLOATING
C4165 S.n3773 VSUBS 0.12fF $ **FLOATING
C4166 S.t130 VSUBS 0.02fF
C4167 S.n3774 VSUBS 0.14fF $ **FLOATING
C4168 S.t581 VSUBS 0.02fF
C4169 S.n3776 VSUBS 0.24fF $ **FLOATING
C4170 S.n3777 VSUBS 0.35fF $ **FLOATING
C4171 S.n3778 VSUBS 0.60fF $ **FLOATING
C4172 S.n3779 VSUBS 0.91fF $ **FLOATING
C4173 S.n3780 VSUBS 0.31fF $ **FLOATING
C4174 S.n3781 VSUBS 0.91fF $ **FLOATING
C4175 S.n3782 VSUBS 1.08fF $ **FLOATING
C4176 S.n3783 VSUBS 0.15fF $ **FLOATING
C4177 S.n3784 VSUBS 4.90fF $ **FLOATING
C4178 S.t521 VSUBS 0.02fF
C4179 S.n3785 VSUBS 0.12fF $ **FLOATING
C4180 S.n3786 VSUBS 0.14fF $ **FLOATING
C4181 S.t611 VSUBS 0.02fF
C4182 S.n3788 VSUBS 0.24fF $ **FLOATING
C4183 S.n3789 VSUBS 0.90fF $ **FLOATING
C4184 S.n3790 VSUBS 0.05fF $ **FLOATING
C4185 S.n3791 VSUBS 1.86fF $ **FLOATING
C4186 S.n3792 VSUBS 2.64fF $ **FLOATING
C4187 S.t64 VSUBS 0.02fF
C4188 S.n3793 VSUBS 0.24fF $ **FLOATING
C4189 S.n3794 VSUBS 0.35fF $ **FLOATING
C4190 S.n3795 VSUBS 0.60fF $ **FLOATING
C4191 S.n3796 VSUBS 0.12fF $ **FLOATING
C4192 S.t1100 VSUBS 0.02fF
C4193 S.n3797 VSUBS 0.14fF $ **FLOATING
C4194 S.n3799 VSUBS 1.86fF $ **FLOATING
C4195 S.n3800 VSUBS 2.64fF $ **FLOATING
C4196 S.t71 VSUBS 0.02fF
C4197 S.n3801 VSUBS 0.24fF $ **FLOATING
C4198 S.n3802 VSUBS 0.35fF $ **FLOATING
C4199 S.n3803 VSUBS 0.60fF $ **FLOATING
C4200 S.t199 VSUBS 0.02fF
C4201 S.n3804 VSUBS 0.24fF $ **FLOATING
C4202 S.n3805 VSUBS 0.90fF $ **FLOATING
C4203 S.n3806 VSUBS 0.05fF $ **FLOATING
C4204 S.t94 VSUBS 0.02fF
C4205 S.n3807 VSUBS 0.12fF $ **FLOATING
C4206 S.n3808 VSUBS 0.14fF $ **FLOATING
C4207 S.n3810 VSUBS 0.12fF $ **FLOATING
C4208 S.t882 VSUBS 0.02fF
C4209 S.n3811 VSUBS 0.14fF $ **FLOATING
C4210 S.n3813 VSUBS 2.27fF $ **FLOATING
C4211 S.n3814 VSUBS 2.91fF $ **FLOATING
C4212 S.n3815 VSUBS 5.10fF $ **FLOATING
C4213 S.t915 VSUBS 0.02fF
C4214 S.n3816 VSUBS 0.12fF $ **FLOATING
C4215 S.n3817 VSUBS 0.14fF $ **FLOATING
C4216 S.t267 VSUBS 0.02fF
C4217 S.n3819 VSUBS 0.24fF $ **FLOATING
C4218 S.n3820 VSUBS 0.90fF $ **FLOATING
C4219 S.n3821 VSUBS 0.05fF $ **FLOATING
C4220 S.n3822 VSUBS 1.86fF $ **FLOATING
C4221 S.n3823 VSUBS 2.64fF $ **FLOATING
C4222 S.t428 VSUBS 0.02fF
C4223 S.n3824 VSUBS 0.24fF $ **FLOATING
C4224 S.n3825 VSUBS 0.35fF $ **FLOATING
C4225 S.n3826 VSUBS 0.60fF $ **FLOATING
C4226 S.n3827 VSUBS 0.12fF $ **FLOATING
C4227 S.t330 VSUBS 0.02fF
C4228 S.n3828 VSUBS 0.14fF $ **FLOATING
C4229 S.n3830 VSUBS 5.11fF $ **FLOATING
C4230 S.t717 VSUBS 0.02fF
C4231 S.n3831 VSUBS 0.12fF $ **FLOATING
C4232 S.n3832 VSUBS 0.14fF $ **FLOATING
C4233 S.t614 VSUBS 0.02fF
C4234 S.n3834 VSUBS 0.24fF $ **FLOATING
C4235 S.n3835 VSUBS 0.90fF $ **FLOATING
C4236 S.n3836 VSUBS 0.05fF $ **FLOATING
C4237 S.n3837 VSUBS 1.86fF $ **FLOATING
C4238 S.n3838 VSUBS 2.64fF $ **FLOATING
C4239 S.t767 VSUBS 0.02fF
C4240 S.n3839 VSUBS 0.24fF $ **FLOATING
C4241 S.n3840 VSUBS 0.35fF $ **FLOATING
C4242 S.n3841 VSUBS 0.60fF $ **FLOATING
C4243 S.n3842 VSUBS 0.12fF $ **FLOATING
C4244 S.t674 VSUBS 0.02fF
C4245 S.n3843 VSUBS 0.14fF $ **FLOATING
C4246 S.n3845 VSUBS 5.11fF $ **FLOATING
C4247 S.t1053 VSUBS 0.02fF
C4248 S.n3846 VSUBS 0.12fF $ **FLOATING
C4249 S.n3847 VSUBS 0.14fF $ **FLOATING
C4250 S.t965 VSUBS 0.02fF
C4251 S.n3849 VSUBS 0.24fF $ **FLOATING
C4252 S.n3850 VSUBS 0.90fF $ **FLOATING
C4253 S.n3851 VSUBS 0.05fF $ **FLOATING
C4254 S.n3852 VSUBS 1.86fF $ **FLOATING
C4255 S.n3853 VSUBS 2.64fF $ **FLOATING
C4256 S.t1108 VSUBS 0.02fF
C4257 S.n3854 VSUBS 0.24fF $ **FLOATING
C4258 S.n3855 VSUBS 0.35fF $ **FLOATING
C4259 S.n3856 VSUBS 0.60fF $ **FLOATING
C4260 S.n3857 VSUBS 0.12fF $ **FLOATING
C4261 S.t1020 VSUBS 0.02fF
C4262 S.n3858 VSUBS 0.14fF $ **FLOATING
C4263 S.n3860 VSUBS 4.84fF $ **FLOATING
C4264 S.t293 VSUBS 0.02fF
C4265 S.n3861 VSUBS 0.12fF $ **FLOATING
C4266 S.n3862 VSUBS 0.14fF $ **FLOATING
C4267 S.t202 VSUBS 0.02fF
C4268 S.n3864 VSUBS 0.24fF $ **FLOATING
C4269 S.n3865 VSUBS 0.90fF $ **FLOATING
C4270 S.n3866 VSUBS 0.05fF $ **FLOATING
C4271 S.n3867 VSUBS 1.86fF $ **FLOATING
C4272 S.n3868 VSUBS 2.64fF $ **FLOATING
C4273 S.t343 VSUBS 0.02fF
C4274 S.n3869 VSUBS 0.24fF $ **FLOATING
C4275 S.n3870 VSUBS 0.35fF $ **FLOATING
C4276 S.n3871 VSUBS 0.60fF $ **FLOATING
C4277 S.n3872 VSUBS 0.12fF $ **FLOATING
C4278 S.t255 VSUBS 0.02fF
C4279 S.n3873 VSUBS 0.14fF $ **FLOATING
C4280 S.n3875 VSUBS 5.38fF $ **FLOATING
C4281 S.t637 VSUBS 0.02fF
C4282 S.n3876 VSUBS 0.12fF $ **FLOATING
C4283 S.n3877 VSUBS 0.14fF $ **FLOATING
C4284 S.t549 VSUBS 0.02fF
C4285 S.n3879 VSUBS 0.24fF $ **FLOATING
C4286 S.n3880 VSUBS 0.90fF $ **FLOATING
C4287 S.n3881 VSUBS 0.05fF $ **FLOATING
C4288 S.t129 VSUBS 31.95fF
C4289 S.t276 VSUBS 0.02fF
C4290 S.n3882 VSUBS 0.01fF $ **FLOATING
C4291 S.n3883 VSUBS 0.25fF $ **FLOATING
C4292 S.t331 VSUBS 0.02fF
C4293 S.n3885 VSUBS 1.18fF $ **FLOATING
C4294 S.n3886 VSUBS 0.05fF $ **FLOATING
C4295 S.t299 VSUBS 0.02fF
C4296 S.n3887 VSUBS 0.63fF $ **FLOATING
C4297 S.n3888 VSUBS 0.60fF $ **FLOATING
C4298 S.n3889 VSUBS 8.88fF $ **FLOATING
C4299 S.n3890 VSUBS 8.88fF $ **FLOATING
C4300 S.n3891 VSUBS 0.59fF $ **FLOATING
C4301 S.n3892 VSUBS 0.21fF $ **FLOATING
C4302 S.n3893 VSUBS 0.59fF $ **FLOATING
C4303 S.n3894 VSUBS 2.55fF $ **FLOATING
C4304 S.n3895 VSUBS 0.28fF $ **FLOATING
C4305 S.t10 VSUBS 14.53fF
C4306 S.n3896 VSUBS 15.80fF $ **FLOATING
C4307 S.n3897 VSUBS 0.76fF $ **FLOATING
C4308 S.n3898 VSUBS 0.27fF $ **FLOATING
C4309 S.n3899 VSUBS 3.96fF $ **FLOATING
C4310 S.n3900 VSUBS 1.34fF $ **FLOATING
C4311 S.n3901 VSUBS 0.01fF $ **FLOATING
C4312 S.n3902 VSUBS 0.02fF $ **FLOATING
C4313 S.n3903 VSUBS 0.03fF $ **FLOATING
C4314 S.n3904 VSUBS 0.04fF $ **FLOATING
C4315 S.n3905 VSUBS 0.17fF $ **FLOATING
C4316 S.n3906 VSUBS 0.01fF $ **FLOATING
C4317 S.n3907 VSUBS 0.02fF $ **FLOATING
C4318 S.n3908 VSUBS 0.01fF $ **FLOATING
C4319 S.n3909 VSUBS 0.01fF $ **FLOATING
C4320 S.n3910 VSUBS 0.01fF $ **FLOATING
C4321 S.n3911 VSUBS 0.01fF $ **FLOATING
C4322 S.n3912 VSUBS 0.01fF $ **FLOATING
C4323 S.n3913 VSUBS 0.01fF $ **FLOATING
C4324 S.n3914 VSUBS 0.02fF $ **FLOATING
C4325 S.n3915 VSUBS 0.05fF $ **FLOATING
C4326 S.n3916 VSUBS 0.04fF $ **FLOATING
C4327 S.n3917 VSUBS 0.11fF $ **FLOATING
C4328 S.n3918 VSUBS 0.37fF $ **FLOATING
C4329 S.n3919 VSUBS 0.20fF $ **FLOATING
C4330 S.n3920 VSUBS 4.34fF $ **FLOATING
C4331 S.n3921 VSUBS 0.24fF $ **FLOATING
C4332 S.n3922 VSUBS 1.48fF $ **FLOATING
C4333 S.n3923 VSUBS 1.29fF $ **FLOATING
C4334 S.n3924 VSUBS 0.27fF $ **FLOATING
C4335 S.n3925 VSUBS 1.86fF $ **FLOATING
C4336 S.n3926 VSUBS 0.45fF $ **FLOATING
C4337 S.n3927 VSUBS 0.22fF $ **FLOATING
C4338 S.n3928 VSUBS 0.38fF $ **FLOATING
C4339 S.n3929 VSUBS 0.16fF $ **FLOATING
C4340 S.n3930 VSUBS 0.28fF $ **FLOATING
C4341 S.n3931 VSUBS 0.21fF $ **FLOATING
C4342 S.n3932 VSUBS 0.30fF $ **FLOATING
C4343 S.n3933 VSUBS 0.41fF $ **FLOATING
C4344 S.n3934 VSUBS 0.20fF $ **FLOATING
C4345 S.t573 VSUBS 0.02fF
C4346 S.n3935 VSUBS 0.24fF $ **FLOATING
C4347 S.n3936 VSUBS 0.35fF $ **FLOATING
C4348 S.n3937 VSUBS 0.60fF $ **FLOATING
C4349 S.n3938 VSUBS 0.12fF $ **FLOATING
C4350 S.t214 VSUBS 0.02fF
C4351 S.n3939 VSUBS 0.14fF $ **FLOATING
C4352 S.n3941 VSUBS 0.04fF $ **FLOATING
C4353 S.n3942 VSUBS 0.03fF $ **FLOATING
C4354 S.n3943 VSUBS 0.03fF $ **FLOATING
C4355 S.n3944 VSUBS 0.10fF $ **FLOATING
C4356 S.n3945 VSUBS 0.36fF $ **FLOATING
C4357 S.n3946 VSUBS 0.37fF $ **FLOATING
C4358 S.n3947 VSUBS 0.10fF $ **FLOATING
C4359 S.n3948 VSUBS 0.12fF $ **FLOATING
C4360 S.n3949 VSUBS 0.07fF $ **FLOATING
C4361 S.n3950 VSUBS 0.12fF $ **FLOATING
C4362 S.n3951 VSUBS 0.18fF $ **FLOATING
C4363 S.n3952 VSUBS 3.95fF $ **FLOATING
C4364 S.t690 VSUBS 0.02fF
C4365 S.n3953 VSUBS 0.24fF $ **FLOATING
C4366 S.n3954 VSUBS 0.90fF $ **FLOATING
C4367 S.n3955 VSUBS 0.05fF $ **FLOATING
C4368 S.t594 VSUBS 0.02fF
C4369 S.n3956 VSUBS 0.12fF $ **FLOATING
C4370 S.n3957 VSUBS 0.14fF $ **FLOATING
C4371 S.n3959 VSUBS 0.25fF $ **FLOATING
C4372 S.n3960 VSUBS 0.09fF $ **FLOATING
C4373 S.n3961 VSUBS 0.21fF $ **FLOATING
C4374 S.n3962 VSUBS 1.27fF $ **FLOATING
C4375 S.n3963 VSUBS 0.52fF $ **FLOATING
C4376 S.n3964 VSUBS 1.86fF $ **FLOATING
C4377 S.n3965 VSUBS 0.12fF $ **FLOATING
C4378 S.t24 VSUBS 0.02fF
C4379 S.n3966 VSUBS 0.14fF $ **FLOATING
C4380 S.t413 VSUBS 0.02fF
C4381 S.n3968 VSUBS 0.24fF $ **FLOATING
C4382 S.n3969 VSUBS 0.35fF $ **FLOATING
C4383 S.n3970 VSUBS 0.60fF $ **FLOATING
C4384 S.n3971 VSUBS 1.56fF $ **FLOATING
C4385 S.n3972 VSUBS 2.42fF $ **FLOATING
C4386 S.t536 VSUBS 0.02fF
C4387 S.n3973 VSUBS 0.24fF $ **FLOATING
C4388 S.n3974 VSUBS 0.90fF $ **FLOATING
C4389 S.n3975 VSUBS 0.05fF $ **FLOATING
C4390 S.t435 VSUBS 0.02fF
C4391 S.n3976 VSUBS 0.12fF $ **FLOATING
C4392 S.n3977 VSUBS 0.14fF $ **FLOATING
C4393 S.n3979 VSUBS 1.87fF $ **FLOATING
C4394 S.n3980 VSUBS 0.06fF $ **FLOATING
C4395 S.n3981 VSUBS 0.03fF $ **FLOATING
C4396 S.n3982 VSUBS 0.03fF $ **FLOATING
C4397 S.n3983 VSUBS 0.98fF $ **FLOATING
C4398 S.n3984 VSUBS 0.02fF $ **FLOATING
C4399 S.n3985 VSUBS 0.01fF $ **FLOATING
C4400 S.n3986 VSUBS 0.02fF $ **FLOATING
C4401 S.n3987 VSUBS 0.08fF $ **FLOATING
C4402 S.n3988 VSUBS 0.36fF $ **FLOATING
C4403 S.n3989 VSUBS 1.83fF $ **FLOATING
C4404 S.t755 VSUBS 0.02fF
C4405 S.n3990 VSUBS 0.24fF $ **FLOATING
C4406 S.n3991 VSUBS 0.35fF $ **FLOATING
C4407 S.n3992 VSUBS 0.60fF $ **FLOATING
C4408 S.n3993 VSUBS 0.12fF $ **FLOATING
C4409 S.t398 VSUBS 0.02fF
C4410 S.n3994 VSUBS 0.14fF $ **FLOATING
C4411 S.n3996 VSUBS 0.69fF $ **FLOATING
C4412 S.n3997 VSUBS 0.22fF $ **FLOATING
C4413 S.n3998 VSUBS 0.22fF $ **FLOATING
C4414 S.n3999 VSUBS 0.69fF $ **FLOATING
C4415 S.n4000 VSUBS 1.14fF $ **FLOATING
C4416 S.n4001 VSUBS 0.22fF $ **FLOATING
C4417 S.n4002 VSUBS 0.25fF $ **FLOATING
C4418 S.n4003 VSUBS 0.09fF $ **FLOATING
C4419 S.n4004 VSUBS 1.86fF $ **FLOATING
C4420 S.t879 VSUBS 0.02fF
C4421 S.n4005 VSUBS 0.24fF $ **FLOATING
C4422 S.n4006 VSUBS 0.90fF $ **FLOATING
C4423 S.n4007 VSUBS 0.05fF $ **FLOATING
C4424 S.t777 VSUBS 0.02fF
C4425 S.n4008 VSUBS 0.12fF $ **FLOATING
C4426 S.n4009 VSUBS 0.14fF $ **FLOATING
C4427 S.n4011 VSUBS 14.09fF $ **FLOATING
C4428 S.n4012 VSUBS 1.70fF $ **FLOATING
C4429 S.n4013 VSUBS 0.65fF $ **FLOATING
C4430 S.n4014 VSUBS 0.68fF $ **FLOATING
C4431 S.n4015 VSUBS 0.71fF $ **FLOATING
C4432 S.n4016 VSUBS 0.36fF $ **FLOATING
C4433 S.t177 VSUBS 0.02fF
C4434 S.n4017 VSUBS 0.24fF $ **FLOATING
C4435 S.n4018 VSUBS 0.35fF $ **FLOATING
C4436 S.n4019 VSUBS 0.60fF $ **FLOATING
C4437 S.n4020 VSUBS 0.12fF $ **FLOATING
C4438 S.t923 VSUBS 0.02fF
C4439 S.n4021 VSUBS 0.14fF $ **FLOATING
C4440 S.n4023 VSUBS 0.31fF $ **FLOATING
C4441 S.n4024 VSUBS 0.22fF $ **FLOATING
C4442 S.n4025 VSUBS 0.65fF $ **FLOATING
C4443 S.n4026 VSUBS 0.94fF $ **FLOATING
C4444 S.n4027 VSUBS 0.22fF $ **FLOATING
C4445 S.n4028 VSUBS 0.20fF $ **FLOATING
C4446 S.n4029 VSUBS 0.20fF $ **FLOATING
C4447 S.n4030 VSUBS 0.06fF $ **FLOATING
C4448 S.n4031 VSUBS 0.09fF $ **FLOATING
C4449 S.n4032 VSUBS 0.09fF $ **FLOATING
C4450 S.n4033 VSUBS 1.65fF $ **FLOATING
C4451 S.t197 VSUBS 0.02fF
C4452 S.n4034 VSUBS 0.12fF $ **FLOATING
C4453 S.n4035 VSUBS 0.14fF $ **FLOATING
C4454 S.t290 VSUBS 0.02fF
C4455 S.n4037 VSUBS 0.24fF $ **FLOATING
C4456 S.n4038 VSUBS 0.90fF $ **FLOATING
C4457 S.n4039 VSUBS 0.05fF $ **FLOATING
C4458 S.n4040 VSUBS 1.86fF $ **FLOATING
C4459 S.n4041 VSUBS 0.12fF $ **FLOATING
C4460 S.t984 VSUBS 0.02fF
C4461 S.n4042 VSUBS 0.14fF $ **FLOATING
C4462 S.t253 VSUBS 0.02fF
C4463 S.n4044 VSUBS 0.12fF $ **FLOATING
C4464 S.n4045 VSUBS 0.14fF $ **FLOATING
C4465 S.t375 VSUBS 0.02fF
C4466 S.n4047 VSUBS 0.24fF $ **FLOATING
C4467 S.n4048 VSUBS 0.90fF $ **FLOATING
C4468 S.n4049 VSUBS 0.05fF $ **FLOATING
C4469 S.t239 VSUBS 0.02fF
C4470 S.n4050 VSUBS 0.24fF $ **FLOATING
C4471 S.n4051 VSUBS 0.35fF $ **FLOATING
C4472 S.n4052 VSUBS 0.60fF $ **FLOATING
C4473 S.n4053 VSUBS 0.31fF $ **FLOATING
C4474 S.n4054 VSUBS 1.08fF $ **FLOATING
C4475 S.n4055 VSUBS 0.15fF $ **FLOATING
C4476 S.n4056 VSUBS 2.08fF $ **FLOATING
C4477 S.n4057 VSUBS 2.91fF $ **FLOATING
C4478 S.n4058 VSUBS 1.86fF $ **FLOATING
C4479 S.n4059 VSUBS 0.12fF $ **FLOATING
C4480 S.t738 VSUBS 0.02fF
C4481 S.n4060 VSUBS 0.14fF $ **FLOATING
C4482 S.t1092 VSUBS 0.02fF
C4483 S.n4062 VSUBS 0.24fF $ **FLOATING
C4484 S.n4063 VSUBS 0.35fF $ **FLOATING
C4485 S.n4064 VSUBS 0.60fF $ **FLOATING
C4486 S.n4065 VSUBS 0.91fF $ **FLOATING
C4487 S.n4066 VSUBS 0.31fF $ **FLOATING
C4488 S.n4067 VSUBS 0.91fF $ **FLOATING
C4489 S.n4068 VSUBS 1.08fF $ **FLOATING
C4490 S.n4069 VSUBS 0.15fF $ **FLOATING
C4491 S.n4070 VSUBS 4.90fF $ **FLOATING
C4492 S.t1121 VSUBS 0.02fF
C4493 S.n4071 VSUBS 0.12fF $ **FLOATING
C4494 S.n4072 VSUBS 0.14fF $ **FLOATING
C4495 S.t110 VSUBS 0.02fF
C4496 S.n4074 VSUBS 0.24fF $ **FLOATING
C4497 S.n4075 VSUBS 0.90fF $ **FLOATING
C4498 S.n4076 VSUBS 0.05fF $ **FLOATING
C4499 S.n4077 VSUBS 1.86fF $ **FLOATING
C4500 S.n4078 VSUBS 2.64fF $ **FLOATING
C4501 S.t325 VSUBS 0.02fF
C4502 S.n4079 VSUBS 0.24fF $ **FLOATING
C4503 S.n4080 VSUBS 0.35fF $ **FLOATING
C4504 S.n4081 VSUBS 0.60fF $ **FLOATING
C4505 S.n4082 VSUBS 0.12fF $ **FLOATING
C4506 S.t1073 VSUBS 0.02fF
C4507 S.n4083 VSUBS 0.14fF $ **FLOATING
C4508 S.n4085 VSUBS 1.86fF $ **FLOATING
C4509 S.n4086 VSUBS 2.64fF $ **FLOATING
C4510 S.t588 VSUBS 0.02fF
C4511 S.n4087 VSUBS 0.24fF $ **FLOATING
C4512 S.n4088 VSUBS 0.35fF $ **FLOATING
C4513 S.n4089 VSUBS 0.60fF $ **FLOATING
C4514 S.t707 VSUBS 0.02fF
C4515 S.n4090 VSUBS 0.24fF $ **FLOATING
C4516 S.n4091 VSUBS 0.90fF $ **FLOATING
C4517 S.n4092 VSUBS 0.05fF $ **FLOATING
C4518 S.t604 VSUBS 0.02fF
C4519 S.n4093 VSUBS 0.12fF $ **FLOATING
C4520 S.n4094 VSUBS 0.14fF $ **FLOATING
C4521 S.n4096 VSUBS 0.12fF $ **FLOATING
C4522 S.t223 VSUBS 0.02fF
C4523 S.n4097 VSUBS 0.14fF $ **FLOATING
C4524 S.n4099 VSUBS 2.27fF $ **FLOATING
C4525 S.n4100 VSUBS 2.91fF $ **FLOATING
C4526 S.n4101 VSUBS 5.10fF $ **FLOATING
C4527 S.t353 VSUBS 0.02fF
C4528 S.n4102 VSUBS 0.12fF $ **FLOATING
C4529 S.n4103 VSUBS 0.14fF $ **FLOATING
C4530 S.t468 VSUBS 0.02fF
C4531 S.n4105 VSUBS 0.24fF $ **FLOATING
C4532 S.n4106 VSUBS 0.90fF $ **FLOATING
C4533 S.n4107 VSUBS 0.05fF $ **FLOATING
C4534 S.n4108 VSUBS 1.86fF $ **FLOATING
C4535 S.n4109 VSUBS 2.64fF $ **FLOATING
C4536 S.t450 VSUBS 0.02fF
C4537 S.n4110 VSUBS 0.24fF $ **FLOATING
C4538 S.n4111 VSUBS 0.35fF $ **FLOATING
C4539 S.n4112 VSUBS 0.60fF $ **FLOATING
C4540 S.n4113 VSUBS 0.12fF $ **FLOATING
C4541 S.t535 VSUBS 0.02fF
C4542 S.n4114 VSUBS 0.14fF $ **FLOATING
C4543 S.n4116 VSUBS 5.11fF $ **FLOATING
C4544 S.t759 VSUBS 0.02fF
C4545 S.n4117 VSUBS 0.12fF $ **FLOATING
C4546 S.n4118 VSUBS 0.14fF $ **FLOATING
C4547 S.t816 VSUBS 0.02fF
C4548 S.n4120 VSUBS 0.24fF $ **FLOATING
C4549 S.n4121 VSUBS 0.90fF $ **FLOATING
C4550 S.n4122 VSUBS 0.05fF $ **FLOATING
C4551 S.n4123 VSUBS 1.86fF $ **FLOATING
C4552 S.n4124 VSUBS 2.64fF $ **FLOATING
C4553 S.t793 VSUBS 0.02fF
C4554 S.n4125 VSUBS 0.24fF $ **FLOATING
C4555 S.n4126 VSUBS 0.35fF $ **FLOATING
C4556 S.n4127 VSUBS 0.60fF $ **FLOATING
C4557 S.n4128 VSUBS 0.12fF $ **FLOATING
C4558 S.t878 VSUBS 0.02fF
C4559 S.n4129 VSUBS 0.14fF $ **FLOATING
C4560 S.n4131 VSUBS 5.11fF $ **FLOATING
C4561 S.t147 VSUBS 0.02fF
C4562 S.n4132 VSUBS 0.12fF $ **FLOATING
C4563 S.n4133 VSUBS 0.14fF $ **FLOATING
C4564 S.t28 VSUBS 0.02fF
C4565 S.n4135 VSUBS 0.24fF $ **FLOATING
C4566 S.n4136 VSUBS 0.90fF $ **FLOATING
C4567 S.n4137 VSUBS 0.05fF $ **FLOATING
C4568 S.n4138 VSUBS 1.86fF $ **FLOATING
C4569 S.n4139 VSUBS 2.64fF $ **FLOATING
C4570 S.t1133 VSUBS 0.02fF
C4571 S.n4140 VSUBS 0.24fF $ **FLOATING
C4572 S.n4141 VSUBS 0.35fF $ **FLOATING
C4573 S.n4142 VSUBS 0.60fF $ **FLOATING
C4574 S.n4143 VSUBS 0.12fF $ **FLOATING
C4575 S.t109 VSUBS 0.02fF
C4576 S.n4144 VSUBS 0.14fF $ **FLOATING
C4577 S.n4146 VSUBS 5.11fF $ **FLOATING
C4578 S.t505 VSUBS 0.02fF
C4579 S.n4147 VSUBS 0.12fF $ **FLOATING
C4580 S.n4148 VSUBS 0.14fF $ **FLOATING
C4581 S.t399 VSUBS 0.02fF
C4582 S.n4150 VSUBS 0.24fF $ **FLOATING
C4583 S.n4151 VSUBS 0.90fF $ **FLOATING
C4584 S.n4152 VSUBS 0.05fF $ **FLOATING
C4585 S.n4153 VSUBS 1.86fF $ **FLOATING
C4586 S.n4154 VSUBS 2.64fF $ **FLOATING
C4587 S.t373 VSUBS 0.02fF
C4588 S.n4155 VSUBS 0.24fF $ **FLOATING
C4589 S.n4156 VSUBS 0.35fF $ **FLOATING
C4590 S.n4157 VSUBS 0.60fF $ **FLOATING
C4591 S.n4158 VSUBS 0.12fF $ **FLOATING
C4592 S.t467 VSUBS 0.02fF
C4593 S.n4159 VSUBS 0.14fF $ **FLOATING
C4594 S.n4161 VSUBS 4.84fF $ **FLOATING
C4595 S.t845 VSUBS 0.02fF
C4596 S.n4162 VSUBS 0.12fF $ **FLOATING
C4597 S.n4163 VSUBS 0.14fF $ **FLOATING
C4598 S.t740 VSUBS 0.02fF
C4599 S.n4165 VSUBS 0.24fF $ **FLOATING
C4600 S.n4166 VSUBS 0.90fF $ **FLOATING
C4601 S.n4167 VSUBS 0.05fF $ **FLOATING
C4602 S.n4168 VSUBS 1.86fF $ **FLOATING
C4603 S.n4169 VSUBS 2.64fF $ **FLOATING
C4604 S.t711 VSUBS 0.02fF
C4605 S.n4170 VSUBS 0.24fF $ **FLOATING
C4606 S.n4171 VSUBS 0.35fF $ **FLOATING
C4607 S.n4172 VSUBS 0.60fF $ **FLOATING
C4608 S.n4173 VSUBS 0.12fF $ **FLOATING
C4609 S.t805 VSUBS 0.02fF
C4610 S.n4174 VSUBS 0.14fF $ **FLOATING
C4611 S.n4176 VSUBS 1.86fF $ **FLOATING
C4612 S.n4177 VSUBS 2.65fF $ **FLOATING
C4613 S.t723 VSUBS 0.02fF
C4614 S.n4178 VSUBS 0.24fF $ **FLOATING
C4615 S.n4179 VSUBS 0.35fF $ **FLOATING
C4616 S.n4180 VSUBS 0.60fF $ **FLOATING
C4617 S.t441 VSUBS 0.02fF
C4618 S.n4181 VSUBS 1.20fF $ **FLOATING
C4619 S.n4182 VSUBS 0.60fF $ **FLOATING
C4620 S.n4183 VSUBS 1.14fF $ **FLOATING
C4621 S.n4184 VSUBS 2.15fF $ **FLOATING
C4622 S.n4185 VSUBS 0.01fF $ **FLOATING
C4623 S.n4186 VSUBS 0.96fF $ **FLOATING
C4624 S.t4 VSUBS 14.53fF
C4625 S.n4187 VSUBS 14.40fF $ **FLOATING
C4626 S.n4189 VSUBS 0.37fF $ **FLOATING
C4627 S.n4190 VSUBS 0.23fF $ **FLOATING
C4628 S.n4191 VSUBS 2.85fF $ **FLOATING
C4629 S.n4192 VSUBS 2.43fF $ **FLOATING
C4630 S.n4193 VSUBS 2.50fF $ **FLOATING
C4631 S.n4194 VSUBS 3.90fF $ **FLOATING
C4632 S.n4195 VSUBS 0.25fF $ **FLOATING
C4633 S.n4196 VSUBS 0.01fF $ **FLOATING
C4634 S.t67 VSUBS 0.02fF
C4635 S.n4197 VSUBS 0.25fF $ **FLOATING
C4636 S.t558 VSUBS 0.02fF
C4637 S.n4198 VSUBS 0.94fF $ **FLOATING
C4638 S.n4199 VSUBS 0.70fF $ **FLOATING
C4639 S.n4200 VSUBS 1.86fF $ **FLOATING
C4640 S.n4201 VSUBS 0.47fF $ **FLOATING
C4641 S.n4202 VSUBS 0.09fF $ **FLOATING
C4642 S.n4203 VSUBS 0.32fF $ **FLOATING
C4643 S.n4204 VSUBS 0.30fF $ **FLOATING
C4644 S.n4205 VSUBS 0.76fF $ **FLOATING
C4645 S.n4206 VSUBS 0.58fF $ **FLOATING
C4646 S.t780 VSUBS 0.02fF
C4647 S.n4207 VSUBS 0.24fF $ **FLOATING
C4648 S.n4208 VSUBS 0.35fF $ **FLOATING
C4649 S.n4209 VSUBS 0.60fF $ **FLOATING
C4650 S.n4210 VSUBS 0.12fF $ **FLOATING
C4651 S.t481 VSUBS 0.02fF
C4652 S.n4211 VSUBS 0.14fF $ **FLOATING
C4653 S.n4213 VSUBS 1.42fF $ **FLOATING
C4654 S.n4214 VSUBS 2.13fF $ **FLOATING
C4655 S.t905 VSUBS 0.02fF
C4656 S.n4215 VSUBS 0.24fF $ **FLOATING
C4657 S.n4216 VSUBS 0.90fF $ **FLOATING
C4658 S.n4217 VSUBS 0.05fF $ **FLOATING
C4659 S.t801 VSUBS 0.02fF
C4660 S.n4218 VSUBS 0.12fF $ **FLOATING
C4661 S.n4219 VSUBS 0.14fF $ **FLOATING
C4662 S.n4221 VSUBS 0.77fF $ **FLOATING
C4663 S.n4222 VSUBS 2.27fF $ **FLOATING
C4664 S.n4223 VSUBS 1.86fF $ **FLOATING
C4665 S.n4224 VSUBS 0.12fF $ **FLOATING
C4666 S.t291 VSUBS 0.02fF
C4667 S.n4225 VSUBS 0.14fF $ **FLOATING
C4668 S.t650 VSUBS 0.02fF
C4669 S.n4227 VSUBS 0.24fF $ **FLOATING
C4670 S.n4228 VSUBS 0.35fF $ **FLOATING
C4671 S.n4229 VSUBS 0.60fF $ **FLOATING
C4672 S.n4230 VSUBS 1.37fF $ **FLOATING
C4673 S.n4231 VSUBS 0.70fF $ **FLOATING
C4674 S.n4232 VSUBS 1.13fF $ **FLOATING
C4675 S.n4233 VSUBS 0.35fF $ **FLOATING
C4676 S.n4234 VSUBS 2.00fF $ **FLOATING
C4677 S.t790 VSUBS 0.02fF
C4678 S.n4235 VSUBS 0.24fF $ **FLOATING
C4679 S.n4236 VSUBS 0.90fF $ **FLOATING
C4680 S.n4237 VSUBS 0.05fF $ **FLOATING
C4681 S.t84 VSUBS 0.02fF
C4682 S.n4238 VSUBS 0.12fF $ **FLOATING
C4683 S.n4239 VSUBS 0.14fF $ **FLOATING
C4684 S.n4241 VSUBS 1.87fF $ **FLOATING
C4685 S.n4242 VSUBS 1.86fF $ **FLOATING
C4686 S.t996 VSUBS 0.02fF
C4687 S.n4243 VSUBS 0.24fF $ **FLOATING
C4688 S.n4244 VSUBS 0.35fF $ **FLOATING
C4689 S.n4245 VSUBS 0.60fF $ **FLOATING
C4690 S.n4246 VSUBS 0.12fF $ **FLOATING
C4691 S.t636 VSUBS 0.02fF
C4692 S.n4247 VSUBS 0.14fF $ **FLOATING
C4693 S.n4249 VSUBS 1.14fF $ **FLOATING
C4694 S.n4250 VSUBS 0.22fF $ **FLOATING
C4695 S.n4251 VSUBS 0.25fF $ **FLOATING
C4696 S.n4252 VSUBS 0.09fF $ **FLOATING
C4697 S.n4253 VSUBS 1.86fF $ **FLOATING
C4698 S.t1135 VSUBS 0.02fF
C4699 S.n4254 VSUBS 0.24fF $ **FLOATING
C4700 S.n4255 VSUBS 0.90fF $ **FLOATING
C4701 S.n4256 VSUBS 0.05fF $ **FLOATING
C4702 S.t1019 VSUBS 0.02fF
C4703 S.n4257 VSUBS 0.12fF $ **FLOATING
C4704 S.n4258 VSUBS 0.14fF $ **FLOATING
C4705 S.n4260 VSUBS 14.09fF $ **FLOATING
C4706 S.n4261 VSUBS 1.86fF $ **FLOATING
C4707 S.n4262 VSUBS 2.64fF $ **FLOATING
C4708 S.t933 VSUBS 0.02fF
C4709 S.n4263 VSUBS 0.24fF $ **FLOATING
C4710 S.n4264 VSUBS 0.35fF $ **FLOATING
C4711 S.n4265 VSUBS 0.60fF $ **FLOATING
C4712 S.n4266 VSUBS 0.12fF $ **FLOATING
C4713 S.t620 VSUBS 0.02fF
C4714 S.n4267 VSUBS 0.14fF $ **FLOATING
C4715 S.n4269 VSUBS 2.77fF $ **FLOATING
C4716 S.n4270 VSUBS 2.27fF $ **FLOATING
C4717 S.t949 VSUBS 0.02fF
C4718 S.n4271 VSUBS 0.12fF $ **FLOATING
C4719 S.n4272 VSUBS 0.14fF $ **FLOATING
C4720 S.t1049 VSUBS 0.02fF
C4721 S.n4274 VSUBS 0.24fF $ **FLOATING
C4722 S.n4275 VSUBS 0.90fF $ **FLOATING
C4723 S.n4276 VSUBS 0.05fF $ **FLOATING
C4724 S.n4277 VSUBS 1.86fF $ **FLOATING
C4725 S.n4278 VSUBS 2.64fF $ **FLOATING
C4726 S.t798 VSUBS 0.02fF
C4727 S.n4279 VSUBS 0.24fF $ **FLOATING
C4728 S.n4280 VSUBS 0.35fF $ **FLOATING
C4729 S.n4281 VSUBS 0.60fF $ **FLOATING
C4730 S.n4282 VSUBS 0.12fF $ **FLOATING
C4731 S.t889 VSUBS 0.02fF
C4732 S.n4283 VSUBS 0.14fF $ **FLOATING
C4733 S.n4285 VSUBS 2.77fF $ **FLOATING
C4734 S.n4286 VSUBS 2.27fF $ **FLOATING
C4735 S.t161 VSUBS 0.02fF
C4736 S.n4287 VSUBS 0.12fF $ **FLOATING
C4737 S.n4288 VSUBS 0.14fF $ **FLOATING
C4738 S.t46 VSUBS 0.02fF
C4739 S.n4290 VSUBS 0.24fF $ **FLOATING
C4740 S.n4291 VSUBS 0.90fF $ **FLOATING
C4741 S.n4292 VSUBS 0.05fF $ **FLOATING
C4742 S.n4293 VSUBS 1.86fF $ **FLOATING
C4743 S.n4294 VSUBS 2.64fF $ **FLOATING
C4744 S.t5 VSUBS 0.02fF
C4745 S.n4295 VSUBS 0.24fF $ **FLOATING
C4746 S.n4296 VSUBS 0.35fF $ **FLOATING
C4747 S.n4297 VSUBS 0.60fF $ **FLOATING
C4748 S.n4298 VSUBS 0.12fF $ **FLOATING
C4749 S.t118 VSUBS 0.02fF
C4750 S.n4299 VSUBS 0.14fF $ **FLOATING
C4751 S.n4301 VSUBS 2.77fF $ **FLOATING
C4752 S.n4302 VSUBS 2.27fF $ **FLOATING
C4753 S.t513 VSUBS 0.02fF
C4754 S.n4303 VSUBS 0.12fF $ **FLOATING
C4755 S.n4304 VSUBS 0.14fF $ **FLOATING
C4756 S.t415 VSUBS 0.02fF
C4757 S.n4306 VSUBS 0.24fF $ **FLOATING
C4758 S.n4307 VSUBS 0.90fF $ **FLOATING
C4759 S.n4308 VSUBS 0.05fF $ **FLOATING
C4760 S.n4309 VSUBS 1.86fF $ **FLOATING
C4761 S.n4310 VSUBS 2.64fF $ **FLOATING
C4762 S.t382 VSUBS 0.02fF
C4763 S.n4311 VSUBS 0.24fF $ **FLOATING
C4764 S.n4312 VSUBS 0.35fF $ **FLOATING
C4765 S.n4313 VSUBS 0.60fF $ **FLOATING
C4766 S.n4314 VSUBS 0.12fF $ **FLOATING
C4767 S.t479 VSUBS 0.02fF
C4768 S.n4315 VSUBS 0.14fF $ **FLOATING
C4769 S.n4317 VSUBS 2.77fF $ **FLOATING
C4770 S.n4318 VSUBS 2.27fF $ **FLOATING
C4771 S.t856 VSUBS 0.02fF
C4772 S.n4319 VSUBS 0.12fF $ **FLOATING
C4773 S.n4320 VSUBS 0.14fF $ **FLOATING
C4774 S.t753 VSUBS 0.02fF
C4775 S.n4322 VSUBS 0.24fF $ **FLOATING
C4776 S.n4323 VSUBS 0.90fF $ **FLOATING
C4777 S.n4324 VSUBS 0.05fF $ **FLOATING
C4778 S.n4325 VSUBS 2.70fF $ **FLOATING
C4779 S.n4326 VSUBS 1.58fF $ **FLOATING
C4780 S.n4327 VSUBS 0.12fF $ **FLOATING
C4781 S.t396 VSUBS 0.02fF
C4782 S.n4328 VSUBS 0.14fF $ **FLOATING
C4783 S.t357 VSUBS 0.02fF
C4784 S.n4330 VSUBS 0.24fF $ **FLOATING
C4785 S.n4331 VSUBS 0.35fF $ **FLOATING
C4786 S.n4332 VSUBS 0.60fF $ **FLOATING
C4787 S.n4333 VSUBS 0.07fF $ **FLOATING
C4788 S.n4334 VSUBS 0.01fF $ **FLOATING
C4789 S.n4335 VSUBS 0.23fF $ **FLOATING
C4790 S.n4336 VSUBS 1.15fF $ **FLOATING
C4791 S.n4337 VSUBS 1.33fF $ **FLOATING
C4792 S.n4338 VSUBS 2.27fF $ **FLOATING
C4793 S.t443 VSUBS 0.02fF
C4794 S.n4339 VSUBS 0.12fF $ **FLOATING
C4795 S.n4340 VSUBS 0.14fF $ **FLOATING
C4796 S.t971 VSUBS 0.02fF
C4797 S.n4342 VSUBS 0.24fF $ **FLOATING
C4798 S.n4343 VSUBS 0.90fF $ **FLOATING
C4799 S.n4344 VSUBS 0.05fF $ **FLOATING
C4800 S.t66 VSUBS 32.33fF
C4801 S.t1094 VSUBS 0.02fF
C4802 S.n4345 VSUBS 0.24fF $ **FLOATING
C4803 S.n4346 VSUBS 0.90fF $ **FLOATING
C4804 S.n4347 VSUBS 0.05fF $ **FLOATING
C4805 S.t82 VSUBS 0.02fF
C4806 S.n4348 VSUBS 0.12fF $ **FLOATING
C4807 S.n4349 VSUBS 0.14fF $ **FLOATING
C4808 S.n4351 VSUBS 0.12fF $ **FLOATING
C4809 S.t820 VSUBS 0.02fF
C4810 S.n4352 VSUBS 0.14fF $ **FLOATING
C4811 S.n4354 VSUBS 5.11fF $ **FLOATING
C4812 S.n4355 VSUBS 5.38fF $ **FLOATING
C4813 S.t69 VSUBS 0.02fF
C4814 S.n4356 VSUBS 0.12fF $ **FLOATING
C4815 S.n4357 VSUBS 0.14fF $ **FLOATING
C4816 S.t1077 VSUBS 0.02fF
C4817 S.n4359 VSUBS 0.24fF $ **FLOATING
C4818 S.n4360 VSUBS 0.90fF $ **FLOATING
C4819 S.n4361 VSUBS 0.05fF $ **FLOATING
C4820 S.t23 VSUBS 31.95fF
C4821 S.t982 VSUBS 0.02fF
C4822 S.n4362 VSUBS 0.01fF $ **FLOATING
C4823 S.n4363 VSUBS 0.25fF $ **FLOATING
C4824 S.t183 VSUBS 0.02fF
C4825 S.n4365 VSUBS 1.18fF $ **FLOATING
C4826 S.n4366 VSUBS 0.05fF $ **FLOATING
C4827 S.t38 VSUBS 0.02fF
C4828 S.n4367 VSUBS 0.63fF $ **FLOATING
C4829 S.n4368 VSUBS 0.60fF $ **FLOATING
C4830 S.n4369 VSUBS 0.59fF $ **FLOATING
C4831 S.n4370 VSUBS 0.21fF $ **FLOATING
C4832 S.n4371 VSUBS 0.59fF $ **FLOATING
C4833 S.n4372 VSUBS 2.55fF $ **FLOATING
C4834 S.n4373 VSUBS 0.28fF $ **FLOATING
C4835 S.t37 VSUBS 14.53fF
C4836 S.n4374 VSUBS 15.80fF $ **FLOATING
C4837 S.n4375 VSUBS 0.76fF $ **FLOATING
C4838 S.n4376 VSUBS 0.27fF $ **FLOATING
C4839 S.n4377 VSUBS 3.96fF $ **FLOATING
C4840 S.n4378 VSUBS 1.34fF $ **FLOATING
C4841 S.n4379 VSUBS 0.01fF $ **FLOATING
C4842 S.n4380 VSUBS 0.02fF $ **FLOATING
C4843 S.n4381 VSUBS 0.03fF $ **FLOATING
C4844 S.n4382 VSUBS 0.04fF $ **FLOATING
C4845 S.n4383 VSUBS 0.17fF $ **FLOATING
C4846 S.n4384 VSUBS 0.01fF $ **FLOATING
C4847 S.n4385 VSUBS 0.02fF $ **FLOATING
C4848 S.n4386 VSUBS 0.01fF $ **FLOATING
C4849 S.n4387 VSUBS 0.01fF $ **FLOATING
C4850 S.n4388 VSUBS 0.01fF $ **FLOATING
C4851 S.n4389 VSUBS 0.01fF $ **FLOATING
C4852 S.n4390 VSUBS 0.01fF $ **FLOATING
C4853 S.n4391 VSUBS 0.01fF $ **FLOATING
C4854 S.n4392 VSUBS 0.02fF $ **FLOATING
C4855 S.n4393 VSUBS 0.05fF $ **FLOATING
C4856 S.n4394 VSUBS 0.04fF $ **FLOATING
C4857 S.n4395 VSUBS 0.11fF $ **FLOATING
C4858 S.n4396 VSUBS 0.37fF $ **FLOATING
C4859 S.n4397 VSUBS 0.20fF $ **FLOATING
C4860 S.n4398 VSUBS 4.34fF $ **FLOATING
C4861 S.n4399 VSUBS 0.24fF $ **FLOATING
C4862 S.n4400 VSUBS 1.48fF $ **FLOATING
C4863 S.n4401 VSUBS 1.24fF $ **FLOATING
C4864 S.n4402 VSUBS 0.27fF $ **FLOATING
C4865 S.n4403 VSUBS 0.25fF $ **FLOATING
C4866 S.n4404 VSUBS 0.09fF $ **FLOATING
C4867 S.n4405 VSUBS 0.21fF $ **FLOATING
C4868 S.n4406 VSUBS 1.27fF $ **FLOATING
C4869 S.n4407 VSUBS 0.52fF $ **FLOATING
C4870 S.n4408 VSUBS 1.86fF $ **FLOATING
C4871 S.n4409 VSUBS 0.12fF $ **FLOATING
C4872 S.t1064 VSUBS 0.02fF
C4873 S.n4410 VSUBS 0.14fF $ **FLOATING
C4874 S.t313 VSUBS 0.02fF
C4875 S.n4412 VSUBS 0.24fF $ **FLOATING
C4876 S.n4413 VSUBS 0.35fF $ **FLOATING
C4877 S.n4414 VSUBS 0.60fF $ **FLOATING
C4878 S.n4415 VSUBS 1.56fF $ **FLOATING
C4879 S.n4416 VSUBS 2.42fF $ **FLOATING
C4880 S.t458 VSUBS 0.02fF
C4881 S.n4417 VSUBS 0.24fF $ **FLOATING
C4882 S.n4418 VSUBS 0.90fF $ **FLOATING
C4883 S.n4419 VSUBS 0.05fF $ **FLOATING
C4884 S.t344 VSUBS 0.02fF
C4885 S.n4420 VSUBS 0.12fF $ **FLOATING
C4886 S.n4421 VSUBS 0.14fF $ **FLOATING
C4887 S.n4423 VSUBS 1.87fF $ **FLOATING
C4888 S.n4424 VSUBS 0.06fF $ **FLOATING
C4889 S.n4425 VSUBS 0.03fF $ **FLOATING
C4890 S.n4426 VSUBS 0.03fF $ **FLOATING
C4891 S.n4427 VSUBS 0.98fF $ **FLOATING
C4892 S.n4428 VSUBS 0.02fF $ **FLOATING
C4893 S.n4429 VSUBS 0.01fF $ **FLOATING
C4894 S.n4430 VSUBS 0.02fF $ **FLOATING
C4895 S.n4431 VSUBS 0.08fF $ **FLOATING
C4896 S.n4432 VSUBS 0.36fF $ **FLOATING
C4897 S.n4433 VSUBS 1.83fF $ **FLOATING
C4898 S.t153 VSUBS 0.02fF
C4899 S.n4434 VSUBS 0.24fF $ **FLOATING
C4900 S.n4435 VSUBS 0.35fF $ **FLOATING
C4901 S.n4436 VSUBS 0.60fF $ **FLOATING
C4902 S.n4437 VSUBS 0.12fF $ **FLOATING
C4903 S.t908 VSUBS 0.02fF
C4904 S.n4438 VSUBS 0.14fF $ **FLOATING
C4905 S.n4440 VSUBS 0.69fF $ **FLOATING
C4906 S.n4441 VSUBS 0.22fF $ **FLOATING
C4907 S.n4442 VSUBS 0.22fF $ **FLOATING
C4908 S.n4443 VSUBS 0.69fF $ **FLOATING
C4909 S.n4444 VSUBS 1.14fF $ **FLOATING
C4910 S.n4445 VSUBS 0.22fF $ **FLOATING
C4911 S.n4446 VSUBS 0.25fF $ **FLOATING
C4912 S.n4447 VSUBS 0.09fF $ **FLOATING
C4913 S.n4448 VSUBS 1.86fF $ **FLOATING
C4914 S.t269 VSUBS 0.02fF
C4915 S.n4449 VSUBS 0.24fF $ **FLOATING
C4916 S.n4450 VSUBS 0.90fF $ **FLOATING
C4917 S.n4451 VSUBS 0.05fF $ **FLOATING
C4918 S.t179 VSUBS 0.02fF
C4919 S.n4452 VSUBS 0.12fF $ **FLOATING
C4920 S.n4453 VSUBS 0.14fF $ **FLOATING
C4921 S.n4455 VSUBS 14.09fF $ **FLOATING
C4922 S.n4456 VSUBS 2.36fF $ **FLOATING
C4923 S.n4457 VSUBS 0.45fF $ **FLOATING
C4924 S.n4458 VSUBS 0.22fF $ **FLOATING
C4925 S.n4459 VSUBS 0.38fF $ **FLOATING
C4926 S.n4460 VSUBS 0.16fF $ **FLOATING
C4927 S.n4461 VSUBS 0.28fF $ **FLOATING
C4928 S.n4462 VSUBS 0.21fF $ **FLOATING
C4929 S.n4463 VSUBS 0.30fF $ **FLOATING
C4930 S.n4464 VSUBS 0.20fF $ **FLOATING
C4931 S.t1021 VSUBS 0.02fF
C4932 S.n4465 VSUBS 0.24fF $ **FLOATING
C4933 S.n4466 VSUBS 0.35fF $ **FLOATING
C4934 S.n4467 VSUBS 0.60fF $ **FLOATING
C4935 S.n4468 VSUBS 0.12fF $ **FLOATING
C4936 S.t661 VSUBS 0.02fF
C4937 S.n4469 VSUBS 0.14fF $ **FLOATING
C4938 S.n4471 VSUBS 0.19fF $ **FLOATING
C4939 S.n4472 VSUBS 1.56fF $ **FLOATING
C4940 S.n4473 VSUBS 2.18fF $ **FLOATING
C4941 S.n4474 VSUBS 0.32fF $ **FLOATING
C4942 S.n4475 VSUBS 2.36fF $ **FLOATING
C4943 S.t1043 VSUBS 0.02fF
C4944 S.n4476 VSUBS 0.12fF $ **FLOATING
C4945 S.n4477 VSUBS 0.14fF $ **FLOATING
C4946 S.t29 VSUBS 0.02fF
C4947 S.n4479 VSUBS 0.24fF $ **FLOATING
C4948 S.n4480 VSUBS 0.90fF $ **FLOATING
C4949 S.n4481 VSUBS 0.05fF $ **FLOATING
C4950 S.n4482 VSUBS 1.86fF $ **FLOATING
C4951 S.n4483 VSUBS 0.12fF $ **FLOATING
C4952 S.t404 VSUBS 0.02fF
C4953 S.n4484 VSUBS 0.14fF $ **FLOATING
C4954 S.t783 VSUBS 0.02fF
C4955 S.n4486 VSUBS 0.12fF $ **FLOATING
C4956 S.n4487 VSUBS 0.14fF $ **FLOATING
C4957 S.t881 VSUBS 0.02fF
C4958 S.n4489 VSUBS 0.24fF $ **FLOATING
C4959 S.n4490 VSUBS 0.90fF $ **FLOATING
C4960 S.n4491 VSUBS 0.05fF $ **FLOATING
C4961 S.t758 VSUBS 0.02fF
C4962 S.n4492 VSUBS 0.24fF $ **FLOATING
C4963 S.n4493 VSUBS 0.35fF $ **FLOATING
C4964 S.n4494 VSUBS 0.60fF $ **FLOATING
C4965 S.n4495 VSUBS 0.31fF $ **FLOATING
C4966 S.n4496 VSUBS 1.08fF $ **FLOATING
C4967 S.n4497 VSUBS 0.15fF $ **FLOATING
C4968 S.n4498 VSUBS 2.08fF $ **FLOATING
C4969 S.n4499 VSUBS 2.91fF $ **FLOATING
C4970 S.n4500 VSUBS 1.86fF $ **FLOATING
C4971 S.n4501 VSUBS 0.12fF $ **FLOATING
C4972 S.t137 VSUBS 0.02fF
C4973 S.n4502 VSUBS 0.14fF $ **FLOATING
C4974 S.t509 VSUBS 0.02fF
C4975 S.n4504 VSUBS 0.24fF $ **FLOATING
C4976 S.n4505 VSUBS 0.35fF $ **FLOATING
C4977 S.n4506 VSUBS 0.60fF $ **FLOATING
C4978 S.n4507 VSUBS 0.91fF $ **FLOATING
C4979 S.n4508 VSUBS 0.31fF $ **FLOATING
C4980 S.n4509 VSUBS 0.91fF $ **FLOATING
C4981 S.n4510 VSUBS 1.08fF $ **FLOATING
C4982 S.n4511 VSUBS 0.15fF $ **FLOATING
C4983 S.n4512 VSUBS 4.90fF $ **FLOATING
C4984 S.t528 VSUBS 0.02fF
C4985 S.n4513 VSUBS 0.12fF $ **FLOATING
C4986 S.n4514 VSUBS 0.14fF $ **FLOATING
C4987 S.t616 VSUBS 0.02fF
C4988 S.n4516 VSUBS 0.24fF $ **FLOATING
C4989 S.n4517 VSUBS 0.90fF $ **FLOATING
C4990 S.n4518 VSUBS 0.05fF $ **FLOATING
C4991 S.n4519 VSUBS 1.86fF $ **FLOATING
C4992 S.n4520 VSUBS 2.64fF $ **FLOATING
C4993 S.t852 VSUBS 0.02fF
C4994 S.n4521 VSUBS 0.24fF $ **FLOATING
C4995 S.n4522 VSUBS 0.35fF $ **FLOATING
C4996 S.n4523 VSUBS 0.60fF $ **FLOATING
C4997 S.n4524 VSUBS 0.12fF $ **FLOATING
C4998 S.t497 VSUBS 0.02fF
C4999 S.n4525 VSUBS 0.14fF $ **FLOATING
C5000 S.n4527 VSUBS 1.86fF $ **FLOATING
C5001 S.n4528 VSUBS 2.64fF $ **FLOATING
C5002 S.t1099 VSUBS 0.02fF
C5003 S.n4529 VSUBS 0.24fF $ **FLOATING
C5004 S.n4530 VSUBS 0.35fF $ **FLOATING
C5005 S.n4531 VSUBS 0.60fF $ **FLOATING
C5006 S.t115 VSUBS 0.02fF
C5007 S.n4532 VSUBS 0.24fF $ **FLOATING
C5008 S.n4533 VSUBS 0.90fF $ **FLOATING
C5009 S.n4534 VSUBS 0.05fF $ **FLOATING
C5010 S.t1125 VSUBS 0.02fF
C5011 S.n4535 VSUBS 0.12fF $ **FLOATING
C5012 S.n4536 VSUBS 0.14fF $ **FLOATING
C5013 S.n4538 VSUBS 0.12fF $ **FLOATING
C5014 S.t745 VSUBS 0.02fF
C5015 S.n4539 VSUBS 0.14fF $ **FLOATING
C5016 S.n4541 VSUBS 2.27fF $ **FLOATING
C5017 S.n4542 VSUBS 2.91fF $ **FLOATING
C5018 S.n4543 VSUBS 5.10fF $ **FLOATING
C5019 S.t871 VSUBS 0.02fF
C5020 S.n4544 VSUBS 0.12fF $ **FLOATING
C5021 S.n4545 VSUBS 0.14fF $ **FLOATING
C5022 S.t966 VSUBS 0.02fF
C5023 S.n4547 VSUBS 0.24fF $ **FLOATING
C5024 S.n4548 VSUBS 0.90fF $ **FLOATING
C5025 S.n4549 VSUBS 0.05fF $ **FLOATING
C5026 S.n4550 VSUBS 1.86fF $ **FLOATING
C5027 S.n4551 VSUBS 2.64fF $ **FLOATING
C5028 S.t75 VSUBS 0.02fF
C5029 S.n4552 VSUBS 0.24fF $ **FLOATING
C5030 S.n4553 VSUBS 0.35fF $ **FLOATING
C5031 S.n4554 VSUBS 0.60fF $ **FLOATING
C5032 S.n4555 VSUBS 0.12fF $ **FLOATING
C5033 S.t834 VSUBS 0.02fF
C5034 S.n4556 VSUBS 0.14fF $ **FLOATING
C5035 S.n4558 VSUBS 5.11fF $ **FLOATING
C5036 S.t98 VSUBS 0.02fF
C5037 S.n4559 VSUBS 0.12fF $ **FLOATING
C5038 S.n4560 VSUBS 0.14fF $ **FLOATING
C5039 S.t207 VSUBS 0.02fF
C5040 S.n4562 VSUBS 0.24fF $ **FLOATING
C5041 S.n4563 VSUBS 0.90fF $ **FLOATING
C5042 S.n4564 VSUBS 0.05fF $ **FLOATING
C5043 S.n4565 VSUBS 1.86fF $ **FLOATING
C5044 S.n4566 VSUBS 2.64fF $ **FLOATING
C5045 S.t812 VSUBS 0.02fF
C5046 S.n4567 VSUBS 0.24fF $ **FLOATING
C5047 S.n4568 VSUBS 0.35fF $ **FLOATING
C5048 S.n4569 VSUBS 0.60fF $ **FLOATING
C5049 S.n4570 VSUBS 0.12fF $ **FLOATING
C5050 S.t896 VSUBS 0.02fF
C5051 S.n4571 VSUBS 0.14fF $ **FLOATING
C5052 S.n4573 VSUBS 5.11fF $ **FLOATING
C5053 S.t514 VSUBS 0.02fF
C5054 S.n4574 VSUBS 0.12fF $ **FLOATING
C5055 S.n4575 VSUBS 0.14fF $ **FLOATING
C5056 S.t58 VSUBS 0.02fF
C5057 S.n4577 VSUBS 0.24fF $ **FLOATING
C5058 S.n4578 VSUBS 0.90fF $ **FLOATING
C5059 S.n4579 VSUBS 0.05fF $ **FLOATING
C5060 S.n4580 VSUBS 1.86fF $ **FLOATING
C5061 S.n4581 VSUBS 2.64fF $ **FLOATING
C5062 S.t20 VSUBS 0.02fF
C5063 S.n4582 VSUBS 0.24fF $ **FLOATING
C5064 S.n4583 VSUBS 0.35fF $ **FLOATING
C5065 S.n4584 VSUBS 0.60fF $ **FLOATING
C5066 S.n4585 VSUBS 0.12fF $ **FLOATING
C5067 S.t132 VSUBS 0.02fF
C5068 S.n4586 VSUBS 0.14fF $ **FLOATING
C5069 S.n4588 VSUBS 5.11fF $ **FLOATING
C5070 S.t522 VSUBS 0.02fF
C5071 S.n4589 VSUBS 0.12fF $ **FLOATING
C5072 S.n4590 VSUBS 0.14fF $ **FLOATING
C5073 S.t424 VSUBS 0.02fF
C5074 S.n4592 VSUBS 0.24fF $ **FLOATING
C5075 S.n4593 VSUBS 0.90fF $ **FLOATING
C5076 S.n4594 VSUBS 0.05fF $ **FLOATING
C5077 S.n4595 VSUBS 1.86fF $ **FLOATING
C5078 S.n4596 VSUBS 2.64fF $ **FLOATING
C5079 S.t395 VSUBS 0.02fF
C5080 S.n4597 VSUBS 0.24fF $ **FLOATING
C5081 S.n4598 VSUBS 0.35fF $ **FLOATING
C5082 S.n4599 VSUBS 0.60fF $ **FLOATING
C5083 S.n4600 VSUBS 0.12fF $ **FLOATING
C5084 S.t486 VSUBS 0.02fF
C5085 S.n4601 VSUBS 0.14fF $ **FLOATING
C5086 S.n4603 VSUBS 5.11fF $ **FLOATING
C5087 S.t864 VSUBS 0.02fF
C5088 S.n4604 VSUBS 0.12fF $ **FLOATING
C5089 S.n4605 VSUBS 0.14fF $ **FLOATING
C5090 S.t764 VSUBS 0.02fF
C5091 S.n4607 VSUBS 0.24fF $ **FLOATING
C5092 S.n4608 VSUBS 0.90fF $ **FLOATING
C5093 S.n4609 VSUBS 0.05fF $ **FLOATING
C5094 S.n4610 VSUBS 1.86fF $ **FLOATING
C5095 S.n4611 VSUBS 2.64fF $ **FLOATING
C5096 S.t736 VSUBS 0.02fF
C5097 S.n4612 VSUBS 0.24fF $ **FLOATING
C5098 S.n4613 VSUBS 0.35fF $ **FLOATING
C5099 S.n4614 VSUBS 0.60fF $ **FLOATING
C5100 S.n4615 VSUBS 0.12fF $ **FLOATING
C5101 S.t830 VSUBS 0.02fF
C5102 S.n4616 VSUBS 0.14fF $ **FLOATING
C5103 S.n4618 VSUBS 4.84fF $ **FLOATING
C5104 S.t91 VSUBS 0.02fF
C5105 S.n4619 VSUBS 0.12fF $ **FLOATING
C5106 S.n4620 VSUBS 0.14fF $ **FLOATING
C5107 S.t1106 VSUBS 0.02fF
C5108 S.n4622 VSUBS 0.24fF $ **FLOATING
C5109 S.n4623 VSUBS 0.90fF $ **FLOATING
C5110 S.n4624 VSUBS 0.05fF $ **FLOATING
C5111 S.n4625 VSUBS 1.86fF $ **FLOATING
C5112 S.n4626 VSUBS 2.64fF $ **FLOATING
C5113 S.t1072 VSUBS 0.02fF
C5114 S.n4627 VSUBS 0.24fF $ **FLOATING
C5115 S.n4628 VSUBS 0.35fF $ **FLOATING
C5116 S.n4629 VSUBS 0.60fF $ **FLOATING
C5117 S.n4630 VSUBS 0.12fF $ **FLOATING
C5118 S.t51 VSUBS 0.02fF
C5119 S.n4631 VSUBS 0.14fF $ **FLOATING
C5120 S.n4633 VSUBS 1.86fF $ **FLOATING
C5121 S.n4634 VSUBS 2.65fF $ **FLOATING
C5122 S.t1090 VSUBS 0.02fF
C5123 S.n4635 VSUBS 0.24fF $ **FLOATING
C5124 S.n4636 VSUBS 0.35fF $ **FLOATING
C5125 S.n4637 VSUBS 0.60fF $ **FLOATING
C5126 S.t181 VSUBS 0.02fF
C5127 S.n4638 VSUBS 1.20fF $ **FLOATING
C5128 S.n4639 VSUBS 0.41fF $ **FLOATING
C5129 S.n4640 VSUBS 0.44fF $ **FLOATING
C5130 S.n4641 VSUBS 0.36fF $ **FLOATING
C5131 S.n4642 VSUBS 0.20fF $ **FLOATING
C5132 S.n4643 VSUBS 0.25fF $ **FLOATING
C5133 S.n4644 VSUBS 1.27fF $ **FLOATING
C5134 S.n4645 VSUBS 1.98fF $ **FLOATING
C5135 S.n4646 VSUBS 4.03fF $ **FLOATING
C5136 S.n4647 VSUBS 0.25fF $ **FLOATING
C5137 S.n4648 VSUBS 0.01fF $ **FLOATING
C5138 S.t926 VSUBS 0.02fF
C5139 S.n4649 VSUBS 0.25fF $ **FLOATING
C5140 S.t296 VSUBS 0.02fF
C5141 S.n4650 VSUBS 0.94fF $ **FLOATING
C5142 S.n4651 VSUBS 0.70fF $ **FLOATING
C5143 S.n4652 VSUBS 0.77fF $ **FLOATING
C5144 S.n4653 VSUBS 2.24fF $ **FLOATING
C5145 S.n4654 VSUBS 1.86fF $ **FLOATING
C5146 S.n4655 VSUBS 0.12fF $ **FLOATING
C5147 S.t219 VSUBS 0.02fF
C5148 S.n4656 VSUBS 0.14fF $ **FLOATING
C5149 S.t532 VSUBS 0.02fF
C5150 S.n4658 VSUBS 0.24fF $ **FLOATING
C5151 S.n4659 VSUBS 0.35fF $ **FLOATING
C5152 S.n4660 VSUBS 0.60fF $ **FLOATING
C5153 S.n4661 VSUBS 1.37fF $ **FLOATING
C5154 S.n4662 VSUBS 0.70fF $ **FLOATING
C5155 S.n4663 VSUBS 1.13fF $ **FLOATING
C5156 S.n4664 VSUBS 0.35fF $ **FLOATING
C5157 S.n4665 VSUBS 2.00fF $ **FLOATING
C5158 S.t639 VSUBS 0.02fF
C5159 S.n4666 VSUBS 0.24fF $ **FLOATING
C5160 S.n4667 VSUBS 0.90fF $ **FLOATING
C5161 S.n4668 VSUBS 0.05fF $ **FLOATING
C5162 S.t548 VSUBS 0.02fF
C5163 S.n4669 VSUBS 0.12fF $ **FLOATING
C5164 S.n4670 VSUBS 0.14fF $ **FLOATING
C5165 S.n4672 VSUBS 1.87fF $ **FLOATING
C5166 S.n4673 VSUBS 1.86fF $ **FLOATING
C5167 S.t418 VSUBS 0.02fF
C5168 S.n4674 VSUBS 0.24fF $ **FLOATING
C5169 S.n4675 VSUBS 0.35fF $ **FLOATING
C5170 S.n4676 VSUBS 0.60fF $ **FLOATING
C5171 S.n4677 VSUBS 0.12fF $ **FLOATING
C5172 S.t32 VSUBS 0.02fF
C5173 S.n4678 VSUBS 0.14fF $ **FLOATING
C5174 S.n4680 VSUBS 1.14fF $ **FLOATING
C5175 S.n4681 VSUBS 0.22fF $ **FLOATING
C5176 S.n4682 VSUBS 0.25fF $ **FLOATING
C5177 S.n4683 VSUBS 0.09fF $ **FLOATING
C5178 S.n4684 VSUBS 1.86fF $ **FLOATING
C5179 S.t539 VSUBS 0.02fF
C5180 S.n4685 VSUBS 0.24fF $ **FLOATING
C5181 S.n4686 VSUBS 0.90fF $ **FLOATING
C5182 S.n4687 VSUBS 0.05fF $ **FLOATING
C5183 S.t945 VSUBS 0.02fF
C5184 S.n4688 VSUBS 0.12fF $ **FLOATING
C5185 S.n4689 VSUBS 0.14fF $ **FLOATING
C5186 S.n4691 VSUBS 1.86fF $ **FLOATING
C5187 S.n4692 VSUBS 2.64fF $ **FLOATING
C5188 S.t328 VSUBS 0.02fF
C5189 S.n4693 VSUBS 0.24fF $ **FLOATING
C5190 S.n4694 VSUBS 0.35fF $ **FLOATING
C5191 S.n4695 VSUBS 0.60fF $ **FLOATING
C5192 S.n4696 VSUBS 0.12fF $ **FLOATING
C5193 S.t1081 VSUBS 0.02fF
C5194 S.n4697 VSUBS 0.14fF $ **FLOATING
C5195 S.n4699 VSUBS 2.77fF $ **FLOATING
C5196 S.n4700 VSUBS 2.27fF $ **FLOATING
C5197 S.t363 VSUBS 0.02fF
C5198 S.n4701 VSUBS 0.12fF $ **FLOATING
C5199 S.n4702 VSUBS 0.14fF $ **FLOATING
C5200 S.t471 VSUBS 0.02fF
C5201 S.n4704 VSUBS 0.24fF $ **FLOATING
C5202 S.n4705 VSUBS 0.90fF $ **FLOATING
C5203 S.n4706 VSUBS 0.05fF $ **FLOATING
C5204 S.n4707 VSUBS 1.86fF $ **FLOATING
C5205 S.n4708 VSUBS 2.64fF $ **FLOATING
C5206 S.t672 VSUBS 0.02fF
C5207 S.n4709 VSUBS 0.24fF $ **FLOATING
C5208 S.n4710 VSUBS 0.35fF $ **FLOATING
C5209 S.n4711 VSUBS 0.60fF $ **FLOATING
C5210 S.n4712 VSUBS 0.12fF $ **FLOATING
C5211 S.t384 VSUBS 0.02fF
C5212 S.n4713 VSUBS 0.14fF $ **FLOATING
C5213 S.n4715 VSUBS 2.77fF $ **FLOATING
C5214 S.n4716 VSUBS 2.27fF $ **FLOATING
C5215 S.t694 VSUBS 0.02fF
C5216 S.n4717 VSUBS 0.12fF $ **FLOATING
C5217 S.n4718 VSUBS 0.14fF $ **FLOATING
C5218 S.t813 VSUBS 0.02fF
C5219 S.n4720 VSUBS 0.24fF $ **FLOATING
C5220 S.n4721 VSUBS 0.90fF $ **FLOATING
C5221 S.n4722 VSUBS 0.05fF $ **FLOATING
C5222 S.n4723 VSUBS 1.86fF $ **FLOATING
C5223 S.n4724 VSUBS 2.64fF $ **FLOATING
C5224 S.t39 VSUBS 0.02fF
C5225 S.n4725 VSUBS 0.24fF $ **FLOATING
C5226 S.n4726 VSUBS 0.35fF $ **FLOATING
C5227 S.n4727 VSUBS 0.60fF $ **FLOATING
C5228 S.n4728 VSUBS 0.12fF $ **FLOATING
C5229 S.t144 VSUBS 0.02fF
C5230 S.n4729 VSUBS 0.14fF $ **FLOATING
C5231 S.n4731 VSUBS 2.77fF $ **FLOATING
C5232 S.n4732 VSUBS 2.27fF $ **FLOATING
C5233 S.t533 VSUBS 0.02fF
C5234 S.n4733 VSUBS 0.12fF $ **FLOATING
C5235 S.n4734 VSUBS 0.14fF $ **FLOATING
C5236 S.t434 VSUBS 0.02fF
C5237 S.n4736 VSUBS 0.24fF $ **FLOATING
C5238 S.n4737 VSUBS 0.90fF $ **FLOATING
C5239 S.n4738 VSUBS 0.05fF $ **FLOATING
C5240 S.n4739 VSUBS 1.86fF $ **FLOATING
C5241 S.n4740 VSUBS 2.64fF $ **FLOATING
C5242 S.t411 VSUBS 0.02fF
C5243 S.n4741 VSUBS 0.24fF $ **FLOATING
C5244 S.n4742 VSUBS 0.35fF $ **FLOATING
C5245 S.n4743 VSUBS 0.60fF $ **FLOATING
C5246 S.n4744 VSUBS 0.12fF $ **FLOATING
C5247 S.t502 VSUBS 0.02fF
C5248 S.n4745 VSUBS 0.14fF $ **FLOATING
C5249 S.n4747 VSUBS 2.77fF $ **FLOATING
C5250 S.n4748 VSUBS 2.27fF $ **FLOATING
C5251 S.t877 VSUBS 0.02fF
C5252 S.n4749 VSUBS 0.12fF $ **FLOATING
C5253 S.n4750 VSUBS 0.14fF $ **FLOATING
C5254 S.t775 VSUBS 0.02fF
C5255 S.n4752 VSUBS 0.24fF $ **FLOATING
C5256 S.n4753 VSUBS 0.90fF $ **FLOATING
C5257 S.n4754 VSUBS 0.05fF $ **FLOATING
C5258 S.n4755 VSUBS 1.86fF $ **FLOATING
C5259 S.n4756 VSUBS 2.64fF $ **FLOATING
C5260 S.t751 VSUBS 0.02fF
C5261 S.n4757 VSUBS 0.24fF $ **FLOATING
C5262 S.n4758 VSUBS 0.35fF $ **FLOATING
C5263 S.n4759 VSUBS 0.60fF $ **FLOATING
C5264 S.n4760 VSUBS 0.12fF $ **FLOATING
C5265 S.t842 VSUBS 0.02fF
C5266 S.n4761 VSUBS 0.14fF $ **FLOATING
C5267 S.n4763 VSUBS 2.77fF $ **FLOATING
C5268 S.n4764 VSUBS 2.27fF $ **FLOATING
C5269 S.t104 VSUBS 0.02fF
C5270 S.n4765 VSUBS 0.12fF $ **FLOATING
C5271 S.n4766 VSUBS 0.14fF $ **FLOATING
C5272 S.t1120 VSUBS 0.02fF
C5273 S.n4768 VSUBS 0.24fF $ **FLOATING
C5274 S.n4769 VSUBS 0.90fF $ **FLOATING
C5275 S.n4770 VSUBS 0.05fF $ **FLOATING
C5276 S.n4771 VSUBS 0.12fF $ **FLOATING
C5277 S.t288 VSUBS 0.02fF
C5278 S.n4772 VSUBS 0.14fF $ **FLOATING
C5279 S.t232 VSUBS 0.02fF
C5280 S.n4774 VSUBS 0.24fF $ **FLOATING
C5281 S.n4775 VSUBS 0.35fF $ **FLOATING
C5282 S.n4776 VSUBS 0.60fF $ **FLOATING
C5283 S.n4777 VSUBS 1.58fF $ **FLOATING
C5284 S.n4778 VSUBS 0.03fF $ **FLOATING
C5285 S.n4779 VSUBS 0.14fF $ **FLOATING
C5286 S.n4780 VSUBS 0.58fF $ **FLOATING
C5287 S.n4781 VSUBS 0.12fF $ **FLOATING
C5288 S.n4782 VSUBS 0.53fF $ **FLOATING
C5289 S.n4783 VSUBS 0.41fF $ **FLOATING
C5290 S.n4784 VSUBS 0.24fF $ **FLOATING
C5291 S.n4785 VSUBS 0.24fF $ **FLOATING
C5292 S.n4786 VSUBS 0.67fF $ **FLOATING
C5293 S.n4787 VSUBS 1.95fF $ **FLOATING
C5294 S.t803 VSUBS 0.02fF
C5295 S.n4788 VSUBS 0.12fF $ **FLOATING
C5296 S.n4789 VSUBS 0.14fF $ **FLOATING
C5297 S.t858 VSUBS 0.02fF
C5298 S.n4791 VSUBS 0.24fF $ **FLOATING
C5299 S.n4792 VSUBS 0.90fF $ **FLOATING
C5300 S.n4793 VSUBS 0.05fF $ **FLOATING
C5301 S.t31 VSUBS 32.33fF
C5302 S.t351 VSUBS 0.02fF
C5303 S.n4794 VSUBS 0.24fF $ **FLOATING
C5304 S.n4795 VSUBS 0.90fF $ **FLOATING
C5305 S.n4796 VSUBS 0.05fF $ **FLOATING
C5306 S.t465 VSUBS 0.02fF
C5307 S.n4797 VSUBS 0.12fF $ **FLOATING
C5308 S.n4798 VSUBS 0.14fF $ **FLOATING
C5309 S.n4800 VSUBS 0.12fF $ **FLOATING
C5310 S.t68 VSUBS 0.02fF
C5311 S.n4801 VSUBS 0.14fF $ **FLOATING
C5312 S.n4803 VSUBS 5.11fF $ **FLOATING
C5313 S.n4804 VSUBS 5.38fF $ **FLOATING
C5314 S.t455 VSUBS 0.02fF
C5315 S.n4805 VSUBS 0.12fF $ **FLOATING
C5316 S.n4806 VSUBS 0.14fF $ **FLOATING
C5317 S.t340 VSUBS 0.02fF
C5318 S.n4808 VSUBS 0.24fF $ **FLOATING
C5319 S.n4809 VSUBS 0.90fF $ **FLOATING
C5320 S.n4810 VSUBS 0.05fF $ **FLOATING
C5321 S.t50 VSUBS 31.95fF
C5322 S.t899 VSUBS 0.02fF
C5323 S.n4811 VSUBS 0.01fF $ **FLOATING
C5324 S.n4812 VSUBS 0.25fF $ **FLOATING
C5325 S.t1029 VSUBS 0.02fF
C5326 S.n4814 VSUBS 1.18fF $ **FLOATING
C5327 S.n4815 VSUBS 0.05fF $ **FLOATING
C5328 S.t914 VSUBS 0.02fF
C5329 S.n4816 VSUBS 0.63fF $ **FLOATING
C5330 S.n4817 VSUBS 0.60fF $ **FLOATING
C5331 S.n4818 VSUBS 0.56fF $ **FLOATING
C5332 S.n4819 VSUBS 0.03fF $ **FLOATING
C5333 S.n4820 VSUBS 0.85fF $ **FLOATING
C5334 S.n4821 VSUBS 0.22fF $ **FLOATING
C5335 S.n4822 VSUBS 0.14fF $ **FLOATING
C5336 S.n4823 VSUBS 0.76fF $ **FLOATING
C5337 S.n4824 VSUBS 0.27fF $ **FLOATING
C5338 S.n4825 VSUBS 3.96fF $ **FLOATING
C5339 S.n4826 VSUBS 1.13fF $ **FLOATING
C5340 S.n4827 VSUBS 0.02fF $ **FLOATING
C5341 S.n4828 VSUBS 0.03fF $ **FLOATING
C5342 S.n4829 VSUBS 0.24fF $ **FLOATING
C5343 S.n4830 VSUBS 0.13fF $ **FLOATING
C5344 S.n4831 VSUBS 4.33fF $ **FLOATING
C5345 S.n4832 VSUBS 1.87fF $ **FLOATING
C5346 S.n4833 VSUBS 0.06fF $ **FLOATING
C5347 S.n4834 VSUBS 0.03fF $ **FLOATING
C5348 S.n4835 VSUBS 0.03fF $ **FLOATING
C5349 S.n4836 VSUBS 0.98fF $ **FLOATING
C5350 S.n4837 VSUBS 0.02fF $ **FLOATING
C5351 S.n4838 VSUBS 0.01fF $ **FLOATING
C5352 S.n4839 VSUBS 0.02fF $ **FLOATING
C5353 S.n4840 VSUBS 0.08fF $ **FLOATING
C5354 S.n4841 VSUBS 0.36fF $ **FLOATING
C5355 S.n4842 VSUBS 1.83fF $ **FLOATING
C5356 S.t65 VSUBS 0.02fF
C5357 S.n4843 VSUBS 0.24fF $ **FLOATING
C5358 S.n4844 VSUBS 0.35fF $ **FLOATING
C5359 S.n4845 VSUBS 0.60fF $ **FLOATING
C5360 S.n4846 VSUBS 0.12fF $ **FLOATING
C5361 S.t827 VSUBS 0.02fF
C5362 S.n4847 VSUBS 0.14fF $ **FLOATING
C5363 S.n4849 VSUBS 0.69fF $ **FLOATING
C5364 S.n4850 VSUBS 0.22fF $ **FLOATING
C5365 S.n4851 VSUBS 0.22fF $ **FLOATING
C5366 S.n4852 VSUBS 0.69fF $ **FLOATING
C5367 S.n4853 VSUBS 1.14fF $ **FLOATING
C5368 S.n4854 VSUBS 0.22fF $ **FLOATING
C5369 S.n4855 VSUBS 0.25fF $ **FLOATING
C5370 S.n4856 VSUBS 0.09fF $ **FLOATING
C5371 S.n4857 VSUBS 1.86fF $ **FLOATING
C5372 S.t196 VSUBS 0.02fF
C5373 S.n4858 VSUBS 0.24fF $ **FLOATING
C5374 S.n4859 VSUBS 0.90fF $ **FLOATING
C5375 S.n4860 VSUBS 0.05fF $ **FLOATING
C5376 S.t89 VSUBS 0.02fF
C5377 S.n4861 VSUBS 0.12fF $ **FLOATING
C5378 S.n4862 VSUBS 0.14fF $ **FLOATING
C5379 S.n4864 VSUBS 0.09fF $ **FLOATING
C5380 S.n4865 VSUBS 0.20fF $ **FLOATING
C5381 S.n4866 VSUBS 0.07fF $ **FLOATING
C5382 S.n4867 VSUBS 0.06fF $ **FLOATING
C5383 S.n4868 VSUBS 0.07fF $ **FLOATING
C5384 S.n4869 VSUBS 0.18fF $ **FLOATING
C5385 S.n4870 VSUBS 0.19fF $ **FLOATING
C5386 S.n4871 VSUBS 1.02fF $ **FLOATING
C5387 S.n4872 VSUBS 0.53fF $ **FLOATING
C5388 S.n4873 VSUBS 2.31fF $ **FLOATING
C5389 S.n4874 VSUBS 0.12fF $ **FLOATING
C5390 S.t430 VSUBS 0.02fF
C5391 S.n4875 VSUBS 0.14fF $ **FLOATING
C5392 S.t785 VSUBS 0.02fF
C5393 S.n4877 VSUBS 0.24fF $ **FLOATING
C5394 S.n4878 VSUBS 0.35fF $ **FLOATING
C5395 S.n4879 VSUBS 0.60fF $ **FLOATING
C5396 S.n4880 VSUBS 1.71fF $ **FLOATING
C5397 S.n4881 VSUBS 2.41fF $ **FLOATING
C5398 S.t807 VSUBS 0.02fF
C5399 S.n4882 VSUBS 0.12fF $ **FLOATING
C5400 S.n4883 VSUBS 0.14fF $ **FLOATING
C5401 S.t909 VSUBS 0.02fF
C5402 S.n4885 VSUBS 0.24fF $ **FLOATING
C5403 S.n4886 VSUBS 0.90fF $ **FLOATING
C5404 S.n4887 VSUBS 0.05fF $ **FLOATING
C5405 S.n4888 VSUBS 2.91fF $ **FLOATING
C5406 S.n4889 VSUBS 1.86fF $ **FLOATING
C5407 S.n4890 VSUBS 0.12fF $ **FLOATING
C5408 S.t642 VSUBS 0.02fF
C5409 S.n4891 VSUBS 0.14fF $ **FLOATING
C5410 S.t1002 VSUBS 0.02fF
C5411 S.n4893 VSUBS 0.24fF $ **FLOATING
C5412 S.n4894 VSUBS 0.35fF $ **FLOATING
C5413 S.n4895 VSUBS 0.60fF $ **FLOATING
C5414 S.n4896 VSUBS 0.91fF $ **FLOATING
C5415 S.n4897 VSUBS 0.31fF $ **FLOATING
C5416 S.n4898 VSUBS 0.91fF $ **FLOATING
C5417 S.n4899 VSUBS 1.08fF $ **FLOATING
C5418 S.n4900 VSUBS 0.15fF $ **FLOATING
C5419 S.n4901 VSUBS 4.90fF $ **FLOATING
C5420 S.t1024 VSUBS 0.02fF
C5421 S.n4902 VSUBS 0.12fF $ **FLOATING
C5422 S.n4903 VSUBS 0.14fF $ **FLOATING
C5423 S.t1139 VSUBS 0.02fF
C5424 S.n4905 VSUBS 0.24fF $ **FLOATING
C5425 S.n4906 VSUBS 0.90fF $ **FLOATING
C5426 S.n4907 VSUBS 0.05fF $ **FLOATING
C5427 S.n4908 VSUBS 1.86fF $ **FLOATING
C5428 S.n4909 VSUBS 2.64fF $ **FLOATING
C5429 S.t241 VSUBS 0.02fF
C5430 S.n4910 VSUBS 0.24fF $ **FLOATING
C5431 S.n4911 VSUBS 0.35fF $ **FLOATING
C5432 S.n4912 VSUBS 0.60fF $ **FLOATING
C5433 S.n4913 VSUBS 0.12fF $ **FLOATING
C5434 S.t989 VSUBS 0.02fF
C5435 S.n4914 VSUBS 0.14fF $ **FLOATING
C5436 S.n4916 VSUBS 2.91fF $ **FLOATING
C5437 S.n4917 VSUBS 5.10fF $ **FLOATING
C5438 S.t260 VSUBS 0.02fF
C5439 S.n4918 VSUBS 0.12fF $ **FLOATING
C5440 S.n4919 VSUBS 0.14fF $ **FLOATING
C5441 S.t377 VSUBS 0.02fF
C5442 S.n4921 VSUBS 0.24fF $ **FLOATING
C5443 S.n4922 VSUBS 0.90fF $ **FLOATING
C5444 S.n4923 VSUBS 0.05fF $ **FLOATING
C5445 S.n4924 VSUBS 1.86fF $ **FLOATING
C5446 S.n4925 VSUBS 2.64fF $ **FLOATING
C5447 S.t593 VSUBS 0.02fF
C5448 S.n4926 VSUBS 0.24fF $ **FLOATING
C5449 S.n4927 VSUBS 0.35fF $ **FLOATING
C5450 S.n4928 VSUBS 0.60fF $ **FLOATING
C5451 S.n4929 VSUBS 0.12fF $ **FLOATING
C5452 S.t230 VSUBS 0.02fF
C5453 S.n4930 VSUBS 0.14fF $ **FLOATING
C5454 S.n4932 VSUBS 5.11fF $ **FLOATING
C5455 S.t610 VSUBS 0.02fF
C5456 S.n4933 VSUBS 0.12fF $ **FLOATING
C5457 S.n4934 VSUBS 0.14fF $ **FLOATING
C5458 S.t716 VSUBS 0.02fF
C5459 S.n4936 VSUBS 0.24fF $ **FLOATING
C5460 S.n4937 VSUBS 0.90fF $ **FLOATING
C5461 S.n4938 VSUBS 0.05fF $ **FLOATING
C5462 S.n4939 VSUBS 1.86fF $ **FLOATING
C5463 S.n4940 VSUBS 2.64fF $ **FLOATING
C5464 S.t938 VSUBS 0.02fF
C5465 S.n4941 VSUBS 0.24fF $ **FLOATING
C5466 S.n4942 VSUBS 0.35fF $ **FLOATING
C5467 S.n4943 VSUBS 0.60fF $ **FLOATING
C5468 S.n4944 VSUBS 0.12fF $ **FLOATING
C5469 S.t577 VSUBS 0.02fF
C5470 S.n4945 VSUBS 0.14fF $ **FLOATING
C5471 S.n4947 VSUBS 5.11fF $ **FLOATING
C5472 S.t957 VSUBS 0.02fF
C5473 S.n4948 VSUBS 0.12fF $ **FLOATING
C5474 S.n4949 VSUBS 0.14fF $ **FLOATING
C5475 S.t1052 VSUBS 0.02fF
C5476 S.n4951 VSUBS 0.24fF $ **FLOATING
C5477 S.n4952 VSUBS 0.90fF $ **FLOATING
C5478 S.n4953 VSUBS 0.05fF $ **FLOATING
C5479 S.n4954 VSUBS 1.86fF $ **FLOATING
C5480 S.n4955 VSUBS 2.64fF $ **FLOATING
C5481 S.t57 VSUBS 0.02fF
C5482 S.n4956 VSUBS 0.24fF $ **FLOATING
C5483 S.n4957 VSUBS 0.35fF $ **FLOATING
C5484 S.n4958 VSUBS 0.60fF $ **FLOATING
C5485 S.n4959 VSUBS 0.12fF $ **FLOATING
C5486 S.t158 VSUBS 0.02fF
C5487 S.n4960 VSUBS 0.14fF $ **FLOATING
C5488 S.n4962 VSUBS 5.11fF $ **FLOATING
C5489 S.t243 VSUBS 0.02fF
C5490 S.n4963 VSUBS 0.12fF $ **FLOATING
C5491 S.n4964 VSUBS 0.14fF $ **FLOATING
C5492 S.t448 VSUBS 0.02fF
C5493 S.n4966 VSUBS 0.24fF $ **FLOATING
C5494 S.n4967 VSUBS 0.90fF $ **FLOATING
C5495 S.n4968 VSUBS 0.05fF $ **FLOATING
C5496 S.n4969 VSUBS 1.86fF $ **FLOATING
C5497 S.n4970 VSUBS 2.64fF $ **FLOATING
C5498 S.t423 VSUBS 0.02fF
C5499 S.n4971 VSUBS 0.24fF $ **FLOATING
C5500 S.n4972 VSUBS 0.35fF $ **FLOATING
C5501 S.n4973 VSUBS 0.60fF $ **FLOATING
C5502 S.n4974 VSUBS 0.12fF $ **FLOATING
C5503 S.t511 VSUBS 0.02fF
C5504 S.n4975 VSUBS 0.14fF $ **FLOATING
C5505 S.n4977 VSUBS 5.11fF $ **FLOATING
C5506 S.t886 VSUBS 0.02fF
C5507 S.n4978 VSUBS 0.12fF $ **FLOATING
C5508 S.n4979 VSUBS 0.14fF $ **FLOATING
C5509 S.t789 VSUBS 0.02fF
C5510 S.n4981 VSUBS 0.24fF $ **FLOATING
C5511 S.n4982 VSUBS 0.90fF $ **FLOATING
C5512 S.n4983 VSUBS 0.05fF $ **FLOATING
C5513 S.n4984 VSUBS 1.86fF $ **FLOATING
C5514 S.n4985 VSUBS 2.64fF $ **FLOATING
C5515 S.t763 VSUBS 0.02fF
C5516 S.n4986 VSUBS 0.24fF $ **FLOATING
C5517 S.n4987 VSUBS 0.35fF $ **FLOATING
C5518 S.n4988 VSUBS 0.60fF $ **FLOATING
C5519 S.n4989 VSUBS 0.12fF $ **FLOATING
C5520 S.t853 VSUBS 0.02fF
C5521 S.n4990 VSUBS 0.14fF $ **FLOATING
C5522 S.n4992 VSUBS 5.11fF $ **FLOATING
C5523 S.t116 VSUBS 0.02fF
C5524 S.n4993 VSUBS 0.12fF $ **FLOATING
C5525 S.n4994 VSUBS 0.14fF $ **FLOATING
C5526 S.t1129 VSUBS 0.02fF
C5527 S.n4996 VSUBS 0.24fF $ **FLOATING
C5528 S.n4997 VSUBS 0.90fF $ **FLOATING
C5529 S.n4998 VSUBS 0.05fF $ **FLOATING
C5530 S.n4999 VSUBS 1.86fF $ **FLOATING
C5531 S.n5000 VSUBS 2.64fF $ **FLOATING
C5532 S.t1101 VSUBS 0.02fF
C5533 S.n5001 VSUBS 0.24fF $ **FLOATING
C5534 S.n5002 VSUBS 0.35fF $ **FLOATING
C5535 S.n5003 VSUBS 0.60fF $ **FLOATING
C5536 S.n5004 VSUBS 0.12fF $ **FLOATING
C5537 S.t80 VSUBS 0.02fF
C5538 S.n5005 VSUBS 0.14fF $ **FLOATING
C5539 S.n5007 VSUBS 4.84fF $ **FLOATING
C5540 S.t474 VSUBS 0.02fF
C5541 S.n5008 VSUBS 0.12fF $ **FLOATING
C5542 S.n5009 VSUBS 0.14fF $ **FLOATING
C5543 S.t370 VSUBS 0.02fF
C5544 S.n5011 VSUBS 0.24fF $ **FLOATING
C5545 S.n5012 VSUBS 0.90fF $ **FLOATING
C5546 S.n5013 VSUBS 0.05fF $ **FLOATING
C5547 S.n5014 VSUBS 0.10fF $ **FLOATING
C5548 S.n5015 VSUBS 0.12fF $ **FLOATING
C5549 S.n5016 VSUBS 0.09fF $ **FLOATING
C5550 S.n5017 VSUBS 0.12fF $ **FLOATING
C5551 S.n5018 VSUBS 0.18fF $ **FLOATING
C5552 S.n5019 VSUBS 1.86fF $ **FLOATING
C5553 S.n5020 VSUBS 0.12fF $ **FLOATING
C5554 S.t453 VSUBS 0.02fF
C5555 S.n5021 VSUBS 0.14fF $ **FLOATING
C5556 S.t1026 VSUBS 0.02fF
C5557 S.n5023 VSUBS 1.20fF $ **FLOATING
C5558 S.n5024 VSUBS 0.06fF $ **FLOATING
C5559 S.n5025 VSUBS 0.10fF $ **FLOATING
C5560 S.n5026 VSUBS 0.60fF $ **FLOATING
C5561 S.n5027 VSUBS 2.39fF $ **FLOATING
C5562 S.n5028 VSUBS 2.44fF $ **FLOATING
C5563 S.n5029 VSUBS 4.24fF $ **FLOATING
C5564 S.n5030 VSUBS 0.25fF $ **FLOATING
C5565 S.n5031 VSUBS 0.01fF $ **FLOATING
C5566 S.t667 VSUBS 0.02fF
C5567 S.n5032 VSUBS 0.25fF $ **FLOATING
C5568 S.t35 VSUBS 0.02fF
C5569 S.n5033 VSUBS 0.94fF $ **FLOATING
C5570 S.n5034 VSUBS 0.70fF $ **FLOATING
C5571 S.n5035 VSUBS 1.87fF $ **FLOATING
C5572 S.n5036 VSUBS 1.86fF $ **FLOATING
C5573 S.t263 VSUBS 0.02fF
C5574 S.n5037 VSUBS 0.24fF $ **FLOATING
C5575 S.n5038 VSUBS 0.35fF $ **FLOATING
C5576 S.n5039 VSUBS 0.60fF $ **FLOATING
C5577 S.n5040 VSUBS 0.12fF $ **FLOATING
C5578 S.t1066 VSUBS 0.02fF
C5579 S.n5041 VSUBS 0.14fF $ **FLOATING
C5580 S.n5043 VSUBS 1.14fF $ **FLOATING
C5581 S.n5044 VSUBS 0.22fF $ **FLOATING
C5582 S.n5045 VSUBS 0.25fF $ **FLOATING
C5583 S.n5046 VSUBS 0.09fF $ **FLOATING
C5584 S.n5047 VSUBS 1.86fF $ **FLOATING
C5585 S.t406 VSUBS 0.02fF
C5586 S.n5048 VSUBS 0.24fF $ **FLOATING
C5587 S.n5049 VSUBS 0.90fF $ **FLOATING
C5588 S.n5050 VSUBS 0.05fF $ **FLOATING
C5589 S.t286 VSUBS 0.02fF
C5590 S.n5051 VSUBS 0.12fF $ **FLOATING
C5591 S.n5052 VSUBS 0.14fF $ **FLOATING
C5592 S.n5054 VSUBS 0.76fF $ **FLOATING
C5593 S.n5055 VSUBS 0.44fF $ **FLOATING
C5594 S.n5056 VSUBS 1.58fF $ **FLOATING
C5595 S.n5057 VSUBS 0.12fF $ **FLOATING
C5596 S.t203 VSUBS 0.02fF
C5597 S.n5058 VSUBS 0.14fF $ **FLOATING
C5598 S.t113 VSUBS 0.02fF
C5599 S.n5060 VSUBS 0.24fF $ **FLOATING
C5600 S.n5061 VSUBS 0.35fF $ **FLOATING
C5601 S.n5062 VSUBS 0.60fF $ **FLOATING
C5602 S.n5063 VSUBS 0.01fF $ **FLOATING
C5603 S.n5064 VSUBS 0.07fF $ **FLOATING
C5604 S.n5065 VSUBS 0.01fF $ **FLOATING
C5605 S.n5066 VSUBS 0.01fF $ **FLOATING
C5606 S.n5067 VSUBS 0.01fF $ **FLOATING
C5607 S.n5068 VSUBS 0.24fF $ **FLOATING
C5608 S.n5069 VSUBS 1.15fF $ **FLOATING
C5609 S.n5070 VSUBS 1.33fF $ **FLOATING
C5610 S.n5071 VSUBS 1.97fF $ **FLOATING
C5611 S.t729 VSUBS 0.02fF
C5612 S.n5072 VSUBS 0.24fF $ **FLOATING
C5613 S.n5073 VSUBS 0.90fF $ **FLOATING
C5614 S.n5074 VSUBS 0.05fF $ **FLOATING
C5615 S.t45 VSUBS 0.02fF
C5616 S.n5075 VSUBS 0.12fF $ **FLOATING
C5617 S.n5076 VSUBS 0.14fF $ **FLOATING
C5618 S.n5078 VSUBS 1.86fF $ **FLOATING
C5619 S.n5079 VSUBS 0.12fF $ **FLOATING
C5620 S.t910 VSUBS 0.02fF
C5621 S.n5080 VSUBS 0.14fF $ **FLOATING
C5622 S.t160 VSUBS 0.02fF
C5623 S.n5082 VSUBS 0.24fF $ **FLOATING
C5624 S.n5083 VSUBS 0.35fF $ **FLOATING
C5625 S.n5084 VSUBS 0.60fF $ **FLOATING
C5626 S.n5085 VSUBS 0.31fF $ **FLOATING
C5627 S.n5086 VSUBS 1.08fF $ **FLOATING
C5628 S.n5087 VSUBS 0.15fF $ **FLOATING
C5629 S.n5088 VSUBS 2.08fF $ **FLOATING
C5630 S.t686 VSUBS 0.02fF
C5631 S.n5089 VSUBS 0.12fF $ **FLOATING
C5632 S.n5090 VSUBS 0.14fF $ **FLOATING
C5633 S.t273 VSUBS 0.02fF
C5634 S.n5092 VSUBS 0.24fF $ **FLOATING
C5635 S.n5093 VSUBS 0.90fF $ **FLOATING
C5636 S.n5094 VSUBS 0.05fF $ **FLOATING
C5637 S.n5095 VSUBS 1.86fF $ **FLOATING
C5638 S.n5096 VSUBS 2.64fF $ **FLOATING
C5639 S.t512 VSUBS 0.02fF
C5640 S.n5097 VSUBS 0.24fF $ **FLOATING
C5641 S.n5098 VSUBS 0.35fF $ **FLOATING
C5642 S.n5099 VSUBS 0.60fF $ **FLOATING
C5643 S.n5100 VSUBS 0.12fF $ **FLOATING
C5644 S.t143 VSUBS 0.02fF
C5645 S.n5101 VSUBS 0.14fF $ **FLOATING
C5646 S.n5103 VSUBS 2.27fF $ **FLOATING
C5647 S.t534 VSUBS 0.02fF
C5648 S.n5104 VSUBS 0.12fF $ **FLOATING
C5649 S.n5105 VSUBS 0.14fF $ **FLOATING
C5650 S.t619 VSUBS 0.02fF
C5651 S.n5107 VSUBS 0.24fF $ **FLOATING
C5652 S.n5108 VSUBS 0.90fF $ **FLOATING
C5653 S.n5109 VSUBS 0.05fF $ **FLOATING
C5654 S.n5110 VSUBS 1.86fF $ **FLOATING
C5655 S.n5111 VSUBS 2.64fF $ **FLOATING
C5656 S.t855 VSUBS 0.02fF
C5657 S.n5112 VSUBS 0.24fF $ **FLOATING
C5658 S.n5113 VSUBS 0.35fF $ **FLOATING
C5659 S.n5114 VSUBS 0.60fF $ **FLOATING
C5660 S.n5115 VSUBS 0.12fF $ **FLOATING
C5661 S.t504 VSUBS 0.02fF
C5662 S.n5116 VSUBS 0.14fF $ **FLOATING
C5663 S.n5118 VSUBS 2.77fF $ **FLOATING
C5664 S.n5119 VSUBS 2.27fF $ **FLOATING
C5665 S.t876 VSUBS 0.02fF
C5666 S.n5120 VSUBS 0.12fF $ **FLOATING
C5667 S.n5121 VSUBS 0.14fF $ **FLOATING
C5668 S.t970 VSUBS 0.02fF
C5669 S.n5123 VSUBS 0.24fF $ **FLOATING
C5670 S.n5124 VSUBS 0.90fF $ **FLOATING
C5671 S.n5125 VSUBS 0.05fF $ **FLOATING
C5672 S.n5126 VSUBS 1.86fF $ **FLOATING
C5673 S.n5127 VSUBS 2.64fF $ **FLOATING
C5674 S.t81 VSUBS 0.02fF
C5675 S.n5128 VSUBS 0.24fF $ **FLOATING
C5676 S.n5129 VSUBS 0.35fF $ **FLOATING
C5677 S.n5130 VSUBS 0.60fF $ **FLOATING
C5678 S.n5131 VSUBS 0.12fF $ **FLOATING
C5679 S.t838 VSUBS 0.02fF
C5680 S.n5132 VSUBS 0.14fF $ **FLOATING
C5681 S.n5134 VSUBS 2.77fF $ **FLOATING
C5682 S.n5135 VSUBS 2.27fF $ **FLOATING
C5683 S.t106 VSUBS 0.02fF
C5684 S.n5136 VSUBS 0.12fF $ **FLOATING
C5685 S.n5137 VSUBS 0.14fF $ **FLOATING
C5686 S.t210 VSUBS 0.02fF
C5687 S.n5139 VSUBS 0.24fF $ **FLOATING
C5688 S.n5140 VSUBS 0.90fF $ **FLOATING
C5689 S.n5141 VSUBS 0.05fF $ **FLOATING
C5690 S.n5142 VSUBS 1.86fF $ **FLOATING
C5691 S.n5143 VSUBS 2.64fF $ **FLOATING
C5692 S.t444 VSUBS 0.02fF
C5693 S.n5144 VSUBS 0.24fF $ **FLOATING
C5694 S.n5145 VSUBS 0.35fF $ **FLOATING
C5695 S.n5146 VSUBS 0.60fF $ **FLOATING
C5696 S.n5147 VSUBS 0.12fF $ **FLOATING
C5697 S.t121 VSUBS 0.02fF
C5698 S.n5148 VSUBS 0.14fF $ **FLOATING
C5699 S.n5150 VSUBS 2.77fF $ **FLOATING
C5700 S.n5151 VSUBS 2.27fF $ **FLOATING
C5701 S.t461 VSUBS 0.02fF
C5702 S.n5152 VSUBS 0.12fF $ **FLOATING
C5703 S.n5153 VSUBS 0.14fF $ **FLOATING
C5704 S.t559 VSUBS 0.02fF
C5705 S.n5155 VSUBS 0.24fF $ **FLOATING
C5706 S.n5156 VSUBS 0.90fF $ **FLOATING
C5707 S.n5157 VSUBS 0.05fF $ **FLOATING
C5708 S.n5158 VSUBS 1.86fF $ **FLOATING
C5709 S.n5159 VSUBS 2.64fF $ **FLOATING
C5710 S.t431 VSUBS 0.02fF
C5711 S.n5160 VSUBS 0.24fF $ **FLOATING
C5712 S.n5161 VSUBS 0.35fF $ **FLOATING
C5713 S.n5162 VSUBS 0.60fF $ **FLOATING
C5714 S.n5163 VSUBS 0.12fF $ **FLOATING
C5715 S.t519 VSUBS 0.02fF
C5716 S.n5164 VSUBS 0.14fF $ **FLOATING
C5717 S.n5166 VSUBS 2.77fF $ **FLOATING
C5718 S.n5167 VSUBS 2.27fF $ **FLOATING
C5719 S.t894 VSUBS 0.02fF
C5720 S.n5168 VSUBS 0.12fF $ **FLOATING
C5721 S.n5169 VSUBS 0.14fF $ **FLOATING
C5722 S.t796 VSUBS 0.02fF
C5723 S.n5171 VSUBS 0.24fF $ **FLOATING
C5724 S.n5172 VSUBS 0.90fF $ **FLOATING
C5725 S.n5173 VSUBS 0.05fF $ **FLOATING
C5726 S.n5174 VSUBS 1.86fF $ **FLOATING
C5727 S.n5175 VSUBS 2.64fF $ **FLOATING
C5728 S.t773 VSUBS 0.02fF
C5729 S.n5176 VSUBS 0.24fF $ **FLOATING
C5730 S.n5177 VSUBS 0.35fF $ **FLOATING
C5731 S.n5178 VSUBS 0.60fF $ **FLOATING
C5732 S.n5179 VSUBS 0.12fF $ **FLOATING
C5733 S.t861 VSUBS 0.02fF
C5734 S.n5180 VSUBS 0.14fF $ **FLOATING
C5735 S.n5182 VSUBS 2.77fF $ **FLOATING
C5736 S.n5183 VSUBS 2.27fF $ **FLOATING
C5737 S.t126 VSUBS 0.02fF
C5738 S.n5184 VSUBS 0.12fF $ **FLOATING
C5739 S.n5185 VSUBS 0.14fF $ **FLOATING
C5740 S.t1 VSUBS 0.02fF
C5741 S.n5187 VSUBS 0.24fF $ **FLOATING
C5742 S.n5188 VSUBS 0.90fF $ **FLOATING
C5743 S.n5189 VSUBS 0.05fF $ **FLOATING
C5744 S.n5190 VSUBS 1.86fF $ **FLOATING
C5745 S.n5191 VSUBS 2.64fF $ **FLOATING
C5746 S.t1116 VSUBS 0.02fF
C5747 S.n5192 VSUBS 0.24fF $ **FLOATING
C5748 S.n5193 VSUBS 0.35fF $ **FLOATING
C5749 S.n5194 VSUBS 0.60fF $ **FLOATING
C5750 S.n5195 VSUBS 0.12fF $ **FLOATING
C5751 S.t88 VSUBS 0.02fF
C5752 S.n5196 VSUBS 0.14fF $ **FLOATING
C5753 S.n5198 VSUBS 2.77fF $ **FLOATING
C5754 S.n5199 VSUBS 2.27fF $ **FLOATING
C5755 S.t484 VSUBS 0.02fF
C5756 S.n5200 VSUBS 0.12fF $ **FLOATING
C5757 S.n5201 VSUBS 0.14fF $ **FLOATING
C5758 S.t379 VSUBS 0.02fF
C5759 S.n5203 VSUBS 0.24fF $ **FLOATING
C5760 S.n5204 VSUBS 0.90fF $ **FLOATING
C5761 S.n5205 VSUBS 0.05fF $ **FLOATING
C5762 S.t44 VSUBS 32.33fF
C5763 S.t828 VSUBS 0.02fF
C5764 S.n5206 VSUBS 0.12fF $ **FLOATING
C5765 S.n5207 VSUBS 0.14fF $ **FLOATING
C5766 S.t719 VSUBS 0.02fF
C5767 S.n5209 VSUBS 0.24fF $ **FLOATING
C5768 S.n5210 VSUBS 0.90fF $ **FLOATING
C5769 S.n5211 VSUBS 0.05fF $ **FLOATING
C5770 S.t348 VSUBS 0.02fF
C5771 S.n5212 VSUBS 0.24fF $ **FLOATING
C5772 S.n5213 VSUBS 0.35fF $ **FLOATING
C5773 S.n5214 VSUBS 0.60fF $ **FLOATING
C5774 S.n5215 VSUBS 2.63fF $ **FLOATING
C5775 S.n5216 VSUBS 3.24fF $ **FLOATING
C5776 S.n5217 VSUBS 0.10fF $ **FLOATING
C5777 S.n5218 VSUBS 0.35fF $ **FLOATING
C5778 S.n5219 VSUBS 0.46fF $ **FLOATING
C5779 S.n5220 VSUBS 1.12fF $ **FLOATING
C5780 S.n5221 VSUBS 1.85fF $ **FLOATING
C5781 S.n5222 VSUBS 0.12fF $ **FLOATING
C5782 S.t438 VSUBS 0.02fF
C5783 S.n5223 VSUBS 0.14fF $ **FLOATING
C5784 S.t336 VSUBS 0.02fF
C5785 S.n5225 VSUBS 0.24fF $ **FLOATING
C5786 S.n5226 VSUBS 0.35fF $ **FLOATING
C5787 S.n5227 VSUBS 0.60fF $ **FLOATING
C5788 S.n5228 VSUBS 1.25fF $ **FLOATING
C5789 S.n5229 VSUBS 2.36fF $ **FLOATING
C5790 S.n5230 VSUBS 4.15fF $ **FLOATING
C5791 S.t819 VSUBS 0.02fF
C5792 S.n5231 VSUBS 0.12fF $ **FLOATING
C5793 S.n5232 VSUBS 0.14fF $ **FLOATING
C5794 S.t706 VSUBS 0.02fF
C5795 S.n5234 VSUBS 0.24fF $ **FLOATING
C5796 S.n5235 VSUBS 0.90fF $ **FLOATING
C5797 S.n5236 VSUBS 0.05fF $ **FLOATING
C5798 S.t79 VSUBS 31.95fF
C5799 S.t808 VSUBS 0.02fF
C5800 S.n5237 VSUBS 0.01fF $ **FLOATING
C5801 S.n5238 VSUBS 0.25fF $ **FLOATING
C5802 S.t792 VSUBS 0.02fF
C5803 S.n5240 VSUBS 1.18fF $ **FLOATING
C5804 S.n5241 VSUBS 0.05fF $ **FLOATING
C5805 S.t652 VSUBS 0.02fF
C5806 S.n5242 VSUBS 0.63fF $ **FLOATING
C5807 S.n5243 VSUBS 0.60fF $ **FLOATING
C5808 S.n5244 VSUBS 2.77fF $ **FLOATING
C5809 S.n5245 VSUBS 1.48fF $ **FLOATING
C5810 S.n5246 VSUBS 0.02fF $ **FLOATING
C5811 S.n5247 VSUBS 0.01fF $ **FLOATING
C5812 S.n5248 VSUBS 0.01fF $ **FLOATING
C5813 S.n5249 VSUBS 0.01fF $ **FLOATING
C5814 S.n5250 VSUBS 0.01fF $ **FLOATING
C5815 S.n5251 VSUBS 0.02fF $ **FLOATING
C5816 S.n5252 VSUBS 0.02fF $ **FLOATING
C5817 S.n5253 VSUBS 0.04fF $ **FLOATING
C5818 S.n5254 VSUBS 0.16fF $ **FLOATING
C5819 S.n5255 VSUBS 0.10fF $ **FLOATING
C5820 S.n5256 VSUBS 0.16fF $ **FLOATING
C5821 S.n5257 VSUBS 0.14fF $ **FLOATING
C5822 S.n5258 VSUBS 0.27fF $ **FLOATING
C5823 S.n5259 VSUBS 0.24fF $ **FLOATING
C5824 S.n5260 VSUBS 4.63fF $ **FLOATING
C5825 S.t496 VSUBS 0.02fF
C5826 S.n5261 VSUBS 0.88fF $ **FLOATING
C5827 S.t872 VSUBS 0.02fF
C5828 S.n5262 VSUBS 0.88fF $ **FLOATING
C5829 S.t1006 VSUBS 0.02fF
C5830 S.n5263 VSUBS 0.02fF $ **FLOATING
C5831 S.n5264 VSUBS 0.37fF $ **FLOATING
C5832 S.t903 VSUBS 0.02fF
C5833 S.n5265 VSUBS 0.88fF $ **FLOATING
C5834 S.t277 VSUBS 0.02fF
C5835 S.n5266 VSUBS 0.02fF $ **FLOATING
C5836 S.n5267 VSUBS 0.37fF $ **FLOATING
C5837 S.t527 VSUBS 0.02fF
C5838 S.n5268 VSUBS 0.88fF $ **FLOATING
C5839 S.t190 VSUBS 0.02fF
C5840 S.n5269 VSUBS 0.88fF $ **FLOATING
C5841 S.t676 VSUBS 0.02fF
C5842 S.n5270 VSUBS 0.02fF $ **FLOATING
C5843 S.n5271 VSUBS 0.37fF $ **FLOATING
C5844 S.t918 VSUBS 0.02fF
C5845 S.n5272 VSUBS 0.88fF $ **FLOATING
C5846 S.t1131 VSUBS 0.02fF
C5847 S.n5273 VSUBS 0.88fF $ **FLOATING
C5848 S.t524 VSUBS 0.02fF
C5849 S.n5274 VSUBS 0.02fF $ **FLOATING
C5850 S.n5275 VSUBS 0.37fF $ **FLOATING
C5851 S.t752 VSUBS 0.02fF
C5852 S.n5276 VSUBS 0.88fF $ **FLOATING
C5853 S.t372 VSUBS 0.02fF
C5854 S.n5277 VSUBS 0.88fF $ **FLOATING
C5855 S.t866 VSUBS 0.02fF
C5856 S.n5278 VSUBS 0.02fF $ **FLOATING
C5857 S.n5279 VSUBS 0.37fF $ **FLOATING
C5858 S.t1093 VSUBS 0.02fF
C5859 S.n5280 VSUBS 0.88fF $ **FLOATING
C5860 S.t708 VSUBS 0.02fF
C5861 S.n5281 VSUBS 0.88fF $ **FLOATING
C5862 S.t92 VSUBS 0.02fF
C5863 S.n5282 VSUBS 0.02fF $ **FLOATING
C5864 S.n5283 VSUBS 0.37fF $ **FLOATING
C5865 S.t322 VSUBS 0.02fF
C5866 S.n5284 VSUBS 0.88fF $ **FLOATING
C5867 S.t1046 VSUBS 0.02fF
C5868 S.n5285 VSUBS 0.88fF $ **FLOATING
C5869 S.t454 VSUBS 0.02fF
C5870 S.n5286 VSUBS 0.02fF $ **FLOATING
C5871 S.n5287 VSUBS 0.37fF $ **FLOATING
C5872 S.t665 VSUBS 0.02fF
C5873 S.n5288 VSUBS 0.88fF $ **FLOATING
C5874 S.t345 VSUBS 0.02fF
C5875 S.n5289 VSUBS 0.88fF $ **FLOATING
C5876 S.t744 VSUBS 0.02fF
C5877 S.n5290 VSUBS 0.02fF $ **FLOATING
C5878 S.n5291 VSUBS 0.37fF $ **FLOATING
C5879 S.t211 VSUBS 0.02fF
C5880 S.n5292 VSUBS 0.88fF $ **FLOATING
C5881 S.t939 VSUBS 0.02fF
C5882 S.n5293 VSUBS 0.88fF $ **FLOATING
C5883 S.t1080 VSUBS 0.02fF
C5884 S.n5294 VSUBS 0.02fF $ **FLOATING
C5885 S.n5295 VSUBS 0.37fF $ **FLOATING
C5886 S.t561 VSUBS 0.02fF
C5887 S.n5296 VSUBS 0.88fF $ **FLOATING
C5888 S.t178 VSUBS 0.02fF
C5889 S.n5297 VSUBS 0.88fF $ **FLOATING
C5890 S.t312 VSUBS 0.02fF
C5891 S.n5298 VSUBS 0.02fF $ **FLOATING
C5892 S.n5299 VSUBS 0.37fF $ **FLOATING
C5893 S.t906 VSUBS 0.02fF
C5894 S.n5300 VSUBS 0.88fF $ **FLOATING
C5895 S.t529 VSUBS 0.02fF
C5896 S.n5301 VSUBS 0.88fF $ **FLOATING
C5897 S.t659 VSUBS 0.02fF
C5898 S.n5302 VSUBS 0.02fF $ **FLOATING
C5899 S.n5303 VSUBS 0.37fF $ **FLOATING
C5900 S.t138 VSUBS 0.02fF
C5901 S.n5304 VSUBS 0.88fF $ **FLOATING
C5902 S.t112 VSUBS 0.02fF
C5903 S.n5305 VSUBS 0.44fF $ **FLOATING
C5904 S.t0 VSUBS 969.03fF
C5905 S.t170 VSUBS 0.02fF
C5906 S.n5306 VSUBS 1.30fF $ **FLOATING
C5907 S.n5307 VSUBS 0.24fF $ **FLOATING
C5908 S.n5308 VSUBS 6.68fF $ **FLOATING
C5909 S.n5309 VSUBS 2.89fF $ **FLOATING
C5910 S.n5310 VSUBS 0.25fF $ **FLOATING
C5911 S.n5311 VSUBS 0.09fF $ **FLOATING
C5912 S.n5312 VSUBS 0.20fF $ **FLOATING
C5913 S.n5313 VSUBS 0.77fF $ **FLOATING
C5914 S.n5314 VSUBS 1.91fF $ **FLOATING
C5915 S.n5315 VSUBS 1.86fF $ **FLOATING
C5916 S.n5316 VSUBS 0.12fF $ **FLOATING
C5917 S.t797 VSUBS 0.02fF
C5918 S.n5317 VSUBS 0.14fF $ **FLOATING
C5919 S.t702 VSUBS 0.02fF
C5920 S.n5319 VSUBS 0.24fF $ **FLOATING
C5921 S.n5320 VSUBS 0.35fF $ **FLOATING
C5922 S.n5321 VSUBS 0.60fF $ **FLOATING
C5923 S.n5322 VSUBS 2.64fF $ **FLOATING
C5924 S.n5323 VSUBS 2.96fF $ **FLOATING
C5925 S.t1069 VSUBS 0.02fF
C5926 S.n5324 VSUBS 0.24fF $ **FLOATING
C5927 S.n5325 VSUBS 0.90fF $ **FLOATING
C5928 S.n5326 VSUBS 0.05fF $ **FLOATING
C5929 S.t63 VSUBS 0.02fF
C5930 S.n5327 VSUBS 0.12fF $ **FLOATING
C5931 S.n5328 VSUBS 0.14fF $ **FLOATING
C5932 S.n5330 VSUBS 1.76fF $ **FLOATING
C5933 S.n5331 VSUBS 3.01fF $ **FLOATING
C5934 S.t538 VSUBS 0.02fF
C5935 S.n5332 VSUBS 0.24fF $ **FLOATING
C5936 S.n5333 VSUBS 0.35fF $ **FLOATING
C5937 S.n5334 VSUBS 0.60fF $ **FLOATING
C5938 S.n5335 VSUBS 0.12fF $ **FLOATING
C5939 S.t173 VSUBS 0.02fF
C5940 S.n5336 VSUBS 0.14fF $ **FLOATING
C5941 S.n5338 VSUBS 0.22fF $ **FLOATING
C5942 S.n5339 VSUBS 0.65fF $ **FLOATING
C5943 S.n5340 VSUBS 0.90fF $ **FLOATING
C5944 S.n5341 VSUBS 0.22fF $ **FLOATING
C5945 S.n5342 VSUBS 1.97fF $ **FLOATING
C5946 S.t552 VSUBS 0.02fF
C5947 S.n5343 VSUBS 0.12fF $ **FLOATING
C5948 S.n5344 VSUBS 0.14fF $ **FLOATING
C5949 S.t647 VSUBS 0.02fF
C5950 S.n5346 VSUBS 0.24fF $ **FLOATING
C5951 S.n5347 VSUBS 0.90fF $ **FLOATING
C5952 S.n5348 VSUBS 0.05fF $ **FLOATING
C5953 S.n5349 VSUBS 1.86fF $ **FLOATING
C5954 S.n5350 VSUBS 0.12fF $ **FLOATING
C5955 S.t569 VSUBS 0.02fF
C5956 S.n5351 VSUBS 0.14fF $ **FLOATING
C5957 S.t928 VSUBS 0.02fF
C5958 S.n5353 VSUBS 0.24fF $ **FLOATING
C5959 S.n5354 VSUBS 0.35fF $ **FLOATING
C5960 S.n5355 VSUBS 0.60fF $ **FLOATING
C5961 S.n5356 VSUBS 0.31fF $ **FLOATING
C5962 S.n5357 VSUBS 0.91fF $ **FLOATING
C5963 S.n5358 VSUBS 1.08fF $ **FLOATING
C5964 S.n5359 VSUBS 0.15fF $ **FLOATING
C5965 S.n5360 VSUBS 4.90fF $ **FLOATING
C5966 S.t947 VSUBS 0.02fF
C5967 S.n5361 VSUBS 0.12fF $ **FLOATING
C5968 S.n5362 VSUBS 0.14fF $ **FLOATING
C5969 S.t1042 VSUBS 0.02fF
C5970 S.n5364 VSUBS 0.24fF $ **FLOATING
C5971 S.n5365 VSUBS 0.90fF $ **FLOATING
C5972 S.n5366 VSUBS 0.05fF $ **FLOATING
C5973 S.n5367 VSUBS 1.86fF $ **FLOATING
C5974 S.n5368 VSUBS 2.64fF $ **FLOATING
C5975 S.t762 VSUBS 0.02fF
C5976 S.n5369 VSUBS 0.24fF $ **FLOATING
C5977 S.n5370 VSUBS 0.35fF $ **FLOATING
C5978 S.n5371 VSUBS 0.60fF $ **FLOATING
C5979 S.n5372 VSUBS 0.12fF $ **FLOATING
C5980 S.t407 VSUBS 0.02fF
C5981 S.n5373 VSUBS 0.14fF $ **FLOATING
C5982 S.n5375 VSUBS 5.10fF $ **FLOATING
C5983 S.t787 VSUBS 0.02fF
C5984 S.n5376 VSUBS 0.12fF $ **FLOATING
C5985 S.n5377 VSUBS 0.14fF $ **FLOATING
C5986 S.t887 VSUBS 0.02fF
C5987 S.n5379 VSUBS 0.24fF $ **FLOATING
C5988 S.n5380 VSUBS 0.90fF $ **FLOATING
C5989 S.n5381 VSUBS 0.05fF $ **FLOATING
C5990 S.n5382 VSUBS 1.86fF $ **FLOATING
C5991 S.n5383 VSUBS 2.64fF $ **FLOATING
C5992 S.t1103 VSUBS 0.02fF
C5993 S.n5384 VSUBS 0.24fF $ **FLOATING
C5994 S.n5385 VSUBS 0.35fF $ **FLOATING
C5995 S.n5386 VSUBS 0.60fF $ **FLOATING
C5996 S.n5387 VSUBS 0.12fF $ **FLOATING
C5997 S.t749 VSUBS 0.02fF
C5998 S.n5388 VSUBS 0.14fF $ **FLOATING
C5999 S.n5390 VSUBS 5.11fF $ **FLOATING
C6000 S.t1127 VSUBS 0.02fF
C6001 S.n5391 VSUBS 0.12fF $ **FLOATING
C6002 S.n5392 VSUBS 0.14fF $ **FLOATING
C6003 S.t120 VSUBS 0.02fF
C6004 S.n5394 VSUBS 0.24fF $ **FLOATING
C6005 S.n5395 VSUBS 0.90fF $ **FLOATING
C6006 S.n5396 VSUBS 0.05fF $ **FLOATING
C6007 S.n5397 VSUBS 1.86fF $ **FLOATING
C6008 S.n5398 VSUBS 2.64fF $ **FLOATING
C6009 S.t332 VSUBS 0.02fF
C6010 S.n5399 VSUBS 0.24fF $ **FLOATING
C6011 S.n5400 VSUBS 0.35fF $ **FLOATING
C6012 S.n5401 VSUBS 0.60fF $ **FLOATING
C6013 S.n5402 VSUBS 0.12fF $ **FLOATING
C6014 S.t1087 VSUBS 0.02fF
C6015 S.n5403 VSUBS 0.14fF $ **FLOATING
C6016 S.n5405 VSUBS 5.11fF $ **FLOATING
C6017 S.t368 VSUBS 0.02fF
C6018 S.n5406 VSUBS 0.12fF $ **FLOATING
C6019 S.n5407 VSUBS 0.14fF $ **FLOATING
C6020 S.t477 VSUBS 0.02fF
C6021 S.n5409 VSUBS 0.24fF $ **FLOATING
C6022 S.n5410 VSUBS 0.90fF $ **FLOATING
C6023 S.n5411 VSUBS 0.05fF $ **FLOATING
C6024 S.n5412 VSUBS 1.86fF $ **FLOATING
C6025 S.n5413 VSUBS 2.64fF $ **FLOATING
C6026 S.t679 VSUBS 0.02fF
C6027 S.n5414 VSUBS 0.24fF $ **FLOATING
C6028 S.n5415 VSUBS 0.35fF $ **FLOATING
C6029 S.n5416 VSUBS 0.60fF $ **FLOATING
C6030 S.n5417 VSUBS 0.12fF $ **FLOATING
C6031 S.t317 VSUBS 0.02fF
C6032 S.n5418 VSUBS 0.14fF $ **FLOATING
C6033 S.n5420 VSUBS 5.11fF $ **FLOATING
C6034 S.t698 VSUBS 0.02fF
C6035 S.n5421 VSUBS 0.12fF $ **FLOATING
C6036 S.n5422 VSUBS 0.14fF $ **FLOATING
C6037 S.t822 VSUBS 0.02fF
C6038 S.n5424 VSUBS 0.24fF $ **FLOATING
C6039 S.n5425 VSUBS 0.90fF $ **FLOATING
C6040 S.n5426 VSUBS 0.05fF $ **FLOATING
C6041 S.n5427 VSUBS 1.86fF $ **FLOATING
C6042 S.n5428 VSUBS 2.64fF $ **FLOATING
C6043 S.t446 VSUBS 0.02fF
C6044 S.n5429 VSUBS 0.24fF $ **FLOATING
C6045 S.n5430 VSUBS 0.35fF $ **FLOATING
C6046 S.n5431 VSUBS 0.60fF $ **FLOATING
C6047 S.n5432 VSUBS 0.12fF $ **FLOATING
C6048 S.t531 VSUBS 0.02fF
C6049 S.n5433 VSUBS 0.14fF $ **FLOATING
C6050 S.n5435 VSUBS 5.11fF $ **FLOATING
C6051 S.t1111 VSUBS 0.02fF
C6052 S.n5436 VSUBS 0.12fF $ **FLOATING
C6053 S.n5437 VSUBS 0.14fF $ **FLOATING
C6054 S.t809 VSUBS 0.02fF
C6055 S.n5439 VSUBS 0.24fF $ **FLOATING
C6056 S.n5440 VSUBS 0.90fF $ **FLOATING
C6057 S.n5441 VSUBS 0.05fF $ **FLOATING
C6058 S.n5442 VSUBS 1.86fF $ **FLOATING
C6059 S.n5443 VSUBS 2.64fF $ **FLOATING
C6060 S.t786 VSUBS 0.02fF
C6061 S.n5444 VSUBS 0.24fF $ **FLOATING
C6062 S.n5445 VSUBS 0.35fF $ **FLOATING
C6063 S.n5446 VSUBS 0.60fF $ **FLOATING
C6064 S.n5447 VSUBS 0.12fF $ **FLOATING
C6065 S.t875 VSUBS 0.02fF
C6066 S.n5448 VSUBS 0.14fF $ **FLOATING
C6067 S.n5450 VSUBS 5.11fF $ **FLOATING
C6068 S.t142 VSUBS 0.02fF
C6069 S.n5451 VSUBS 0.12fF $ **FLOATING
C6070 S.n5452 VSUBS 0.14fF $ **FLOATING
C6071 S.t18 VSUBS 0.02fF
C6072 S.n5454 VSUBS 0.24fF $ **FLOATING
C6073 S.n5455 VSUBS 0.90fF $ **FLOATING
C6074 S.n5456 VSUBS 0.05fF $ **FLOATING
C6075 S.n5457 VSUBS 1.86fF $ **FLOATING
C6076 S.n5458 VSUBS 2.64fF $ **FLOATING
C6077 S.t1128 VSUBS 0.02fF
C6078 S.n5459 VSUBS 0.24fF $ **FLOATING
C6079 S.n5460 VSUBS 0.35fF $ **FLOATING
C6080 S.n5461 VSUBS 0.60fF $ **FLOATING
C6081 S.n5462 VSUBS 0.12fF $ **FLOATING
C6082 S.t101 VSUBS 0.02fF
C6083 S.n5463 VSUBS 0.14fF $ **FLOATING
C6084 S.n5465 VSUBS 5.11fF $ **FLOATING
C6085 S.t499 VSUBS 0.02fF
C6086 S.n5466 VSUBS 0.12fF $ **FLOATING
C6087 S.n5467 VSUBS 0.14fF $ **FLOATING
C6088 S.t394 VSUBS 0.02fF
C6089 S.n5469 VSUBS 0.24fF $ **FLOATING
C6090 S.n5470 VSUBS 0.90fF $ **FLOATING
C6091 S.n5471 VSUBS 0.05fF $ **FLOATING
C6092 S.n5472 VSUBS 0.35fF $ **FLOATING
C6093 S.n5473 VSUBS 0.46fF $ **FLOATING
C6094 S.n5474 VSUBS 1.12fF $ **FLOATING
C6095 S.n5475 VSUBS 1.86fF $ **FLOATING
C6096 S.n5476 VSUBS 0.12fF $ **FLOATING
C6097 S.t460 VSUBS 0.02fF
C6098 S.n5477 VSUBS 0.14fF $ **FLOATING
C6099 S.t366 VSUBS 0.02fF
C6100 S.n5479 VSUBS 0.24fF $ **FLOATING
C6101 S.n5480 VSUBS 0.35fF $ **FLOATING
C6102 S.n5481 VSUBS 0.60fF $ **FLOATING
C6103 S.n5482 VSUBS 2.64fF $ **FLOATING
C6104 S.n5483 VSUBS 3.88fF $ **FLOATING
C6105 S.t837 VSUBS 0.02fF
C6106 S.n5484 VSUBS 0.12fF $ **FLOATING
C6107 S.n5485 VSUBS 0.14fF $ **FLOATING
C6108 S.t732 VSUBS 0.02fF
C6109 S.n5487 VSUBS 0.24fF $ **FLOATING
C6110 S.n5488 VSUBS 0.90fF $ **FLOATING
C6111 S.n5489 VSUBS 0.05fF $ **FLOATING
C6112 S.t62 VSUBS 31.95fF
C6113 S.t703 VSUBS 0.02fF
C6114 S.n5490 VSUBS 0.01fF $ **FLOATING
C6115 S.n5491 VSUBS 0.25fF $ **FLOATING
C6116 S.t541 VSUBS 0.02fF
C6117 S.n5493 VSUBS 1.18fF $ **FLOATING
C6118 S.n5494 VSUBS 0.05fF $ **FLOATING
C6119 S.t421 VSUBS 0.02fF
C6120 S.n5495 VSUBS 0.63fF $ **FLOATING
C6121 S.n5496 VSUBS 0.60fF $ **FLOATING
C6122 S.n5497 VSUBS 2.30fF $ **FLOATING
C6123 S.n5498 VSUBS 5.52fF $ **FLOATING
C6124 S.n5499 VSUBS 15.97fF $ **FLOATING
C6125 S.n5500 VSUBS 9.18fF $ **FLOATING
C6126 S.n5501 VSUBS 9.19fF $ **FLOATING
C6127 S.n5502 VSUBS 9.19fF $ **FLOATING
C6128 S.n5503 VSUBS 9.19fF $ **FLOATING
C6129 S.n5504 VSUBS 9.19fF $ **FLOATING
C6130 S.n5505 VSUBS 9.19fF $ **FLOATING
C6131 S.n5506 VSUBS 9.19fF $ **FLOATING
C6132 S.n5507 VSUBS 9.19fF $ **FLOATING
C6133 S.n5508 VSUBS 9.25fF $ **FLOATING
C6134 S.n5509 VSUBS 12.68fF $ **FLOATING
.ends

